PK
     w�O\���gm gm    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_0":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_1":["pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_1"],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_2":["pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_1"],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_3":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_4":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_5":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_6":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_7":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_8":["pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_1"],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_9":["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_1"],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_10":["pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_1"],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_11":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_12":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_13":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_14":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_15":["pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_0"],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_16":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_17":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_18":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_19":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_20":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_21":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_22":["pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_1"],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_23":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_24":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_25":["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_1"],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_26":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_27":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_28":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_29":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_30":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_31":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32":["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_2","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5"],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_33":[],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34":["pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_1","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0"],"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35":["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3"],"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0":["pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34"],"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_1":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_22"],"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2":["pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32"],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0":["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32"],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_1":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_25"],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2":["pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_0"],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_3":[],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_4":[],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_5":[],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6":["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0"],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35"],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_8":[],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_9":[],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_10":[],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_11":[],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_12":[],"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_13":[],"pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35"],"pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32"],"pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_2":[],"pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_3":[],"pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_4":[],"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_0":["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3"],"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_1":["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_4"],"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_2":["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5"],"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35"],"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4":["pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_1"],"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32"],"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0":["pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0"],"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_1":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_2"],"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2":["pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2"],"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0":["pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0"],"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_1":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_10"],"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2":["pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2"],"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0":["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0"],"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_1":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_8"],"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2":["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2"],"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0":["pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_0","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0"],"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_1":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_9"],"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2":["pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_2","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2"],"pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_0":["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0"],"pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_1":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_1"],"pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_2":["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2"],"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_0":["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3"],"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_1":["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_4"],"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_2":["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5"],"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3":["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_0"],"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_4":["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_1"],"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5":["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_2"],"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_0":["pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3"],"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_1":["pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_4"],"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_2":["pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5"],"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3":["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_0"],"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_4":["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_1"],"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5":["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_2"],"pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_0":[],"pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_1":[],"pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_2":[],"pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3":["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_0"],"pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_4":["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_1"],"pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5":["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_2"],"pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_0":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_15"],"pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_1":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34"],"pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_2":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32"],"pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_0":["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2"],"pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_1":["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4"]},"pin_to_color":{"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_0":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_1":"#C28C9F","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_2":"#FF74A3","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_3":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_4":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_5":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_6":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_7":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_8":"#FF029D","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_9":"#5FAD4E","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_10":"#683D3B","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_11":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_12":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_13":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_14":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_15":"#00AE7E","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_16":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_17":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_18":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_19":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_20":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_21":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_22":"#008F9C","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_23":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_24":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_25":"#FFE502","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_26":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_27":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_28":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_29":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_30":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_31":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32":"#BB8800","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_33":"#000000","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34":"#6A826C","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35":"#9E008E","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0":"#6A826C","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_1":"#008F9C","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2":"#BB8800","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0":"#BB8800","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_1":"#FFE502","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2":"#005F39","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_3":"#000000","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_4":"#000000","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_5":"#000000","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6":"#BB8800","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7":"#9E008E","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_8":"#000000","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_9":"#000000","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_10":"#000000","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_11":"#000000","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_12":"#000000","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_13":"#000000","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0":"#9E008E","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1":"#BB8800","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_2":"#000000","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_3":"#000000","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_4":"#000000","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_0":"#FE8900","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_1":"#95003A","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_2":"#BDC6FF","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3":"#9E008E","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4":"#7544B1","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5":"#BB8800","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0":"#6A826C","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_1":"#FF74A3","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2":"#BB8800","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0":"#6A826C","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_1":"#683D3B","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2":"#BB8800","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0":"#6A826C","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_1":"#FF029D","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2":"#BB8800","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0":"#6A826C","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_1":"#5FAD4E","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2":"#BB8800","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_0":"#6A826C","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_1":"#C28C9F","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_2":"#BB8800","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_0":"#01FFFE","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_1":"#FF937E","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_2":"#98FF52","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3":"#FE8900","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_4":"#95003A","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5":"#BDC6FF","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_0":"#A75740","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_1":"#001544","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_2":"#968AE8","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3":"#01FFFE","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_4":"#FF937E","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5":"#98FF52","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_0":"#000000","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_1":"#000000","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_2":"#000000","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3":"#A75740","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_4":"#001544","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5":"#968AE8","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_0":"#00AE7E","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_1":"#6A826C","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_2":"#BB8800","pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_0":"#005F39","pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_1":"#7544B1"},"pin_to_state":{"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_0":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_1":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_2":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_3":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_4":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_5":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_6":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_7":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_8":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_9":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_10":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_11":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_12":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_13":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_14":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_15":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_16":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_17":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_18":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_19":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_20":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_21":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_22":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_23":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_24":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_25":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_26":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_27":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_28":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_29":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_30":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_31":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_33":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34":"neutral","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35":"neutral","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0":"neutral","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_1":"neutral","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_1":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_3":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_4":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_5":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_8":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_9":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_10":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_11":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_12":"neutral","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_13":"neutral","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0":"neutral","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1":"neutral","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_2":"neutral","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_3":"neutral","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_4":"neutral","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_0":"neutral","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_1":"neutral","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_2":"neutral","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3":"neutral","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4":"neutral","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5":"neutral","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0":"neutral","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_1":"neutral","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2":"neutral","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0":"neutral","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_1":"neutral","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2":"neutral","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0":"neutral","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_1":"neutral","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2":"neutral","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0":"neutral","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_1":"neutral","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2":"neutral","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_0":"neutral","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_1":"neutral","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_2":"neutral","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_0":"neutral","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_1":"neutral","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_2":"neutral","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3":"neutral","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_4":"neutral","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5":"neutral","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_0":"neutral","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_1":"neutral","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_2":"neutral","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3":"neutral","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_4":"neutral","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5":"neutral","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_0":"neutral","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_1":"neutral","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_2":"neutral","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3":"neutral","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_4":"neutral","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5":"neutral","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_0":"neutral","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_1":"neutral","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_2":"neutral","pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_0":"neutral","pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_1":"neutral"},"next_color_idx":26,"wires_placed_in_order":[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7"],["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3"],["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5"],["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7"],["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35"],["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_25","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_1"],["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0"],["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4"],["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6"],["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_4","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_1"],["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_4","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_1"],["pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_4","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_1"],["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3"],["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3"],["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3"],["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5"],["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5"],["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5"],["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_2"],["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_0"],["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0"],["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2"],["pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0"],["pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2"],["pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0"],["pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2"],["pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0"],["pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_2"],["pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_1","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0"],["pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_15","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_0"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_1","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_1"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_22","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_1"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_9","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_1"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_8","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_1"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_10","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_1"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_2","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_1"],["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_2","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5"],["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_2","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5"],["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_0","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3"],["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_0","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3"],["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_0","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3"],["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_2","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5"],["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3"],["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32"],["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5"],["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2","pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_0"],["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4","pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_1"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7"]]],[[],[["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3"]]],[[],[["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5"]]],[[],[["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7"]]],[[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7"]],[]],[[],[["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35"]]],[[],[["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32"]]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_25","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_1"]]],[[],[["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0"]]],[[],[["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4"]]],[[],[["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6"]]],[[],[["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_4","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_1"]]],[[],[["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_4","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_1"]]],[[],[["pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_4","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_1"]]],[[],[["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3"]]],[[],[["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3"]]],[[],[["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3"]]],[[],[["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5"]]],[[],[["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5"]]],[[],[["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5"]]],[[],[["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_2"]]],[[],[["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_0"]]],[[],[["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0"]]],[[],[["pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2"]]],[[],[["pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0"]]],[[],[["pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2"]]],[[],[["pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0"]]],[[],[["pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2"]]],[[],[["pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0"]]],[[],[["pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2"]]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_2"]]],[[],[["pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_1","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34"]]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0"]]],[[],[["pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32"]]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_15","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_0"]]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_1","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_1"]]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_22","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_1"]]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_9","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_1"]]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_8","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_1"]]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_10","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_1"]]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_2","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_1"]]],[[["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5"]],[]],[[],[["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_2","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5"]]],[[["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5"]],[]],[[],[["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_2","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5"]]],[[["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3"]],[]],[[],[["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_0","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3"]]],[[["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3"]],[]],[[],[["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_0","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3"]]],[[["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3"]],[]],[[],[["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_0","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3"]]],[[["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5"]],[]],[[],[["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_2","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5"]]],[[["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6"]],[]],[[],[["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6"]]],[[["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7"]],[]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7"]]],[[["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3"]],[]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3"]]],[[["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0"]],[]],[[],[["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32"]]],[[["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5"]],[]],[[],[["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5"]]],[[],[["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2","pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_0"]]],[[],[["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4","pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_1"]]],[[["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2"]],[]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_0":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_1":"0000000000000009","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_2":"0000000000000014","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_3":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_4":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_5":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_6":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_7":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_8":"0000000000000012","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_9":"0000000000000011","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_10":"0000000000000013","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_11":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_12":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_13":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_14":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_15":"0000000000000007","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_16":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_17":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_18":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_19":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_20":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_21":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_22":"0000000000000010","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_23":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_24":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_25":"0000000000000001","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_26":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_27":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_28":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_29":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_30":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_31":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32":"0000000000000002","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_33":"_","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34":"0000000000000008","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35":"0000000000000000","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0":"0000000000000008","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_1":"0000000000000010","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2":"0000000000000002","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0":"0000000000000002","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_1":"0000000000000001","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2":"0000000000000003","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_3":"_","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_4":"_","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_5":"_","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6":"0000000000000002","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7":"0000000000000000","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_8":"_","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_9":"_","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_10":"_","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_11":"_","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_12":"_","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_13":"_","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0":"0000000000000000","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1":"0000000000000002","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_2":"_","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_3":"_","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_4":"_","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_0":"0000000000000019","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_1":"0000000000000004","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_2":"0000000000000020","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3":"0000000000000000","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4":"0000000000000021","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5":"0000000000000002","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0":"0000000000000008","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_1":"0000000000000014","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2":"0000000000000002","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0":"0000000000000008","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_1":"0000000000000013","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2":"0000000000000002","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0":"0000000000000008","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_1":"0000000000000012","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2":"0000000000000002","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0":"0000000000000008","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_1":"0000000000000011","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2":"0000000000000002","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_0":"0000000000000008","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_1":"0000000000000009","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_2":"0000000000000002","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_0":"0000000000000018","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_1":"0000000000000005","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_2":"0000000000000016","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3":"0000000000000019","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_4":"0000000000000004","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5":"0000000000000020","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_0":"0000000000000017","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_1":"0000000000000006","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_2":"0000000000000015","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3":"0000000000000018","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_4":"0000000000000005","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5":"0000000000000016","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_0":"_","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_1":"_","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_2":"_","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3":"0000000000000017","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_4":"0000000000000006","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5":"0000000000000015","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_0":"0000000000000007","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_1":"0000000000000008","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_2":"0000000000000002","pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_0":"0000000000000003","pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_1":"0000000000000021"},"component_id_to_pins":{"74acac88-bdbd-4cf8-a6d0-88a8e37e4339":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33","34","35"],"eec8f51a-d3bf-449e-8d78-eae90dc3b47b":["0","1","2"],"9f8a660b-abfe-4ab0-b928-17d164c70e91":["0","1","2","3","4","5","6","7","8","9","10","11","12","13"],"626afbb9-b6e8-484c-a0c9-73a3153bfa4b":["0","1","2","3","4"],"84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93":["0","1","2","3","4","5"],"b30c19b4-cbcc-4fcb-922a-41036c5c1597":["0","1","2"],"e05342e8-37ba-4805-9f10-65c175bc3b0a":["0","1","2"],"3370895a-3b84-4a37-962a-17eb943a9099":["0","1","2"],"c233f660-2a1e-47b6-a3be-9e7359335c8d":["0","1","2"],"6059ea10-2811-4e34-bdb0-f79b9ba26520":["0","1","2"],"e5987f7a-cd81-40fb-a133-7daaaf14ca65":["0","1","2","3","4","5"],"1de15ba4-c578-435f-a770-003084d8278c":["0","1","2","3","4","5"],"278bdbb6-15d7-48ca-b9a7-98b3768b8b53":["0","1","2","3","4","5"],"d559fc7a-7bf4-428e-897b-06b2c446b856":["0","1","2"],"8b1a8dd9-b28d-4698-be03-bc2e13b1280b":[],"cc2e085a-84a3-44a1-b00d-edfd81716ffb":[],"e34757b9-8443-454a-bfd1-8e46b2a1b931":[],"977fc553-9453-4974-bc2f-c5c683bde336":[],"373db5bb-f7db-4663-b1c6-ca837886b0ef":[],"d1480eaa-3e21-4494-97d1-a6d04570c0ee":["0","1"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3"],"0000000000000002":["pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_2","pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_2","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5"],"0000000000000001":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_25","pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_1"],"0000000000000003":["pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2","pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_0"],"0000000000000004":["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_4","pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_1"],"0000000000000005":["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_4","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_1"],"0000000000000006":["pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_4","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_1"],"0000000000000008":["pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_0","pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_1","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0"],"0000000000000007":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_15","pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_0"],"0000000000000009":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_1","pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_1"],"0000000000000010":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_22","pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_1"],"0000000000000011":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_9","pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_1"],"0000000000000012":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_8","pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_1"],"0000000000000013":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_10","pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_1"],"0000000000000014":["pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_2","pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_1"],"0000000000000015":["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_2","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5"],"0000000000000016":["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_2","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5"],"0000000000000017":["pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_0","pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3"],"0000000000000018":["pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_0","pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3"],"0000000000000019":["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_0","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3"],"0000000000000020":["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_2","pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5"],"0000000000000021":["pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4","pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_1"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000002":"Net 2","0000000000000001":"Net 1","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000008":"Net 8","0000000000000007":"Net 7","0000000000000009":"Net 9","0000000000000010":"Net 10","0000000000000011":"Net 11","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000014":"Net 14","0000000000000015":"Net 15","0000000000000016":"Net 16","0000000000000017":"Net 17","0000000000000018":"Net 18","0000000000000019":"Net 19","0000000000000020":"Net 20","0000000000000021":"Net 21"},"all_breadboard_info_list":[],"breadboard_info_list":[],"componentsData":[{"compProperties":{},"position":[1068.2708245,-721.1528079999999],"typeId":"8c62c73e-11cc-47e9-8a08-93f7b83d583d","componentVersion":1,"instanceId":"74acac88-bdbd-4cf8-a6d0-88a8e37e4339","orientation":"up","circleData":[[1142.5,-595],[1141.9236219999998,-609.9999999999999],[1142.5,-625],[1142.5,-640.576378],[1142.5,-654.9999999999999],[1142.4495655,-669.5673025],[1141.8732475000002,-684.553012],[1142.4495655,-699.5387199999999],[1142.4495655,-714.5244294999999],[1142.4495655,-729.5101974999999],[1142.4495655,-744.4959054999999],[1141.8732475000002,-758.9052355],[1141.2968695,-774.467323],[1142.4495655,-789.4530309999999],[1142.4495655,-805.0151185],[1142.4495655,-818.8481304999999],[1142.4495655,-833.2574604999999],[1142.4495655,-849.3959245],[993.7451769999999,-849.3959245],[993.7451769999999,-834.4102164999999],[993.1687989999999,-818.8481304999999],[993.1687989999999,-803.8624209999999],[993.1687989999999,-790.029409],[993.1687989999999,-773.890945],[993.1687989999999,-758.9052355],[992.592421,-743.9195275],[993.1687989999999,-730.0865739999999],[993.1687989999999,-713.9481024999999],[993.7451769999999,-700.1150905],[993.7451769999999,-684.553012],[993.1687989999999,-669.5673025],[993.1687989999999,-654.5815944999999],[992.592421,-639.5958864999999],[993.7451769999999,-624.6101185],[993.1687989999999,-610.2007869999999],[993.1687989999999,-594.638701]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1376.206567,-1008.6937404999996],"typeId":"3eb2c561-68ea-4550-951c-6dd736f5b9fe","componentVersion":1,"instanceId":"eec8f51a-d3bf-449e-8d78-eae90dc3b47b","orientation":"up","circleData":[[1307.5,-1014.9999999999999],[1306.9866535,-1004.3331369999999],[1306.9866535,-994.3346319999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1108.744858,-438.08225949999996],"typeId":"1e6e3ab1-f6ac-46c9-9e87-56073aaa4ed0","componentVersion":1,"instanceId":"9f8a660b-abfe-4ab0-b928-17d164c70e91","orientation":"up","circleData":[[1052.5,-415],[1072,-415],[1090.75,-415],[1111,-415],[1129,-415],[1147.75,-415],[1167.25,-415],[1052.5,-482.4999999999999],[1072,-482.4999999999999],[1090.75,-482.4999999999999],[1111,-482.4999999999999],[1129,-482.4999999999999],[1147.75,-482.4999999999999],[1167.25,-482.4999999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1562.5000000000005,-984.9999999999995],"typeId":"4d90ceac-9e99-4afa-997d-ea12d0bf78ab","componentVersion":2,"instanceId":"84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93","orientation":"left","circleData":[[1547.5000000000005,-939.9999999999998],[1562.5000000000005,-939.9999999999998],[1577.5000000000005,-939.9999999999998],[1547.5000000000005,-1029.9999999999998],[1562.5000000000005,-1029.9999999999998],[1577.5000000000005,-1029.9999999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1376.206567,-948.6937405000001],"typeId":"3eb2c561-68ea-4550-951c-6dd736f5b9fe","componentVersion":1,"instanceId":"b30c19b4-cbcc-4fcb-922a-41036c5c1597","orientation":"up","circleData":[[1307.5,-955.0000000000001],[1306.9866535,-944.3331370000001],[1306.9866535,-934.334632]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1376.206567,-813.6937404999999],"typeId":"3eb2c561-68ea-4550-951c-6dd736f5b9fe","componentVersion":1,"instanceId":"e05342e8-37ba-4805-9f10-65c175bc3b0a","orientation":"up","circleData":[[1307.5,-819.9999999999999],[1306.9866535,-809.3331369999999],[1306.9866535,-799.3346319999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1376.206567,-723.6937404999999],"typeId":"3eb2c561-68ea-4550-951c-6dd736f5b9fe","componentVersion":1,"instanceId":"3370895a-3b84-4a37-962a-17eb943a9099","orientation":"up","circleData":[[1307.5,-730],[1306.9866535,-719.3331369999999],[1306.9866535,-709.3346319999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1376.206567,-573.6937404999996],"typeId":"3eb2c561-68ea-4550-951c-6dd736f5b9fe","componentVersion":1,"instanceId":"c233f660-2a1e-47b6-a3be-9e7359335c8d","orientation":"up","circleData":[[1307.5,-580],[1306.9866535,-569.3331369999999],[1306.9866535,-559.3346319999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1376.206567,-513.6937404999994],"typeId":"3eb2c561-68ea-4550-951c-6dd736f5b9fe","componentVersion":1,"instanceId":"6059ea10-2811-4e34-bdb0-f79b9ba26520","orientation":"up","circleData":[[1307.5,-519.9999999999998],[1306.9866535,-509.3331369999996],[1306.9866535,-499.3346319999996]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1562.5,-835],"typeId":"4d90ceac-9e99-4afa-997d-ea12d0bf78ab","componentVersion":2,"instanceId":"e5987f7a-cd81-40fb-a133-7daaaf14ca65","orientation":"left","circleData":[[1547.5,-790],[1562.5,-790],[1577.5,-790],[1547.5,-880],[1562.5,-880],[1577.5,-880]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1562.5,-685],"typeId":"4d90ceac-9e99-4afa-997d-ea12d0bf78ab","componentVersion":2,"instanceId":"1de15ba4-c578-435f-a770-003084d8278c","orientation":"left","circleData":[[1547.5,-640],[1562.5,-640],[1577.5,-640],[1547.5,-730],[1562.5,-730],[1577.5,-730]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1562.5,-535],"typeId":"4d90ceac-9e99-4afa-997d-ea12d0bf78ab","componentVersion":2,"instanceId":"278bdbb6-15d7-48ca-b9a7-98b3768b8b53","orientation":"left","circleData":[[1547.5,-490],[1562.5,-490],[1577.5,-490],[1547.5,-580],[1562.5,-580],[1577.5,-580]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1037.4999640000005,-1000.3543165000002],"typeId":"8e39a87a-aa8b-4e7b-b4f9-ffb309d3bd6d","componentVersion":2,"instanceId":"d559fc7a-7bf4-428e-897b-06b2c446b856","orientation":"left","circleData":[[1127.5,-985.0000000000001],[1127.5,-1000.3543300000002],[1127.5,-1016.2992115000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"PIR AM312","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1373.3235491014825,-614.080843588187],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"8b1a8dd9-b28d-4698-be03-bc2e13b1280b","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"SN74AHCT125N","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1241.3991097837843,-446.1850055664984],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"cc2e085a-84a3-44a1-b00d-edfd81716ffb","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"FireBeetle ESP-WROOM-32","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1061.4755430072087,-531.2673966381285],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"977fc553-9453-4974-bc2f-c5c683bde336","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"WS2812B","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1558.1276439176888,-456.817243474783],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"373db5bb-f7db-4663-b1c6-ca837886b0ef","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[539.3530000000001,-828.1929999999998],"typeId":"17f8a068-7d39-4707-9d27-f81c9a96628b","componentVersion":1,"instanceId":"626afbb9-b6e8-484c-a0c9-73a3153bfa4b","orientation":"up","circleData":[[617.5,-580],[553.2280000000001,-591.865],[494.8870000000003,-586.9209999999999],[436.5475,-586.9209999999999],[377.2180000000002,-585.9325]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"HW-486","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1142.9260280148328,-1081.6169160446073],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"e34757b9-8443-454a-bfd1-8e46b2a1b931","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"325","displayFormat":"input","showOnComp":true,"isVisibleToUser":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true}},"position":[1312.9353646483635,-399.90486524040114],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"d1480eaa-3e21-4494-97d1-a6d04570c0ee","orientation":"up","circleData":[[1277.5,-400.00000000000006],[1352.5,-400]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-1133.69300","left":"263.85300","width":"1334.89700","height":"778.59812","x":"263.85300","y":"-1133.69300"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0\",\"endPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35\",\"rawStartPinId\":\"pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_0\",\"rawEndPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"617.5000000000_-580.0000000000\\\",\\\"617.5000000000_-505.0000000000\\\",\\\"947.5000000000_-505.0000000000\\\",\\\"947.5000000000_-595.0000000000\\\",\\\"977.8343995000_-595.0000000000\\\",\\\"977.8343995000_-594.6387010000\\\",\\\"993.1687990000_-594.6387010000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35\",\"endPinId\":\"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35\",\"rawEndPinId\":\"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"993.1687990000_-594.6387010000\\\",\\\"977.8343995000_-594.6387010000\\\",\\\"977.8343995000_-595.0000000000\\\",\\\"947.5000000000_-595.0000000000\\\",\\\"947.5000000000_-940.0000000000\\\",\\\"1187.5000000000_-940.0000000000\\\",\\\"1187.5000000000_-1090.0000000000\\\",\\\"1547.5000000000_-1090.0000000000\\\",\\\"1547.5000000000_-1030.0000000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35\",\"endPinId\":\"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_35\",\"rawEndPinId\":\"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"993.1687990000_-594.6387010000\\\",\\\"970.0000000000_-594.6387010000\\\",\\\"970.0000000000_-482.5000000000\\\",\\\"1052.5000000000_-482.5000000000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2\",\"endPinId\":\"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2\",\"rawStartPinId\":\"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2\",\"rawEndPinId\":\"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1306.9866535000_-709.3346320000\\\",\\\"1288.4933267500_-709.3346320000\\\",\\\"1288.4933267500_-707.5000000000\\\",\\\"1262.5000000000_-707.5000000000\\\",\\\"1262.5000000000_-557.5000000000\\\",\\\"1288.4933267500_-557.5000000000\\\",\\\"1288.4933267500_-559.3346320000\\\",\\\"1306.9866535000_-559.3346320000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2\",\"endPinId\":\"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2\",\"rawStartPinId\":\"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_2\",\"rawEndPinId\":\"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1306.9866535000_-709.3346320000\\\",\\\"1288.4933267500_-709.3346320000\\\",\\\"1288.4933267500_-707.5000000000\\\",\\\"1262.5000000000_-707.5000000000\\\",\\\"1262.5000000000_-797.5000000000\\\",\\\"1288.4933267500_-797.5000000000\\\",\\\"1288.4933267500_-799.3346320000\\\",\\\"1306.9866535000_-799.3346320000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_2\",\"endPinId\":\"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2\",\"rawStartPinId\":\"pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_2\",\"rawEndPinId\":\"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1306.9866535000_-499.3346320000\\\",\\\"1270.0000000000_-499.3346320000\\\",\\\"1270.0000000000_-559.3346320000\\\",\\\"1306.9866535000_-559.3346320000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1\",\"endPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32\",\"rawStartPinId\":\"pin-type-component_626afbb9-b6e8-484c-a0c9-73a3153bfa4b_1\",\"rawEndPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"553.2280000000_-591.8650000000\\\",\\\"553.2280000000_-552.1825000000\\\",\\\"550.0000000000_-552.1825000000\\\",\\\"550.0000000000_-482.5000000000\\\",\\\"741.2500000000_-482.5000000000\\\",\\\"741.2500000000_-497.5000000000\\\",\\\"932.5000000000_-497.5000000000\\\",\\\"932.5000000000_-640.0000000000\\\",\\\"977.5462105000_-640.0000000000\\\",\\\"977.5462105000_-639.5958865000\\\",\\\"992.5924210000_-639.5958865000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32\",\"endPinId\":\"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32\",\"rawEndPinId\":\"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5924210000_-639.5958865000\\\",\\\"977.5462105000_-639.5958865000\\\",\\\"977.5462105000_-640.0000000000\\\",\\\"932.5000000000_-640.0000000000\\\",\\\"932.5000000000_-925.0000000000\\\",\\\"1202.5000000000_-925.0000000000\\\",\\\"1202.5000000000_-1105.0000000000\\\",\\\"1577.5000000000_-1105.0000000000\\\",\\\"1577.5000000000_-1030.0000000000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32\",\"endPinId\":\"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32\",\"rawEndPinId\":\"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5924210000_-639.5958865000\\\",\\\"977.5462105000_-639.5958865000\\\",\\\"977.5462105000_-640.0000000000\\\",\\\"932.5000000000_-640.0000000000\\\",\\\"932.5000000000_-415.0000000000\\\",\\\"1052.5000000000_-415.0000000000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32\",\"endPinId\":\"pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_2\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32\",\"rawEndPinId\":\"pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5924210000_-639.5958865000\\\",\\\"977.5462105000_-639.5958865000\\\",\\\"977.5462105000_-640.0000000000\\\",\\\"932.5000000000_-640.0000000000\\\",\\\"932.5000000000_-910.0000000000\\\",\\\"1157.5000000000_-910.0000000000\\\",\\\"1157.5000000000_-1015.0000000000\\\",\\\"1138.7500000000_-1015.0000000000\\\",\\\"1138.7500000000_-1016.2992115000\\\",\\\"1127.5000000000_-1016.2992115000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32\",\"endPinId\":\"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_32\",\"rawEndPinId\":\"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5924210000_-639.5958865000\\\",\\\"977.5462105000_-639.5958865000\\\",\\\"977.5462105000_-640.0000000000\\\",\\\"955.0000000000_-640.0000000000\\\",\\\"955.0000000000_-932.5000000000\\\",\\\"1210.0000000000_-932.5000000000\\\",\\\"1210.0000000000_-992.5000000000\\\",\\\"1288.4933267500_-992.5000000000\\\",\\\"1288.4933267500_-994.3346320000\\\",\\\"1306.9866535000_-994.3346320000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0\",\"endPinId\":\"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6\",\"rawStartPinId\":\"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_0\",\"rawEndPinId\":\"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1052.5000000000_-415.0000000000\\\",\\\"1052.5000000000_-377.5000000000\\\",\\\"1165.0000000000_-377.5000000000\\\",\\\"1165.0000000000_-415.0000000000\\\",\\\"1167.2500000000_-415.0000000000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2\",\"endPinId\":\"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2\",\"rawStartPinId\":\"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2\",\"rawEndPinId\":\"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1306.9866535000_-934.3346320000\\\",\\\"1288.4933267500_-934.3346320000\\\",\\\"1288.4933267500_-932.5000000000\\\",\\\"1262.5000000000_-932.5000000000\\\",\\\"1262.5000000000_-797.5000000000\\\",\\\"1288.4933267500_-797.5000000000\\\",\\\"1288.4933267500_-799.3346320000\\\",\\\"1306.9866535000_-799.3346320000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2\",\"endPinId\":\"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2\",\"rawStartPinId\":\"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_2\",\"rawEndPinId\":\"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1306.9866535000_-934.3346320000\\\",\\\"1288.4933267500_-934.3346320000\\\",\\\"1288.4933267500_-932.5000000000\\\",\\\"1262.5000000000_-932.5000000000\\\",\\\"1262.5000000000_-992.5000000000\\\",\\\"1288.4933267500_-992.5000000000\\\",\\\"1288.4933267500_-994.3346320000\\\",\\\"1306.9866535000_-994.3346320000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_25\",\"endPinId\":\"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_1\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_25\",\"rawEndPinId\":\"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5924210000_-743.9195275000\\\",\\\"977.5462105000_-743.9195275000\\\",\\\"977.5462105000_-745.0000000000\\\",\\\"872.5000000000_-745.0000000000\\\",\\\"872.5000000000_-340.0000000000\\\",\\\"1075.0000000000_-340.0000000000\\\",\\\"1075.0000000000_-381.2500000000\\\",\\\"1072.0000000000_-381.2500000000\\\",\\\"1072.0000000000_-415.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2\",\"endPinId\":\"pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_0\",\"rawStartPinId\":\"pin-type-component_9f8a660b-abfe-4ab0-b928-17d164c70e91_2\",\"rawEndPinId\":\"pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1090.7500000000_-415.0000000000\\\",\\\"1090.7500000000_-400.0000000000\\\",\\\"1277.5000000000_-400.0000000000\\\"]}\"}","{\"color\":\"#7544B1\",\"startPinId\":\"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4\",\"endPinId\":\"pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_1\",\"rawStartPinId\":\"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_4\",\"rawEndPinId\":\"pin-type-component_d1480eaa-3e21-4494-97d1-a6d04570c0ee_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1562.5000000000_-1030.0000000000\\\",\\\"1562.5000000000_-1045.0000000000\\\",\\\"1607.5000000000_-1045.0000000000\\\",\\\"1607.5000000000_-400.0000000000\\\",\\\"1352.5000000000_-400.0000000000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_1\",\"endPinId\":\"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_4\",\"rawStartPinId\":\"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_1\",\"rawEndPinId\":\"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1562.5000000000_-940.0000000000\\\",\\\"1562.5000000000_-880.0000000000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_4\",\"endPinId\":\"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_1\",\"rawStartPinId\":\"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_4\",\"rawEndPinId\":\"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1562.5000000000_-730.0000000000\\\",\\\"1562.5000000000_-790.0000000000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_1\",\"endPinId\":\"pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_4\",\"rawStartPinId\":\"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_1\",\"rawEndPinId\":\"pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1562.5000000000_-640.0000000000\\\",\\\"1562.5000000000_-580.0000000000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0\",\"endPinId\":\"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0\",\"rawStartPinId\":\"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0\",\"rawEndPinId\":\"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1307.5000000000_-730.0000000000\\\",\\\"1247.5000000000_-730.0000000000\\\",\\\"1247.5000000000_-580.0000000000\\\",\\\"1307.5000000000_-580.0000000000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0\",\"endPinId\":\"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0\",\"rawStartPinId\":\"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_0\",\"rawEndPinId\":\"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1307.5000000000_-730.0000000000\\\",\\\"1247.5000000000_-730.0000000000\\\",\\\"1247.5000000000_-820.0000000000\\\",\\\"1307.5000000000_-820.0000000000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_0\",\"endPinId\":\"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0\",\"rawStartPinId\":\"pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_0\",\"rawEndPinId\":\"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1307.5000000000_-520.0000000000\\\",\\\"1270.0000000000_-520.0000000000\\\",\\\"1270.0000000000_-580.0000000000\\\",\\\"1307.5000000000_-580.0000000000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34\",\"endPinId\":\"pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_1\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34\",\"rawEndPinId\":\"pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"993.1687990000_-610.2007870000\\\",\\\"977.8343995000_-610.2007870000\\\",\\\"977.8343995000_-610.0000000000\\\",\\\"917.5000000000_-610.0000000000\\\",\\\"917.5000000000_-1060.0000000000\\\",\\\"1172.5000000000_-1060.0000000000\\\",\\\"1172.5000000000_-1000.0000000000\\\",\\\"1138.7500000000_-1000.0000000000\\\",\\\"1138.7500000000_-1000.3543300000\\\",\\\"1127.5000000000_-1000.3543300000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34\",\"endPinId\":\"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_34\",\"rawEndPinId\":\"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"993.1687990000_-610.2007870000\\\",\\\"977.8343995000_-610.2007870000\\\",\\\"977.8343995000_-610.0000000000\\\",\\\"917.5000000000_-610.0000000000\\\",\\\"917.5000000000_-1060.0000000000\\\",\\\"1262.5000000000_-1060.0000000000\\\",\\\"1262.5000000000_-1015.0000000000\\\",\\\"1307.5000000000_-1015.0000000000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0\",\"endPinId\":\"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0\",\"rawStartPinId\":\"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0\",\"rawEndPinId\":\"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1307.5000000000_-955.0000000000\\\",\\\"1247.5000000000_-955.0000000000\\\",\\\"1247.5000000000_-820.0000000000\\\",\\\"1307.5000000000_-820.0000000000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0\",\"endPinId\":\"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0\",\"rawStartPinId\":\"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_0\",\"rawEndPinId\":\"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1307.5000000000_-955.0000000000\\\",\\\"1247.5000000000_-955.0000000000\\\",\\\"1247.5000000000_-1015.0000000000\\\",\\\"1307.5000000000_-1015.0000000000\\\"]}\"}","{\"color\":\"#00AE7E\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_15\",\"endPinId\":\"pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_0\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_15\",\"rawEndPinId\":\"pin-type-component_d559fc7a-7bf4-428e-897b-06b2c446b856_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.4495655000_-818.8481305000\\\",\\\"1172.5000000000_-818.8481305000\\\",\\\"1172.5000000000_-985.0000000000\\\",\\\"1127.5000000000_-985.0000000000\\\"]}\"}","{\"color\":\"#C28C9F\",\"startPinId\":\"pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_1\",\"endPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_1\",\"rawStartPinId\":\"pin-type-component_6059ea10-2811-4e34-bdb0-f79b9ba26520_1\",\"rawEndPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1306.9866535000_-509.3331370000\\\",\\\"1288.4933267500_-509.3331370000\\\",\\\"1288.4933267500_-512.5000000000\\\",\\\"1172.5000000000_-512.5000000000\\\",\\\"1172.5000000000_-610.0000000000\\\",\\\"1141.9236220000_-610.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_22\",\"endPinId\":\"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_1\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_22\",\"rawEndPinId\":\"pin-type-component_eec8f51a-d3bf-449e-8d78-eae90dc3b47b_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"993.1687990000_-790.0294090000\\\",\\\"962.5000000000_-790.0294090000\\\",\\\"962.5000000000_-917.5000000000\\\",\\\"1255.0000000000_-917.5000000000\\\",\\\"1255.0000000000_-1007.5000000000\\\",\\\"1288.4933267500_-1007.5000000000\\\",\\\"1288.4933267500_-1004.3331370000\\\",\\\"1306.9866535000_-1004.3331370000\\\"]}\"}","{\"color\":\"#5FAD4E\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_9\",\"endPinId\":\"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_1\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_9\",\"rawEndPinId\":\"pin-type-component_c233f660-2a1e-47b6-a3be-9e7359335c8d_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.4495655000_-729.5101975000\\\",\\\"1157.4747827500_-729.5101975000\\\",\\\"1157.4747827500_-730.0000000000\\\",\\\"1240.0000000000_-730.0000000000\\\",\\\"1240.0000000000_-572.5000000000\\\",\\\"1288.4933267500_-572.5000000000\\\",\\\"1288.4933267500_-569.3331370000\\\",\\\"1306.9866535000_-569.3331370000\\\"]}\"}","{\"color\":\"#FF029D\",\"startPinId\":\"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_1\",\"endPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_8\",\"rawStartPinId\":\"pin-type-component_3370895a-3b84-4a37-962a-17eb943a9099_1\",\"rawEndPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_8\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1306.9866535000_-719.3331370000\\\",\\\"1288.4933267500_-719.3331370000\\\",\\\"1288.4933267500_-722.5000000000\\\",\\\"1157.4747827500_-722.5000000000\\\",\\\"1157.4747827500_-714.5244295000\\\",\\\"1142.4495655000_-714.5244295000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_10\",\"endPinId\":\"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_1\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_10\",\"rawEndPinId\":\"pin-type-component_e05342e8-37ba-4805-9f10-65c175bc3b0a_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.4495655000_-744.4959055000\\\",\\\"1172.5000000000_-744.4959055000\\\",\\\"1172.5000000000_-812.5000000000\\\",\\\"1288.4933267500_-812.5000000000\\\",\\\"1288.4933267500_-809.3331370000\\\",\\\"1306.9866535000_-809.3331370000\\\"]}\"}","{\"color\":\"#FF74A3\",\"startPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_2\",\"endPinId\":\"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_1\",\"rawStartPinId\":\"pin-type-component_74acac88-bdbd-4cf8-a6d0-88a8e37e4339_2\",\"rawEndPinId\":\"pin-type-component_b30c19b4-cbcc-4fcb-922a-41036c5c1597_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.5000000000_-625.0000000000\\\",\\\"1232.5000000000_-625.0000000000\\\",\\\"1232.5000000000_-947.5000000000\\\",\\\"1288.4933267500_-947.5000000000\\\",\\\"1288.4933267500_-944.3331370000\\\",\\\"1306.9866535000_-944.3331370000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_2\",\"endPinId\":\"pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5\",\"rawStartPinId\":\"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_2\",\"rawEndPinId\":\"pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1577.5000000000_-640.0000000000\\\",\\\"1577.5000000000_-580.0000000000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5\",\"endPinId\":\"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_2\",\"rawStartPinId\":\"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_5\",\"rawEndPinId\":\"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1577.5000000000_-730.0000000000\\\",\\\"1577.5000000000_-790.0000000000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_0\",\"endPinId\":\"pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3\",\"rawStartPinId\":\"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_0\",\"rawEndPinId\":\"pin-type-component_278bdbb6-15d7-48ca-b9a7-98b3768b8b53_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1547.5000000000_-640.0000000000\\\",\\\"1547.5000000000_-580.0000000000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3\",\"endPinId\":\"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_0\",\"rawStartPinId\":\"pin-type-component_1de15ba4-c578-435f-a770-003084d8278c_3\",\"rawEndPinId\":\"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1547.5000000000_-730.0000000000\\\",\\\"1547.5000000000_-790.0000000000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_0\",\"endPinId\":\"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3\",\"rawStartPinId\":\"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_0\",\"rawEndPinId\":\"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1547.5000000000_-940.0000000000\\\",\\\"1547.5000000000_-880.0000000000\\\"]}\"}","{\"color\":\"#BDC6FF\",\"startPinId\":\"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_2\",\"endPinId\":\"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5\",\"rawStartPinId\":\"pin-type-component_84e3c7b5-7dfd-4f6a-bb61-ad974b9e9f93_2\",\"rawEndPinId\":\"pin-type-component_e5987f7a-cd81-40fb-a133-7daaaf14ca65_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1577.5000000000_-940.0000000000\\\",\\\"1577.5000000000_-880.0000000000\\\"]}\"}"],"projectDescription":""}PK
     w�O\               jsons/PK
     w�O\�'���d  �d     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"FireBeetle ESP32","category":["User Defined"],"id":"8c62c73e-11cc-47e9-8a08-93f7b83d583d","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"03bee633-62f2-4ed0-b5c1-e772de98cfcb.png","iconPic":"85ff3ff6-223b-4d64-b6b1-3b6b2877ae4f.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"11.41732","numDisplayRows":"22.83465","pins":[{"uniquePinIdString":"0","positionMil":"1065.72717,300.71378","isAnchorPin":true,"label":"RST/EN"},{"uniquePinIdString":"1","positionMil":"1061.88465,400.71378","isAnchorPin":false,"label":"LRCK/IO17"},{"uniquePinIdString":"2","positionMil":"1065.72717,500.71378","isAnchorPin":false,"label":"DI/IO16"},{"uniquePinIdString":"3","positionMil":"1065.72717,604.55630","isAnchorPin":false,"label":"DO/IO4"},{"uniquePinIdString":"4","positionMil":"1065.72717,700.71378","isAnchorPin":false,"label":"MCLK/IO12"},{"uniquePinIdString":"5","positionMil":"1065.39094,797.82913","isAnchorPin":false,"label":"BCLK/IO14"},{"uniquePinIdString":"6","positionMil":"1061.54882,897.73386","isAnchorPin":false,"label":"SCL/IO22"},{"uniquePinIdString":"7","positionMil":"1065.39094,997.63858","isAnchorPin":false,"label":"SDA/IO21"},{"uniquePinIdString":"8","positionMil":"1065.39094,1097.54331","isAnchorPin":false,"label":"MISO/IO19"},{"uniquePinIdString":"9","positionMil":"1065.39094,1197.44843","isAnchorPin":false,"label":"MOSI/IO23"},{"uniquePinIdString":"10","positionMil":"1065.39094,1297.35315","isAnchorPin":false,"label":"SCK/IO18"},{"uniquePinIdString":"11","positionMil":"1061.54882,1393.41535","isAnchorPin":false,"label":"IO0"},{"uniquePinIdString":"12","positionMil":"1057.70630,1497.16260","isAnchorPin":false,"label":"NC"},{"uniquePinIdString":"13","positionMil":"1065.39094,1597.06732","isAnchorPin":false,"label":"A4/IO15"},{"uniquePinIdString":"14","positionMil":"1065.39094,1700.81457","isAnchorPin":false,"label":"A3/IO35"},{"uniquePinIdString":"15","positionMil":"1065.39094,1793.03465","isAnchorPin":false,"label":"A2/IO34"},{"uniquePinIdString":"16","positionMil":"1065.39094,1889.09685","isAnchorPin":false,"label":"A1/IO39/SENSOR_VN"},{"uniquePinIdString":"17","positionMil":"1065.39094,1996.68661","isAnchorPin":false,"label":"A0/IO36/SENSOR_VP"},{"uniquePinIdString":"18","positionMil":"74.02835,1996.68661","isAnchorPin":false,"label":"D0/IO3/RXD"},{"uniquePinIdString":"19","positionMil":"74.02835,1896.78189","isAnchorPin":false,"label":"D1/IO1/TXD"},{"uniquePinIdString":"20","positionMil":"70.18583,1793.03465","isAnchorPin":false,"label":"D2/IO25"},{"uniquePinIdString":"21","positionMil":"70.18583,1693.12992","isAnchorPin":false,"label":"D3/IO26"},{"uniquePinIdString":"22","positionMil":"70.18583,1600.90984","isAnchorPin":false,"label":"D4/IO27"},{"uniquePinIdString":"23","positionMil":"70.18583,1493.32008","isAnchorPin":false,"label":"D5/IO9/SD2"},{"uniquePinIdString":"24","positionMil":"70.18583,1393.41535","isAnchorPin":false,"label":"D6/IO10/SD3"},{"uniquePinIdString":"25","positionMil":"66.34331,1293.51063","isAnchorPin":false,"label":"D7/IO13"},{"uniquePinIdString":"26","positionMil":"70.18583,1201.29094","isAnchorPin":false,"label":"D8/IO5"},{"uniquePinIdString":"27","positionMil":"70.18583,1093.70113","isAnchorPin":false,"label":"D9/IO2"},{"uniquePinIdString":"28","positionMil":"74.02835,1001.48105","isAnchorPin":false,"label":"IO6/CLK"},{"uniquePinIdString":"29","positionMil":"74.02835,897.73386","isAnchorPin":false,"label":"IO7/SD0"},{"uniquePinIdString":"30","positionMil":"70.18583,797.82913","isAnchorPin":false,"label":"IO8/SD1"},{"uniquePinIdString":"31","positionMil":"70.18583,697.92441","isAnchorPin":false,"label":"IO11/SMD"},{"uniquePinIdString":"32","positionMil":"66.34331,598.01969","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"33","positionMil":"74.02835,498.11457","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"34","positionMil":"70.18583,402.05236","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"35","positionMil":"70.18583,298.30512","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"HC-SR505 Mini PIR Motion Sensing Module","category":["User Defined"],"id":"3eb2c561-68ea-4550-951c-6dd736f5b9fe","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"bb2d2ee4-fa83-49b1-89fe-70727f49c778.png","iconPic":"32487380-bef1-4e4f-8e56-19d5eed1120c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"11.81102","numDisplayRows":"7.87402","pins":[{"uniquePinIdString":"0","positionMil":"132.50722,435.74273","isAnchorPin":true,"label":"+"},{"uniquePinIdString":"1","positionMil":"129.08491,364.63031","isAnchorPin":false,"label":"out"},{"uniquePinIdString":"2","positionMil":"129.08491,297.97361","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"SN74AHCT125N ","category":["User Defined"],"id":"1e6e3ab1-f6ac-46c9-9e87-56073aaa4ed0","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"3d684ffe-1f74-462a-8eb5-42254bda90cd.png","iconPic":"6fad6c1f-1fec-41b3-8a64-12aeedea4fac.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"18.74539","numDisplayRows":"9.73165","pins":[{"uniquePinIdString":"0","positionMil":"562.30378,332.70077","isAnchorPin":true,"label":"1OE"},{"uniquePinIdString":"1","positionMil":"692.30378,332.70077","isAnchorPin":false,"label":"1A"},{"uniquePinIdString":"2","positionMil":"817.30378,332.70077","isAnchorPin":false,"label":"1Y"},{"uniquePinIdString":"3","positionMil":"952.30378,332.70077","isAnchorPin":false,"label":"2OE"},{"uniquePinIdString":"4","positionMil":"1072.30378,332.70077","isAnchorPin":false,"label":"2A"},{"uniquePinIdString":"5","positionMil":"1197.30378,332.70077","isAnchorPin":false,"label":"2Y"},{"uniquePinIdString":"6","positionMil":"1327.30378,332.70077","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"562.30378,782.70077","isAnchorPin":false,"label":"Vcc"},{"uniquePinIdString":"8","positionMil":"692.30378,782.70077","isAnchorPin":false,"label":"4OE"},{"uniquePinIdString":"9","positionMil":"817.30378,782.70077","isAnchorPin":false,"label":"4A"},{"uniquePinIdString":"10","positionMil":"952.30378,782.70077","isAnchorPin":false,"label":"4Y"},{"uniquePinIdString":"11","positionMil":"1072.30378,782.70077","isAnchorPin":false,"label":"3OE"},{"uniquePinIdString":"12","positionMil":"1197.30378,782.70077","isAnchorPin":false,"label":"3A"},{"uniquePinIdString":"13","positionMil":"1327.30378,782.70077","isAnchorPin":false,"label":"3Y"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"WS2812B LED","category":["User Defined"],"id":"4d90ceac-9e99-4afa-997d-ea12d0bf78ab","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"80e9010a-c477-4737-bb01-43c9d75c1ab5.png","iconPic":"6a650d67-2f6f-4705-ba20-a1e007a57e5c.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.50000","numDisplayRows":"3.50000","pins":[{"uniquePinIdString":"0","positionMil":"25.00000,275.00000","isAnchorPin":true,"label":"+5V"},{"uniquePinIdString":"1","positionMil":"25.00000,175.00000","isAnchorPin":false,"label":"DO"},{"uniquePinIdString":"2","positionMil":"25.00000,75.00000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"3","positionMil":"625.00000,275.00000","isAnchorPin":false,"label":"+5V"},{"uniquePinIdString":"4","positionMil":"625.00000,175.00000","isAnchorPin":false,"label":"Din"},{"uniquePinIdString":"5","positionMil":"625.00000,75.00000","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"HC-SR505 Mini PIR Motion Sensing Module","category":["User Defined"],"id":"3eb2c561-68ea-4550-951c-6dd736f5b9fe","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"bb2d2ee4-fa83-49b1-89fe-70727f49c778.png","iconPic":"32487380-bef1-4e4f-8e56-19d5eed1120c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"11.81102","numDisplayRows":"7.87402","pins":[{"uniquePinIdString":"0","positionMil":"132.50722,435.74273","isAnchorPin":true,"label":"+"},{"uniquePinIdString":"1","positionMil":"129.08491,364.63031","isAnchorPin":false,"label":"out"},{"uniquePinIdString":"2","positionMil":"129.08491,297.97361","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"HC-SR505 Mini PIR Motion Sensing Module","category":["User Defined"],"id":"3eb2c561-68ea-4550-951c-6dd736f5b9fe","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"bb2d2ee4-fa83-49b1-89fe-70727f49c778.png","iconPic":"32487380-bef1-4e4f-8e56-19d5eed1120c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"11.81102","numDisplayRows":"7.87402","pins":[{"uniquePinIdString":"0","positionMil":"132.50722,435.74273","isAnchorPin":true,"label":"+"},{"uniquePinIdString":"1","positionMil":"129.08491,364.63031","isAnchorPin":false,"label":"out"},{"uniquePinIdString":"2","positionMil":"129.08491,297.97361","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"HC-SR505 Mini PIR Motion Sensing Module","category":["User Defined"],"id":"3eb2c561-68ea-4550-951c-6dd736f5b9fe","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"bb2d2ee4-fa83-49b1-89fe-70727f49c778.png","iconPic":"32487380-bef1-4e4f-8e56-19d5eed1120c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"11.81102","numDisplayRows":"7.87402","pins":[{"uniquePinIdString":"0","positionMil":"132.50722,435.74273","isAnchorPin":true,"label":"+"},{"uniquePinIdString":"1","positionMil":"129.08491,364.63031","isAnchorPin":false,"label":"out"},{"uniquePinIdString":"2","positionMil":"129.08491,297.97361","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"HC-SR505 Mini PIR Motion Sensing Module","category":["User Defined"],"id":"3eb2c561-68ea-4550-951c-6dd736f5b9fe","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"bb2d2ee4-fa83-49b1-89fe-70727f49c778.png","iconPic":"32487380-bef1-4e4f-8e56-19d5eed1120c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"11.81102","numDisplayRows":"7.87402","pins":[{"uniquePinIdString":"0","positionMil":"132.50722,435.74273","isAnchorPin":true,"label":"+"},{"uniquePinIdString":"1","positionMil":"129.08491,364.63031","isAnchorPin":false,"label":"out"},{"uniquePinIdString":"2","positionMil":"129.08491,297.97361","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"HC-SR505 Mini PIR Motion Sensing Module","category":["User Defined"],"id":"3eb2c561-68ea-4550-951c-6dd736f5b9fe","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"bb2d2ee4-fa83-49b1-89fe-70727f49c778.png","iconPic":"32487380-bef1-4e4f-8e56-19d5eed1120c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"11.81102","numDisplayRows":"7.87402","pins":[{"uniquePinIdString":"0","positionMil":"132.50722,435.74273","isAnchorPin":true,"label":"+"},{"uniquePinIdString":"1","positionMil":"129.08491,364.63031","isAnchorPin":false,"label":"out"},{"uniquePinIdString":"2","positionMil":"129.08491,297.97361","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"WS2812B LED","category":["User Defined"],"id":"4d90ceac-9e99-4afa-997d-ea12d0bf78ab","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"80e9010a-c477-4737-bb01-43c9d75c1ab5.png","iconPic":"6a650d67-2f6f-4705-ba20-a1e007a57e5c.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.50000","numDisplayRows":"3.50000","pins":[{"uniquePinIdString":"0","positionMil":"25.00000,275.00000","isAnchorPin":true,"label":"+5V"},{"uniquePinIdString":"1","positionMil":"25.00000,175.00000","isAnchorPin":false,"label":"DO"},{"uniquePinIdString":"2","positionMil":"25.00000,75.00000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"3","positionMil":"625.00000,275.00000","isAnchorPin":false,"label":"+5V"},{"uniquePinIdString":"4","positionMil":"625.00000,175.00000","isAnchorPin":false,"label":"Din"},{"uniquePinIdString":"5","positionMil":"625.00000,75.00000","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"WS2812B LED","category":["User Defined"],"id":"4d90ceac-9e99-4afa-997d-ea12d0bf78ab","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"80e9010a-c477-4737-bb01-43c9d75c1ab5.png","iconPic":"6a650d67-2f6f-4705-ba20-a1e007a57e5c.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.50000","numDisplayRows":"3.50000","pins":[{"uniquePinIdString":"0","positionMil":"25.00000,275.00000","isAnchorPin":true,"label":"+5V"},{"uniquePinIdString":"1","positionMil":"25.00000,175.00000","isAnchorPin":false,"label":"DO"},{"uniquePinIdString":"2","positionMil":"25.00000,75.00000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"3","positionMil":"625.00000,275.00000","isAnchorPin":false,"label":"+5V"},{"uniquePinIdString":"4","positionMil":"625.00000,175.00000","isAnchorPin":false,"label":"Din"},{"uniquePinIdString":"5","positionMil":"625.00000,75.00000","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"WS2812B LED","category":["User Defined"],"id":"4d90ceac-9e99-4afa-997d-ea12d0bf78ab","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"80e9010a-c477-4737-bb01-43c9d75c1ab5.png","iconPic":"6a650d67-2f6f-4705-ba20-a1e007a57e5c.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.50000","numDisplayRows":"3.50000","pins":[{"uniquePinIdString":"0","positionMil":"25.00000,275.00000","isAnchorPin":true,"label":"+5V"},{"uniquePinIdString":"1","positionMil":"25.00000,175.00000","isAnchorPin":false,"label":"DO"},{"uniquePinIdString":"2","positionMil":"25.00000,75.00000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"3","positionMil":"625.00000,275.00000","isAnchorPin":false,"label":"+5V"},{"uniquePinIdString":"4","positionMil":"625.00000,175.00000","isAnchorPin":false,"label":"Din"},{"uniquePinIdString":"5","positionMil":"625.00000,75.00000","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"KY-018 LDR Photo Resistor","category":["User Defined"],"id":"8e39a87a-aa8b-4e7b-b4f9-ffb309d3bd6d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"a65aebfd-90e6-4215-8cb5-f5692b012cc2.png","iconPic":"7e39c2f4-a1af-49ff-bc26-783004b83469.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"5.90551","numDisplayRows":"12.59843","pins":[{"uniquePinIdString":"0","positionMil":"192.91339,29.92126","isAnchorPin":true,"label":"Signal"},{"uniquePinIdString":"1","positionMil":"295.27559,29.92126","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"401.57480,29.92126","isAnchorPin":false,"label":"Ground"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"5V PSU","category":["User Defined"],"id":"17f8a068-7d39-4707-9d27-f81c9a96628b","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"90a26a0e-dc54-4725-bfe3-cfd4e64c35ea.png","iconPic":"5c3bf32d-6880-4472-891e-2d4d904f1ad6.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"35.40000","numDisplayRows":"39.40000","pins":[{"uniquePinIdString":"0","positionMil":"2290.98000,315.38000","isAnchorPin":true,"label":"V+"},{"uniquePinIdString":"1","positionMil":"1862.50000,394.48000","isAnchorPin":false,"label":"V-"},{"uniquePinIdString":"2","positionMil":"1473.56000,361.52000","isAnchorPin":false,"label":"Ground"},{"uniquePinIdString":"3","positionMil":"1084.63000,361.52000","isAnchorPin":false,"label":"Neutral"},{"uniquePinIdString":"4","positionMil":"689.10000,354.93000","isAnchorPin":false,"label":"Line"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     w�O\               images/PK
     w�O\��;�. �. /   images/03bee633-62f2-4ed0-b5c1-e772de98cfcb.png�PNG

   IHDR  -  d   D\w�   	pHYs  �  ��+  ��IDATx���Wy6��ܺw{/�wY���䎻�T�@H�R(	!�H����!@h6c���ɶ,Y�,�$����j����g��=g���ծ�y~��{gΜ93��g��=oq��`Gc#^z�%��=:::p!cڴ���/�$I��(�`�6\*(..Ư~�3�����BFMM,���z˗/K�ƭ��F�x��g�����͸PZR���3x�_��s��b�_�ŗ1e�t\�hkk��Ǐ��k��g?����mm�z��W��_���8.&��t���f�bi9pp��ر㌸~�5�/}�����>NZ��������#,\� ������~;�,Yll�����8z�(8p�`<���_��יP�=����m�ݻ�ǦM������Q�7oƽ���?�_~�e�:p���x	Vw�}dY����8p0��}�v�:u�'O����i�OPWW���̟���'�QPZ���O��`(���Gb8pp�@�$�74`������;�·ǽU��U���b߾}F���X��]��F����"�y�*ܲ�Jԕ((���xd�!�n$v�x=��ēoǳ�<�o���ᮻ��u��P��E��E��@R�ǁ*�����F�q�Z�y��~�ݻv���ɳ!���&-�ǋ��R���?����}+�oX�I**�+��������)ذ�ϼ�*Ξm�����p�5W�wߊ��A�MXw����K�k��>����'�q�e�ѣO��;����ӰH�����wހ�ܹ��QP=rAe~�֮�k��^̜��fM��oo���Ƒ�8��n7�,��;n���nBaY5d_Y���g�r��a֭]��^؆'~�"wa����@�[�w�������
�<�*��ES���%X<!��L��/�و��~8p�`lp�-�⓷�ČUw�W:���q��F9{}�S1oz��'�Á��5�s"���j��/>�+��?�V����-�HaH�r��O��?��|��SQ��.ȅu#�gY�4\���4|���pl�C&-�׋��u5�,�c"�mI��
�/�(ނ8�#��5"�8p0�p�\�����W^���W�a��4\������|���Gp�رs�gȤu��WុnG`����*�ކ������yo/8p0��:u*>q�JLXr'dO`T��x-x��;���w`��@C"����y�r��\	���h�~�J��rinG{[8p0����`�����c4(���WM�;�f`�;Cw�ț�h���U�0m�DȣLX��W��7��c�y8=�#�T��tn�j�B��j�\<x�e���9�Lޤ�p�"\=c�)��|���
����uk�r�`���݇����U:㼜�]�+��0��Z��ګC;6߆s�բ~��!,��	�Vw'N©S'�����ǜ���ƛ�\p^�[0q�σ��COOO���EZ��5X{�J�O�����n&��Z���
8y,[�U��o�I��-��~L�:=;�>./�*+)Ĕ*8�p���ʅS�����݁���9,�f阜�z�JL�܄]#MZ�PS[G�q����1{����>8p0r��7�U�cv~_Q��H|��29��$��2.�e�M�
�QZ6��%������t���*�CIi%פF��<�rxK0V(�z�L��&l�F�Kv��0�ϯ��Q�i y��h�*ʡ&�.�F�8�U8�����aј�_ryQ5i!
�Fp �āy�V��P�}+(}�����,���95f�2a��}C�1΋��Ę�D��g``�8p�`dAd��uv�ί&b�8�x��,B^�u�D+B�^1Q����N>yF�=�������HZ[;�T�� /�
�����Je:(�/�H/��r�5�����E$Fs�e�r�漟���zl�ck^���ı#0gٵ�����]{�~���ԁ�� i0�:��ā�18�@`��^�1y�VWW6lޅ�W�Fɔ+p>��ъ�_��6nކ>����w阼4����;Qܰ������x��Cػw8p0:h>q�=���L??I�h:[N⑟�l���MZG��{�b��w�z=F�Cs�lm<�.�x�q�[��W���dʨ�/Զ��z�;t��!�����'�x��K�஘��D�s6���ش8]tvt��7�b��i()�0�!{J�ǎ���<~n.C������0k�2T�υ$�(����~���sL��8����k[�p�l�R�Ѩ��4�P����&���ͩu�t�n�~��wo�����0��#��`�����uH�*8p0<�����$�jk�d�Bx˦�h�jl ͛���G����ι�֐I��H���K����;�l�ʬe���hw����ݟ<9�T��_��3|��kp�5W P���J����ċ��\�	�\qN�k__/~�����B|��^T�/��h"��x�x�E|㗍ؾ};8p06ؿo��]�a\�|�|r�}�5����v�[?z��������F���>�S���cݢ��T/���ϻ�D<D{�i��ܓx��wq���o:p�@�,�������]�%�̘R���eyOs[Qb��4c׮=xv�^���zn.��D@��dw�nw7�,��eWބy3�Q9a<R��Y)Ǩ��x�q�
6�tc��&���^ٰ1�$`8}=r����X��\�"\w�<��M���
�@eZ{6٭"]M���¾C�Lkj�3��@[��%��u�'��a�����1sJ-V�\��2?�Zv��)
Ƽ5HH>��s��oĖ�=�⢳J����Ď���w�0��C5�Ϟ�%�Va���twB�j���'��/�_�Z;�и� :::�p3�Qg�&R���wwٶϛ'|��������P������?�au����d;8/yV��??������ETV�]rh888�����
i9p����CZ8�����.(8�����
i9p����CZ8�����.(8�����
i9p����CZ8�����.(8����%I�PZZ�ų���n��:A�O�����ذ�]^Q~<�!-.!�������WTBq�q@K(zc�e7\���>��z�5�>s�i9pp	�ƫ�b]�{pŻS��o�ڊrtݹ���s�pHˁ�K��v;��wo��}nFf�݊'g��ѣG1ᐖ�
Q��z�v�p�a-��B!���*\�v�y��};q���Q�[R��>.Hj��\�Y�*�i>�&�����������:,[y%|���;�ی�S'��K����3�9�/��ӈo�����[V�p����g��o�\�?��!�$5dT�����;p�}��,�8X�d)��?�]�})�5g�Φ�� zzFo��_P���J��r�۩Zn��4�>�U�$�O�����ŎZbҗJ�@�0�!�_�X�>� /m:&�;Vf}
QP@_�_p5
�ʫP\\��MFy�M�����o��G�YU\u����W�e�"#�*`7�͟�1�b�f��͗�>0)J�����$5����?S8�� �$])���H���o�_��Sn���Z���+�|��}��|����?ï�!߇�e
���V��?|'k��J.�,	W #YI�a�$�"��*{Yo}&��d�Z�e_�$kc���ɖe���!.��?�������މ�f+���U���K�� U���dl:���f>z�ov�d����&-9�_MT��SۇA�d�,F\eK�n0IPt3Ș���FB���l=�d�ົ��9���R�	���G$i�I4�=��?*��X�	�f�RH��&��*|��Wa��ȴ%&���[$�Ώ}+y/'��ա��yn%��'�v#���J�MjW���
B �')���TEW"l�_a_ �������4o˾��LB*c�8_FF��� &m$�*��D�D[I�x��(\[��k�!|�+�púk1�~%���b<�ү���"�.ܨ��%iA��I{Ά�:T��y�>���P�Iy���\��u�rF8F&;�j�?݈��֔�*'�.A��N�nX��\����5������p¢m�EP����`������Ĺ"�@*I�u-׸�]丐�|-܄B!47��� n&as�U��iИ/|{�sMF�S�c}��7,�X��V5#q��p�*T>�������p��m��t����6�c�&-�	��F}CIEr�0G+)?��i�TM�������&��U��n��`z{�s����(��htK��Z�y��x�($ctvsw�-���NP���YI�vFf��N$$�9����}C#-Ք���"1��X�f̾k�k���AZȢ~��x�%��@R�o���?'��!9I+�v�<$��¿D��KNL���b�)(�&UB��Jz���.틓S���+n�۝�P�<��������S���mj�\Ts���3_W�>	��ζWE�}�\���w�3��(i�YƔ�j���黵�F#ط�Cم]�~Zƙ跡2"Տ��u��*�����G
f��x�iL(�@eL��B�9Ľh��A1\t;7ʓ>�ETqcUM%$	J�-�>�R�
�Sb��e	�@!#.7��E���	i�@��ٹ����_6����ӡ��Pۥ?goo�ޡ�c9��������� .Uۢ�S�ϣ*��J�R��|~*C�YI�*��g3�Nx$�rn�2|��a��{�:�f�W��N{�TekAx�È�|5�^č��۩����4�2�����o�n$�>�+�Z��C�X�$�n(����c���D.��7�HT�������� >@� F5�FU#.�ר�jH&Zi�B�&d0�A��!U������@3�3�fx��W�\�]��܋ؙ�=�;�����&�t�0��o&�mq��'���"�'_�P.aq�QI�\�>�6,M�/�_��=<��$���ߡ�\mE�q����N���<'�J�˂�TW�v��?�#7	�H�is�a&�q���\>��W�D�vw���fA�=�x�;�M����1a�ڳ���"��>�P[��eM�X
W��T�D�y�}�o��U�T|�_�e�e#O����@X���v����6�m�el?78�uq��/��5+��C����6	j��8��/�=+>�mĽ�*���~�,B
#[��K!ۗ�Nĵ���%A6�
4󌢭6�aja�<kS��̈́��?��� �t�L�a��=L4,d�en�5i+�=������B%T4Q��,E��.n�!�J�'z
�-l}ǋ�"P;&V�|�!����;��,Ĝ���M"����/܍@�o��2�j�V�����߭�R���^�͵��y���#���/��e �
��[W弬mHڒ|�L�;��F�b>-bU]�����¸��;/Ex�j+�>}$� <.�6/_� �c�b8���4���!��5�w���]�X�]w'-�K����sG�-�'{��s�7/�
���V��qΣ�� w�����XP�X�A7s'C�Z�'Z�P |DH����T���i�������p�@,R_�V��<�V#o��*���a\|��A�sb�@q��mR����˂j����I�#�U&S��-p�fwnS3;�Z��Y?g�V����q�LZ�CO�]���i��
bn{��W�i+�$�z�o7Ƈ,�9�\Tn<�o�A`��Y����H��Y�\N���Q/:��wJ�� �0�#�ڤ�wc���u��CIUT�Aᐍ��Z�\��Kʥ�9�μw�U���$���=��LZJ�4B;���%	W�t���g�F�cg�=Z��HM��j���G�Y­�n4-�J�o�j��$��&��I�D׹�@�����x�Nc�j6G(m�bK�j�f�� 6AX�&��n�ƥ����݈�<��h�p7"�A���þ�a)�������LZ9P�T�~FX���;�Yw(P9�h�E#ۢ�FY?� +���/��}Z������u���H]�+q�BWь�+{�UwBq�Җ�^�O�$�Q�3�i3��O vj����z$� ޹�i^�y�_6���$�P;S=�>4'8R��*��(WUK�� n�5TAs՞I=�>������f���5�0_���|H~�DV�s�C?���)�)���#1a_R9	�V�	P2�=')!�� k��6�Q^����`�8�51�H:
�j<��;�Ǣ3�.&4�2��i�\YV2���@^�I��*�eD8`ˀ�k4c	���s�W��x��D|���*N�c�z]�P���៥gr*!w!�b��'n)%�d�1���	$��1XA�x��9�E�� /�Ǆ���#4�Ej��A>�v��K_�˛���
�v>�L[?��(hܲ�G��8�ڛu�c�MFr�]����N<��n'�c�������ַ�b�`p �5�\U�Ȅ*�]���8D��@�������Q>�s>���L31_���� o�ھ�4�3���Dn�wv#f|~VW,�nt!=�(s�	`ņͻ-��"_В%!(�<����Z�* #8Rץ�t�\�]�[���}e~��?�������7�����G�G_�Ӽ�M�Z���6h�!O��<m�um}S��u8��P�6E��c����+�2��}z��tg��t�x�Q�ּ��[������#ze".mO(ꐈj<Ÿ�r0���R�I��7U���>�&�N�s�>Y�UI�;퇹e��:��HZ��]��Jɩ-r�"Qi��"5����#Wwi꠸q�mњ��Nm�#�/8j��l�fo��9��J����A5��W6�����XQ�ꥑ<pd����ʡ*yW��7�LMC���Z���X��2}��vϜ9w�v&��8���1N����/�R����:���=�ᨍ;rTͬ��+��e�iͬ�
�av����H �������AQ��Z[+����d٧j�K��.e�B�n���K��M�tJ#$S��s�ĕ�m����	47�0]�2k%U�<U�믻��I(�z�h�ͅR;�ζu�ʻ�p��!��������5z�f�=`ZjG�Ӎ��W�6}��~	ZN.���)�hs6��}�E����i�Z��Q ��j�G���V8qr�UDB1t�_�:�VW3K�H8��t��@3�3��Iղ����z���W���k��e�)/��������.N���<���8r�=�K��o<܅���l�kKbV�~[�f}��O&�E�]�+)�C���_�9���t楼�*t�<����*'�&�˩�J.O{!��X��%\�^*�i�ڪ��d�yf֗�^
i$0	xQ��P4+{�%�;�w��-�o�DJ��e�i
� R�R����( �}H�߰�*��盗˃Q��P
���h�Sy\%��,rf���Q�@M�CK7��<��	1,�)ғi|}?S��#_1{����.1P�\�j�K��J��wN!�xc˩�e��Z�;�W��5!���9��zx�܁�YIK_A�޳��C��$}>�>E���CJ��</���lX�p��7ߤ�c9�)*"	�_��狋�Ja�N�i�M��*��l3���z6��k�NW	M�x�άW�[�nfy9�p�d���VjL�޷��q��Kh���(����D���B�0K�5Ӽb	4��TE}���ZjQC��)�
h?�-L��,�.C�@DE4�](;��s����S�cw���6^Ġb2�
�'E.��S�*�j�� ��$���=%Kf*T$�P�
�6����U�<�f�����Uad�R,e��0y���7`޴
L�T� #�=G�p`�>;֤��3~PT�tk��e�HX��XB���� �g��3�;�w�([�K��x��&z�6���w�'NQ"N)�`����Dfb[��Tgt��PWW�o��x�+�������q��!�����R�g�q���:go���ꊞ�G��n�	_xp-�[��'z�8�C�@�7�GVc��8p`�F~��N�L��R�d�h���]\�j��%���F�p�{�e�	��UH�3
o�(<��=�����00$E���D#�x�i=X�om��)iK��rE¤�ou�������wޅ�_S����CG�!L�XY����������/7�/S닧{��=f1�g&-��fQռ`�ݬ���'n_��gu���w�Zҵ_X^��W�ODq��Q�TL��@n���p�Q�UN�)��HE,	�GUxȩWs�S,Ҟ����]�ۗ�Q���)PjP^���T��L��@h�#/d8�5�`W㳳VO�Nt�e�r��:������A�pT�=�����}�bÒ,�[V��K�E$�p��#�<�����>qn�t޾)c��ZQ��>�jnX�i|��ػ�7�R��|�:#iqw�e�>��M��n���Y;v%��x7>�QF\O�����ԏ��4ʙL͝K%=S��{��8�����$�N���7���c�&���x��a�!<��۶�����^�y����ػ�/��m7�:��[l���+���x���
�Q�j��v�P5��t�����e� �Ve=�a�<�ᵸa����^W�;f��[���N��w v5��YNR��Ղ���WO<o�$,�x*��o���2(����lA��K\�rǻ���]��>��}���$[?YK�^gM�W�z�*�x髖�F7�e����G�1D:{��޾.U�u"�tu����BD�`��� �p8���.��j����U�	Ko�l㒡�7^6��v3�2k�����7��<s)!��o��.%�է��?���[?Ҏȥ���IZz��ǃ�n�BA�Mc�w�(X�es����i��7���܏�8׷�W�Ƌ/��I[�UU�"x:¾ K 4o��)��*�W&U-�Z���j�� 8n�	R�'����b���R%+	��}�,��FX����`�_؎)���mz����M ъk�����ؿo���\���k��Z�*7��E�l�e���(�{�8ք��3�v���l�(�4�x�r�RJ���L�mW<w<�p��
�$\,***0}R;��ź0cZjJ$\6����v�D�8HGm�{�k��R_�25����b\�p
��s?��+w�� �FI��Tm�6C�*��T6Am3&Ua��" (��믄o�'ӎ�;�.��w"v�U����e�X4G#����<b�O�@��� C��Og��2H�5涪2O/_] �RauFU5?.���4��%-��e�K��b>I4�Vuu����a�o+#4�F������n�ml_��i倣6�_�^4~`1�.��%}����e�Ur�m�p<����{8~��f/JVM�ϲ�n�J�CX0{�Q����g�Ր�%��_�Wiyb�X�p~9�T��%-�l���h��V��uH�Bȁ$�ڇ$�$�E���]*�+j�2�2b�~SN$�8o�\_��o��VP��������H]���.+�۳<��
�b�� mF����׾��I�u�_U�����S��缪��<k{�g��\\\��"{��%�a�[�H�R1:���b�M��uUNب�Zh������_���K,�Z��\9��=u+ٻBūsW#���p�s0d8���@�A��p;"�,�'��m7i-kfHB3�ug�{�[U�l��H�b���$r��y�����0�x{#S��gl�ƂP�<�2�	Ѩ~AVY֌���Z��+*Lk9�UC'Oձ��6�8\��5���]L�_�G��Kg��\�H^��!��P�t�>(Eˡx�K8%]�j��V;����(/q�Eҋ\��M��n$�epǻٜD�s�\�J�8�oŁ�v93����n��k?���������J�g�u���VDO�5$$3���j���Up���3@x�jgT���Qp�^��ӫ7g��H���BZ�d���k����sE�������=j�����亟��Q+c�GO��k���5�ؙ��z\ER�*������`�R�kj�P�#��^��9rg_FM���E�1��C(���᩿��:.�+f�0���!�����Z��m��F�S�OH�b�3�%�"'�M̿��ޅ�W�u0rp�Ʊ��L������dn�0-���_Gk^��2�B�`�I�t���gj+E��ׄ��GP��l�i�(�.ԉ����{T���T�_xR�5���S=$GPU����_���ĭh�"ތ��l �ʗ�X %Ԏ��י�h��*lj.��ݻ��R��.VV�G7���vx�0':�-H�1��,�k.$��K:`�|�Q� ���x'Q�*}7�v�<�3�����*���+"D�J{{;�z���S�ro�؉? v�5������.D��P[���8���ы�Z/C�Ǖ%5�lH4zx��ai v�R�'vpfVc���U�v�"�����ӟh^�Z����6n�㨉���?�o�YW�e^ʛ.Ҽ����p˔xbf=8�wp?��#@A=�.�q���a�$����*=���<��G}����BN�S�oQ�Z>;"�t�b�%l�ӄ��܊����?��H��L�S[\x����ј���,�i\���R�^��o��	���k05�Z���������-�j��o뚅��<Q����Iʖ,�
��(Bx�"'.��ٸֿ�u5w�#+��9���S	W��Ȁ��l	8R��1�<��j�bFT���oF��;?��rZ��d��3�xx{�NT�� �udP�g��P(��}��h�n>{�Pҹ��)��7P������[Z<�5cD�?~:d��"�'!��ٓ*��l�ֈo�P[���)F��p/χ�+��[��ߊ-[^�:R���`��ՅCi�������R���Gp�P#�~��Sضk1����'M`�Ro�ވ�%`zo��K%`z4�ػ��~������N�ꦙ�IxsC�>�--�c@�Lw��gtҗC��VOV��hR;3?��"��^z;��g>v3�u�$v�E�=A��Bs�_�{�챌��?沞"#���Q�KT�ѽ�Ei/��w6�f7U�d�@���{Ǐ}�W��$������?Ĥ�<��9\dC3|�D~n�(|�d���6"3
��\��N766�Q۷d�J�J&���0�`$�H^�L��x�������
k��$�7��t$�OMcM?c_\�"�O�д�����J����45�����y�ښZ��OEwwζDoϫ\*3Ϧ��i��5:���Ihj�N�F\AA2�;Bgg'�@���C��� �GKA#i.~A���a��O�VE%".�e����\\�+�P|��I5�p�]��!oک��g̕��40iS��0���d��J�o�ĥ�#�����������W	1�%dG�B웈��2z�-^iG�ɒ�T���yV�Bm2�p#���H�j�^�P���^�y�Ք|�z�C���pt�H]�����K�,Yn�x���d�>���Ǻ�8�Z2��V����<y��y���n��)y_q^��/���dw�%!NLy���+�Ui:+��*��YKŐT�	vNݟ+�o\��}������uk�n�4�
ɶJ����'.��ܛ��ڵd9����ù<����ے��X1�u,�Q�[��i�^4!���EX��t4½-x�����x}Ah>����s��9I�P���^�������PE�s��U��nV�.?󻉬."�BTs8��4�����M��j%�t;}����`Qn@C�?�Ĵ_'�WC������_��/􆖋�Ks�L��kg��i9�������6�8_���:0Һi�t{�t�uR7���*�5wO��'߆G{�BLɉ��4��S哚��@AO�	����a?��RZϙ���@v�rAP]�4ou�ų�r��ݝ@���S�w^�,a�4o�����q����e�'�}�"����(��t�|������Ÿ[���`��:\��]��	�qݝ�9#-3('Y�1�ְ��0lYlU��K�"M��؏�ڑ�ݜtv5+a�'seW���$)n��)|51��*]��^masH)��Rh�vM�O���~��E�L�����ػ)c�c3�$b�� �g��s�֑��[I1Ss}��I�#��&�(|��#3ּ��1�/�����%�QZ�����z��FTW��3�����K=��"O�1�s�]���hA(����q��yx��tm�w0��7m+ʽpqs�hKc�k�c+�<i�G�M_�ύ�J2���J��}P�^�y(�،v��:he%�ݢݘ�i=���q�$&�lOiR�쩺�[�meP��i�UB+��Mۘyt���v%��ğ�V��)-�m���v��9<��,'>X����T�L1���T�}�b)j�u5��d�g)���L��îޘ�|��/�&MM��`-�a�/#�cK�ܨ��UX���q6�d�d�$�FY�Ǩ`��x�&w��9�<�]QNDZ�0#Į�(�+��'R#R�y���È�H���o��H��'�NFt���m�:*�T2Bҷ�X:���a�����o ����Mc�z��د��G䜌>6:�ߗ��D�7�H���3̮ǭ�����q�cmlt�m�Q�WoG����QŮ����7�vgmR��\����E����)��j�:R��4-��i�Q��ff!�����n�D���n$� 4�X�x	�0���y���9]��2#���`i�ˇ�0:��d�X
�L6�:�b*�PL�*-�ȉ&1I5$�(�5���&|kG&�{�M����(�n��4AI���?���H���~��Z�IRPE� <"�nF0D���&1���v?#�0���=F1{_����ȁ������q}�CR:�g��g�)�3���!@ۋb\�dDJd�܎����(�y��5����v�Ml1Ϥro ��"�3z�e�*_���=���Wk�t�W����^12�iAMkd�,�G������=�2P��|�.�����|Z"@�* /�jauÝA2څ��7�3_i�4-�<FϒK=1�dMX"����i�"I ���)>&UXUA�d��I&� $���BoC�H�d%2V�P���ɂ���*�vZ�:��&I#^�dF�{�� B�t�=�f�A!��U��s�8��Z�"��&7س�F4����#���e��U���N:�:�XH��%��n���Bs�@�?Tܮ���dUd��dm2P���ٳ����|�Ş��Q�ن�ѹm�"�dn�������M_�L����.����KZ�z}L(��es�x�\6�
�L{/�xk3�[�ߟ$�Rܠ�@Hp���ϛE7M֗V�ָ�4ܬ�q���O����kK��#�BG�er�\H�	/[&Mf�<yCS&�d��xs���9��%U����/�n�r2�%�&��ٰ��E��&��t$m�t�]*b�5�~;9�>I��Z2��x�+Ɗ���.!]�r��=�� �v"$��i<��iۑ-Q�C*UPn����r��؝������	�f\�)�$ h�E��")�l�o��i�����ʰp�lT&p��+�v�����gp�T��N�*i��\��� ij�b\�^Hu��ɸmU-�_����v��,Jؓ��^4�F����4��d%'S�э�Bi�i�P��2��g�Fhѻ����X9}����p#ރ�'�wl��G4�uC�����/4Y=EC_8 �!5�4�j���qM���D0tnR���ܹRD:$�4r���?��ҵ��1� L#��ںe�D�$]��s�-�`���E�O<1tB	���U�f�ot��%/��h��g�9�(#�8��	W���U���|d�i3R�U�9mI"JZu+".��YXD*���)a�X���[��"(�;���j��"^{��\��~�;w@7�q��!��eFx���l�(+�_~pV�4��`���L�=�_�Lwc��E�Y�<��zK���	7A�)A��%����l:~
���0֭���J!2WU�a.��}�N��e����X��Ξ78'���k��4�iB�j#���OR�p|I�M��N�]#8(�/
d��8i��OD:��)�&+��n�J����&���#	��V7Ip�q�/��Q�i�� A�{<��m�@�1"���8ﻤ(3i�b@k{�Kz�^��`��k�li��Ҧ-��H�L���غ�(v�;�?�6#��#��2���d��W��f�a����+��{&c�����#=U�/�ހ���1�#���x�oZb��nّC=�:�Fw�����?��cv����7N�S�q����7_���b����.�F�ɓ�r�*D��}-m�x��x
��6Z���θ	�&�HH�קX.�V���{�-"&THˎ�.�V�
]��԰p����������އ~,١��h��k�'i��j� �~�@���L�Jg��G��n��'&��I
����5��'�pN+��@�ʊ��$���HMv����������ǰw�N�����AܰEiy�O��*r�^����d]V4U� F��I��˗/��~x&Z�$%˱�G咟�����k��{U8{���"u� �L�
_v��|�,+�if$&�LX���!TA�;��[��Z����3��Ͽ~���9�/*3�%�t������H�����T�$u͚��������|�|>���W���D��YY��FE�Vz�)L��J��'�~����g�ф�JT4��<�mW�	�V'IV�1>Ĉ�Ț�m(lJ�t�t��<�[���:���B��x�"I"�,O]$b�{E�������p�oD`؅��}�e�F\�UUԫc�������ni9�o��jy�yO�Z�9��%؂��'��ŷM����������x�V�I`�#�B��L'M�-�"(�5�,�#�k y��e��E�w��濃��<��l��3�a�vS���Թ��4I²���_��� �.>-��h�����:�����ؙH���������G 5�[h��t��l,d#�.�כ�î$��0d�L5�UD#pRQu?7+H"si�.�vg�Mt��E2#��$_+���*�Iv�5^a��ޫV��٨t�(	�ݞ$TE�a��U/2ͥ�j�zN��z!N@��?�E[uP�5��@���<M;����֋�����!u�fF�$�z|��yP�5�x=c���wZ>˾���P�.��9[v 4�;�&�V:d�a��A�v����V�L��u���x�=�����Cx�H5w�?�8�9��H�Jv-��C
&i��>�V i�k0,���>Ic܃]BΕ8Z�$�7��}.��9D�Kv�J�.D�q����Ɣ�����:��H�&�,*K�9g��L �2z0��O�v"��ma���^�I}UV-h�Lϩ��������=�;v���!8��%���Z�O�q����3$F�3���H!���p%�T�&	{px&߄��)D��o+�ۊ{�� ��������ȘV�&�+aز|�?���\4ra��	��ϕ�P->$�v/�L�.��~���(�����m�U�h.���q�L{���}���=��ȉ�$ ���R��H�!�ӑ�3���&<�I����`	!�䚠DD��K�;|��Dd�'I�k��ѹ�u��H%II'
zȐ���mEi��HJ�����x�c�Zx�A>b��JF�d�������=�i��C]��(�{���������h�܂n,���T��{���i�[�Px��"d�K���^�[�~]��Lc�E�%_#�˙���{�d7��t�"������_�)��ϛ�$�F�����.���g���2�)�b�����LI��;֢��ٔ���b�]ň�c5MYN}j	I��I���{l�^�$������2$H��j��O*'�<���)T�tkg؋�LDN	͑�����M��^g�T��T��O�\,�{b��W��L��t(���V
u5�e��{�⒠���������m�_��P�Rb�7�pW�Q�!=�x'�{����ޡ���E������ic7v��F��r���+ދ�"�)n�[�?e�4P1#�,v*_%۰̝s�7��������%���~�yF�H��?�RW�h��Dv�IO�,$�������E�Bn	��i��IG��섪KF�<�D����/I2]1>��:tu�Mw��1��x��2�˂����\A��j:�D�$��T�ƈ@��m�N΂��dE1�%ڪ ]��s�A��>�!C�u��G|��)���ъ�+�o�Q�nr3�Z�i�q�lX��.MI���[�5K�9����s!ż�8ݙ�������7�;�ƌ�b�R����`���Vf@M�M�F��REU�<�ҫ�U$����jK�
�-�M�L���"HR	����м�iE�8i�T��8:�ȃ�����lZ4V���;IFh݃�
�u����J'Y�F�ib�M�@+�B���q4�霺;IltO�*2I?�^C*tiR)�%��ۑ��MU�vD���tu�8Y��H}ɖ�t�پ3:F�G�ǒ�	����V�JV�}�J�^aZ�@�o��L/�`����aڨ�P��em>����3C{�r�[VDmCv��w�@��e��l��bǞG��z��73�Ʈ�S�����C�	�x�M�3��^��r�4�n��JN���7�b,���+�s��'�fɆ�a�	�RN��ky�e���Աf[Hז�:�="�K>O���VӝO�0n�vR���9vY"]Y�d
@��G)�/"u�����!�8p�/���~���Z
O�*[;�I�J�	D��������7'�9'��F�)�A�=ۀ�	eL_����⠫j!7����06M���}��	������d�喥��x�Yi�탴�����]m8��Szs���*�6���2���ĚܲBm�'���)�^}Z�qi!?����{�+0m���A��n���ײ��k�q�?����3!�Ǝ����ί��F��x]A��U��}�I���LzF�d�i��/!52iK8,��6p{����p�+�eY�FZɃO��d�2�gO籏)='��$ڙn��`<�<8��0:����!R��U|�ɱ���`	�x�-�E�K$�TEQE*��j�p�ct�� S�z� V��2LR6�}J�Dz�"z�EH.!�*�mB��p:6�R�ݘ�S��ܤE/��U��`�	�]���6�H���<�B��K����=���]�'^p5��f���l�F�'/��O-��3\��w�Z[����[ቜB.-�r��q��B�#�!Kq$$��I@E�]��>����`�)0R�S�Z�̖��KVჇ�����ėn��E�"��Cmi��2�����<tC!+�U�!�W����[����s���fb'���uъ�L�Z�؏�޴>̢��a	�Iw]�Njb篞|J�����;�ѪD�{"j"L==�˫����Ӷ���8�`(ƃ�]�P���i�(U�
.��x$�]g����Y��,xA���a;	Q\�����以����z&H]�[L��Qx�8AG�U���{�
�� 6������ˇ���QxŝD��0��L	 ؏���`т�X3w!jK]���1�ġ�h9�wq�L��+�D�i��LE�ٸ�}&=��zly��� ���s]�j�$<��-�FM��T[����wl�s����?��נ��Y���A�b��;���p��ʞ��t"��:�u(�*�ٽX���܌�;K�hF��j5ʘ�PU��S��^�nlĎG�٥2
�R]�2W�j<T0�]LD#���Dً��g�뭍>�鮋��#�8cz�W��2)�E�CT�V\EHo�J�-��+Y���7�Um��+��ő���&˃��#i��%�w��F�'�,�ɕ���������� �'�l�4	Q��%Ex{G/��=�UP=�g��g$��Ӊ�k',��n����
�ڥ�%R:_!��(�J���ԘB���z����I���2��2�0�WFw��A�*J�^��7XG�9������8�����/��L.:�� ��J�D�HBT���$��d��\��H�u)A�>�ŉ��9��C�@�$F.Nt2'.=!���Si�}di⭔�q�;��%Eb%sʤ3�\0��1�IFg;����p������xDq���u��������W�y�EabR�N�mC_�V]��Sӈ�Fp��|2$��6�?a�IGv��Vo���Z��ڲ�M�tJ�?�l\\,�&y�=�[W�Wz��\~!J�}����~�Z\1�� $OY�"�����˿�dc�r�`|��%���[�¹*�zP4S��{�6�#�t݆������jI�15��L�4k8�]���,�uek(����V�aҕK+/�y�e�����[N���f�d�0�A��^X��ǘ�a��t~��0死z5>�h��E<0 ��b������ct��RQZ�C]U���Nc��EM���ԏI�A|�+��W��]��EUM�.�!s	K� 俢'lYP�E*LB2�Di�峮2����+��R"f霱7��d^jH��-[!2 B�ꤞ\P��^<��RR�X߫�q�T�79�IF�`Wc}T�ĝ+�P5N����X�3)\Oh�m�;ց*�d���U7MbK���2T�-�W"�Ef$��F2��t-��I�>X��dʹ��q�)�,f��R����Q\�j���P-2_,�d�7�}���Q�t�J��������E�?��4m�y�'������z�5�mQEj����%\�S����5Ӊ"f�W�*b>����e�D�����'�	�m�ZUh�Q���Lr, w�P#���(�jeZɐ��.bf��	a��H9�
�=<��CZ�?�± t&ko�
D���"�͂s�ymZ��3���C���[ӥ��}�,~Z��|2Om�� ��+e�Z~������ۤT8�ZJ���Oӥ�#��a�J������(����\L �+���Hٔ�w��H��U��|��9N���.l�Y��f�ʑ�L.髍a�@	1$E%8����NXzE٢�b��Ԣ���� Z[[E[�eb�%k���K5�b\���L��Vg1݅���Y�Dh�-C��<lZ\@ �*�ɦ	S��W�{��f����(r9��{	C���ZY�3�**+7���ZZ��n����,.
�� ���<�
�ˬ][[�o�K'FQ*���0��`)z1gCex���x���ЫG����2J˛������ٸ���6.�������A�����f��op��#��\8�C+�\�E��Q:���?m���O�%�(� .Ս��u)G���J������&L�=�\�9�'Q��� 曀~�w��TW�7�[�6,v��<$�Z(�)k�&��:w�\|��U�����_Q�+��Jd\��{��;��ȯ�G$�޶j"n���[tq	�$.nG#��V�|�����Ǐ��G���O�?��U�M��'��E
��'G�D��F1	&(��w��E/���KW<��Y�&�NR����]��r|�#�Pѷ�������.[����|��Æ��%.Ii�k��*�SV4�?w��b��F<M{�Ki5�O����������pXT�����=Us��4b���%�	��Dþ%��x���/�ګ/g�Y�o��ɓq��^��VBl0�j�t�`$p>|��m�3�r�_}�*4�t��W)o��P;��ۈp$jVI��S��=�u���t�����?x>�f���Sډ^��V����ܶ ե���_C,KSn�e��̞3��E��n5W�p�,g�]ʫ�RJU5��w��'p�R�f%�]�67��O�Q3��6.=ɽL��%.q�yT���l�J���`��kol�.�-Y�%e�x��F'`��E�=���e���ĩ��B�Q��2��[��mM���5W�#���c��T������0^8�s�SVSBy� >q�*�w]�om�����s���������]�E;�O�8:����W�B��P�2��Ѧ�=�;ޤ``7>r�b�?6�i0��h�`>�"¯����%.�q���ː��98:�-�K�����9|�N�?�>���&َ�r&mwyy9n�|
ʔ��>�h2
V}�W��<E�=G��=&�4sͪ6ވ?��>������$-U�r�l�rL���5��	0r)��[p[ʈIT馠�>�D�$�D��̟Z�HK܌t�'L?.YH\��=���Z�<|H���V��*�<lToq���MI�_BBq����E.��{������<bJ�KB<��"�*#	�:h��0؇G�HviL�*f��I�p��0\=���^���\Pe��xAf� OB���`�XR&������o�=�N��SfVҲ^BEi��7!�����V2���G��R�ƚ?��l*Dp`@�L���l�oHw\�TT�J������ŋpżbT�r{XY�4�ה��.b_�i�����L��8��]+sKf�bɬZq�{:�r�DT|�Z�9�*ƶ�]xe��F��e��ic��w����U���l�z���
W�D��	����I�ϧ�O������!i�ьI��{[��w͊�G���01qOr/+QT�{���8ie����V�UkG��Ü9s��O��$���������[�Zo�{�M�p��B��)���m���iB�O�A�N��l�f�t��߃��z*��4ye�!Kj�U����{.Q�N���Sw9���'U�./����ym��XW���"�r���NKKk2~m7��H���Bs�Dc����nY�)���}�����­�28pp"�.G�?��V^U�@kэ�3��o-a2��vL�1um�ܜ?�A���>{C'���
�y��WV��Tc�T�QM��O�m�%�v�Q�����a�(��;kOM�+'Oq���y<5Nљ��v�+3�pc�<���?�h�M���,�A-�]osy�����gI8�55��cL���'�<����T^��=�2�����̋jjn���B�@�#G���zi�#�m�A��t]5���M���K�V�(�y���\F�K��f�x�%˄���[+Τ���@�PS�g�3CLMC��2I��x7c�8�Ǡ����>&2��m�=U�ٶ�CE�R�F͎�jG{ѝ(a��Bx�����T�qѓ���9�H����
c�P�ͻ���4�[>��*驔�:���@���4P�1;X�K�9��q(�1�N��Ѫ,�$��_����T@��R��N�������0ӂ^x�y�C�WEs��<W�"�8q��b⤩�����FZ�3�X�|9S��"r��}ք`]q�odRw��mR�R+7�rՎYK.V`��d²=������_2�����EZu���k��b��"dD��B[<����Z�/��4�϶b��B4L(�Oc�����Q��f��p%��;=��'��1O���CGG;�<��δ���C�Q�Ƀ�|�?Q�g��Sz��J�!��@�n���w_�Ђ�u�6���A�B��
h��9��C0���eU1���i��L5�	.*�#v	#)���i���&۳����i��x�ŷ0�kpY�{�D����G�)��ț�����d�#`�w��XjTs�t�U�_���[���=���ys{��b��O��Z:V)��B��4xs�\��M(����q0�����9���I��`���o�[O���V���G�*Z�����t��F�	MG��[�)��������l��y*��s~��1�ut[��lYHK��4���h�?�7]���:xA���q� ~�z�����Ϋg:M&/�X�i^6�i�m��:q��
4T/�=y�P�5��6�'����h�[:p�x�.s�L]�g�8��W���'�o��T�Fm�9Δ-D<��P3e����_Fq��qüy��ޓ\���k�|c�|�%��je���×��q<l�K[
�p�����{ϼ��7ބ��WaŒ��q����xy���q��GH�%V��!k���Y���ĦX�i�Vc�n�7�����h�.��<�5�y����ވ�~�	�vp"=���������7?��{w�?��0�'Q���F'	�&娒�c���'���N�:��}�)�4i2���
�-���
:���BlݺMMGY��qخv��i�aq51�3.(|��%ϓ��ϧ?��g�D>�=T���(��o���TL�Y+}�ݗ)�Rvt<�0�+t�Fz�!���o^x�<:�ݲ>N�l�g��p�A�v;V��O?̼�K����+׊Zx̬��v]�Rͨ..i��������V�R8�x�RU�4�rw�|ہ��j�ے����1
����r5����s�\ϺzH�<IK�'HʭU�Vj��Hto�gj���R���%�7C�'���#��Ă����O�Nh;�ꕋ1����]��٨�*��5�FM����Cwhs�`�`Bu1*J��m�XfN���������w�� )5��0�S�X��|�-S��yŐ��N*=��ٜ��1ē[��(.��X�H�s��Ո'��&��,��C�®�Cꤖ�|���w!Q����
�K�u\��8%�����s,/x�X+ߦ��'�/��u�o���N���q6����e�𙻗%L��E���*Q�U��y�M��_����X�7�a=�=5��,�R��BI�*�^�SS��fw��O�pK��2bLm3U7I��\$�/j�p� u�l`�R̡������F�en�E.y#�}:��Ӻ���·��ck�[���dä�C5����q%�ቶۯ�nE˽��[?x)�2��4�"S�S���F�����������Q�K?=�XK,����`T�՞�A��Lh	�4R����9�� j�;�^_�1���[�����Ō6}t�LD�p��.�F�d5���O�vQ��˗�@Z�᫐�ﴩi4���L�V����(�_�RB,�ʇiR���]�0�e�����Ƶ�G��u��>��H3��1���>qvw�7���:J�2�G���ld<\8�j�t|�; �x���c+��a/�j)j���`W뤬�iR}��.�.�f�TuQ߮�	da5Y��L�y�en�3O�y��]�>����y5!s�
��q������������̫�	�� �N�Q��dU[�$�rwbg'k'�d�������Η����]�$[�eu�eR")�Mb�щ�:�m�W@QI��#@L�3w����s��C���@�lɣ��( �R��M��
�(�᜻H��c�n��B�s>?x8�*<Sb�?�{k�`�5,m��E��b ��P�O�;;����3��f�1Z�f�c�uvME��`�ŻvU��dr�"�CQ.)�٧e�ڋxJ�s���_S�Z�5<sޱ��C[
-k�V�.uu����&Mf��hD��=�9oӔ��O���G��4
�&�� .V��CP�K7Y��^)��F"v} �T]�%����AX����R��B�0" �F�'NM��+�A���̙3�UU�<��-�Ip�����$x���J�8� 4���N��t,
a�U���}�aQ�9�{�̀&���800�w��/����l!�c�b��n�x�t��KT�& ����d���}:�V�XY�lW���]���VQ��N�;�ע.iD��4���$�L~��a�+���!٩i�\�ܟ�C��(��7���z�<�m!�9�i���uF�{���1>>����#;"��д$Ǭ�,B8`ݵ�Z|z]�ӿE`���*;�k�5�\��KV���N������t=7W�L49)*�*j"�5�D�1\ֺ�7nFM���z��g�#�M#�IA.�K�=fQ��^I�wt<������銦(F ����2e=5X�m�6"3��0p�EM� ���hU�}p=n�ه�xR�NW+��wk9p�W��W��ȓ�100 ��V�bN�V���%�[?��F|z����fO(�[&���e�X�z'��w�g�!���ܠ����&!���M��50H���~�<�k��hHa���-Ŋe1<����}�s=�(JQ.Wٶ�N�t���nƑ���mlY'����Ο?�s����6�d��_�̇qgӛ%;�K�U��9c��K��������m���Cj�q�d?��λ�wD�ڷ�uar�,oR�H��#�M4��B�-|����&�H:!NjeC��"�1_ǳm�Y}DZܔ��:��3p�m���P�+F�F��)t����gز{�.�O8G1V�q�}֋#:�����mu��r�dJ	&H���"%4�T�����q�m!^~���$��hfJ�xX�����q��7�|���v�����	�Z��Mx��H�z
��f!���l��g�؉3<�=g%oڎj�����������(Eyw�])tA_{V#T�7mǎӲ<Z0+Y�l/5���l�sʔ��gu9"r�� VYp�->�(3��gݍ��oC���觢�#���+��Z�X,6���;{hF�Ϟ=�6�R� ��_E�f�k�d"��ѺR��f���a�"�9ۉT2��%2F"�R�K�I�A'�ף���h)ZZf��,�L�	ӝ��aQ._�$�ti�=�$kc�#���%K $�hk;�D�T�������J4�vBV�yh�����@)kt�����6t���=���o�SO=9!T�S؂��SY4{2�`3��n� ,�gށt��r�K�h>�]	����)��>�Ӓ(Q� �d��F��Onr�l����	'��(E�������V��)��̚0V<X�"%�fl�7���+�t� ��}� U���W�,�F�B�����@M�ݗYx�g���|Y���G@�HLf�|ZQ�첃�O�[�s9R��-�x�U������r��7mGw���MMs���qϢʆ�XW�B�Z���2�Qá���.JQ.)!�bCm���@��tPFH�G�N����l��0~���^\/�MF��X�,�P��К�t�`	��9��Jp����h`�U�-�HA��=1���D�b$�g@�fkW�#��ی}ӑ��8�ɳ��(JQ.u����E::�Hqw�-0qݒ��G���?ʝP�	��i�\:>�&Jz�O��544UӘag�F����Rْu���G홼��Q$�ܖ^�w�?U3�R jd&+��y�]���R���y�Nh�Y -<��e������U�䠦1�����=M��!�t�V���LT򀖭���eH��N�g˩�O 4��l�<�4.&F�����������ָ�j<y%�G��qV�(E����_u� ZI������0��|�������g!06��Sg_F��j��z���o~˵�{�1LT�<�T��Ǝ7p��{�*ey���!���W�f�O:XG��0�F�鞝H��g��T��&E`H<s 8^�a.jN��.D˝�fgC �r%�H��Eq(Uܵb�C8�8H�����i��'qbd)<�R�ۃ��o ��/.���zb�sa$mM�l������2
�m�5%J%#��ߏ'_�Ǭ^��!N��:�������D�I@=�&��C�c�:ǁ�	2f�́sd��d3���l��|�44����FQ����(E�%P���!B�	��4f<�_ ��]+l&�����Տ�k�P��hx����]iꮲ���@���MZ�O����IV�g���X�z��ż��K��^�?\3!��&��B��d�MF������"T��7s�<���*P��;1K�co"�8>!��w>�(�G�h����I?�e�k=��T{߰����,��5���L��x��-h��1���Yt�Z���'�R�=�Waׁ�X�E�'NK��:�(uq<�'7�D��;qS��.Ϣ���:ۏ����bh��#
a��%v�ծ�]Zֳ/m��K�C������f�:L���R��I
����|k�0#|�3��7�m��yh�/���:E�{&��b�!�!�?�߾�}��#���*�$�e�����;������	��`�x2/`JNj])���3r>JC�cF������,��;_�g��C�����<�<O���^nO���c8f�����b㰠]ʙ�k��y����_��,hnĤJ�A?ej��S�8��rl���J#z�R.�R��s=#��V;�~W,�����ؽ����w���C�{��lj��cS��5Nr!��Ԑ$<���Y�k߈Z� ��KnhG��5t����06��3��m�ٹ�o��A��R�� ʺ�r�,�];108���&���Bl<�C'F�3D�"R^y�F���{�a(aǧD�B

��2/.�j���mg�Yۖ,]�d�?�іb�tQ�ٺ��q�׿� �:��>�[6,R>g��)NMc�5u�����X?��k���F��D1�1D0#-���`���=�&�S�f窳x�J�9�J�G�1 ���N��ބw��	��o]T�����9�̈́Z��r�k^�K_�--^,��'����3�����?v<�A2"&&9��h�T���E��&ċV��D:ӎd^��פs����LS����1Y�'ʊv��r.����l92��%��Pd��#;�����{řâ\�B�i�iH��W����`Rw���.ߒ�H�_mQ7��	y���+��
-�����s򶅁Y>-���Nè���5
yh�X����}l���DT�aj�,�+�kR����4ÃY��b2���>!�����M+����D}��m)G�C�X�^S~��~�L,ݠ(E�Td���n��]�@�ӄ�>p#{7�#�j�����X�� !y�̅jB�quk��;���1�?�*eJA�!�9I���3缻��'8�04�l*1-�����~v�����9'��dS�\�:�P+f��ff,;oi)��y�{���^�y�ZE�leVc�i��0M%!�U:�%K{�g�4�,�ǿV���[h ��x_ �Ą��&��ޭyڊ�� �
�-Dui������`j`N�e�ua�D@�$h��!,��j=��#h������ 9��Z��RN.R�'+JQ.��~-���ď!���O���k�ТKN�V��O�S�;'w�����Y,-cz��@�Kl�����/ǻa���	�Dde�"��9i���6��E����d���2�,������s$�W@�JQ���l&
�b�CQ.�n���H�ގT�B�G�y|�}X�p!�MS�x(���3y0�{<!jI��{�V����_͆��_��jVr�iX $����"b�l��,���8�g�,LE�u$��c���:.1��jX�?�ύJ8Fo�ip&#����b�֢\R�GS%�����R	',�b~�s�D����m��/eY�b�.Z�]�]��M°��r��ʧ��KO��241���7�+�
Q%�eZ�����>z�ZE�l$/pQ.x]E~��*$� j��.�Ж�Q�,[���-�2Ț)d�E�i��Cg0�T�)���VP��:L2��J�5$��N`�;eXNw�Ч}0��ܼd�r{ueom �EZ��\A�aˑۈ�*b_����V���y/k�u<��ñ&30<��Ş�W�l�mZ���+T�!D+��q��!S.�0���U[S���-h�\%��
D�Y��'{��ۇ1J�L��E�0_�3��GK���k���L�ә��O�/h���T7B�3@�\LT�����7R��A,T/!0�"�y��.�C��%g
ࢃ��D),���~#!c֬f4M*Ŵ�;.��N��F���'N@g
��
��}\�������Xv9�V�ǺV`��4<�@z���>��˱`~��[���$mB�in�LV�XS�ދ1�[�/�7�����C$nߠ��p��j/Ѳ�P��\q�DH#�w�H��
MŶ�g��(n��2�.$�Z 9xEE~�CX�ԍ����~�R��p69{��M�q������zQC�J'���}��-��!jpR�(��T�W-��h��:��#ع�RT�H�5�4]�p� Q��4��ؽ?�}�,yM�,�K!�sy1ԡ(���-�h���,c���Ć}x��'����Ɉ����2���܂/޷�Nڇp�R��ԓ�@9��MA�����ǟ�q�����呂@��*��*�O݁��O �p�ۦ&��p?��A)��`E��n_�3m����C)!�O�U�]h���f uN�*\gpp��ih��{��X��+p�M��~��'LMĢ��v��_l8�~�����h/��;��f��o�����j�!�ce���$���F��_�C,��JtQ�/UD �X�l��<�
��C������,�P�w��Їp���ΈN����������z~��-��|A�1��>�����1�].۲�i���%N�JMT���MS���7�h����2]=*WQ�E��Wg�v$���?�=�&�v�z�_II	�c-Z�w���+f@sfNm�(���H0���q�m��?1�>K��d^vk��9��5L �ݱ���IXUV���� =i9R�	}�uKKv`ٲ�ز�5@*��wƚb��8p���$�ԢS�;��4n~��\L� U��X2f�<$�rݒ?䡬�Wψ�L�'�B�@��s�Ԡu�i�	��Db�w�5L����)x��	�ΝCa1\�2��X,���M��qJ$8�.�,�jF9\�pˇ��	Qy�\ł��
葉l�	p�`̣2��EME�����21Qk���4u[;{�4�NB(�5�6/Ӛ���J�E�������j�>Ӕ����,�����������(�:z�knq����z7��dj
R�+

����>�,v�@���F,���߳u��x�!|�[�p��y$��e��+[Qbe�ؖ,���OZ�lѶډ��������X!�.��%LEr,��e�s]M%��c�~��(���UTW��t���y<����(�\�F�����-�$L����2�Zg�Bx�c%���N�=�	�^e��r�Z��<�p�Z�ʊ�@	B��d-F%���h��gQ��a�r����r}�}�3A@�J9�H$�A��3�;KӉ��Ew
�m6A���k��Y'��TU"�����z��T4�r)�.�!�nGt���nM]5>~�J��w��;l���U���<�lL[+!H���+3\�S'|�-C��j��X�-�wH����J}\���|��`�O����@S`�4T��ET*�e&��H�.C�t1���Mu�,�e����H5��zFl��D�`����E���%�"Ӡ��F�f~���X7��N�@�U��w�ݖW�E{��S�J�ת���2F9��u�\�%W	1�r5�W��.Em�(����Ҋ�{a�,�aG>
=!9���������0�!�A�Dc+�,�Y��c����C��T�6��t����$�:ۖ:�$�W#P5'���Gb�wX�i��j`�['X�W��x��i;^�	\)MN��M����X��\Ly[ϓ�A�r��c�B���/����O��z����ǰ<u�c�X�m��R��W��ǻ���i�������(T�N���}����u�q{-#ދ���!���]D�)z����5h��c�������YOf��3x7�:��Y������1�q!�)a\q�U,JQ�3�Q�!�hriFĹ3�+��y����7��JZI:��n�B�7Z����@��P{wZ�~n&v����U!��h�B� �L��'_��_^�����6}�b[�3��b�U�H�@9�)`��"3��M�޽���8��n'����>?����{淀�?Z}��i�kP�灚�����I�aEp+�;"�*V�b+�rBR(5�go���l:*ai�|T'��u��)ķ�W$��P�xF�o�pN%��s������r�쒃�T��38r���a&>{�L�p�-��lc��x��<�̏�J��1� P6�Y��dIC�v���T�`Vk3ܒ�M�ڀH�+�nE@+J��5�V�%�SHoղ����߳<��1��梅����KP.��D4o8���xe,0O��G~�4?���u>�Q��J�g(��s��=�}>��.Ԫ��g7S58X�'��/���5 �h��.S̨Ý��Ƒ��镗pm�z̭CU9e\%jsd
.�A��I�GV��%�p#�ʵ�N*��)<��3�=�w��榦�#��C�>��/��f2fG�2F�hJ��x��0������,E$##��qě�:dn&>�a��{
w��-յX6��ՔQ�k8���'�܌=o@"��I&(�a���P��c�e͙>���4�����^BYI��>$ǘ7oV��ƳO��j���;W�XA����D?\��G�]Q�����mx�;�jC��Y0���Ưs�v���/n|o�­�.�ݍҡ׭����ذ�06����#H��bK�Ҧ��ᨬ2��r&������~������r���F�겼?��g�}ل�
��(Ggr4�0�V��ُ	���=���فfyx7��m�)F��ap$�~�K04<����{�K��<c9pi����~��7��Oee%���������$]@������(ph�'}\aV���8�s ͗'ޚ�`N93ϐV�e���&)���q]��1��^>HP��\�,wڎ�'�5�A�(�����5��cS����h���a]�j<���d$���,Z�W��\�&���(��q��d���^���:�yANG}&5M4FM5�|��͝RP��\IRVZ���<'8��c�"�����j� q��{���L��vts���Z׀pP�=���A1퉚|��i�����F>�X��,��`����H�6C2�/~���><p�tDS�,�K)��(QQo��!����8ږ��^k:Em�(�Ƚ7���\��b�C��~4�L�u��e��@6N�;?|��mlu�b.�U���[A�2��ws�c��W����.�".�o�,a��*�7S1e D+���X�ic�j�I�,@�,���-7��D�����_��@���ZU�=4����;Ԥ\E�'�p �7˃��L�D4��� :F��yH<|?����q�bd���[��|��1��;��4#!�A���h�/\
QZ��0 	g�be�%I �$J���+C�3ǻ�@�/ӏ%��d.e�	���>�5�g����ٮ �ƒ����x��(E��DG:��<�r|е);��f��&NS1���1���aaa��f�#�9���ҭ?���1�N�"eY�gU���ȝ�+��A4,��*��yy�U�B��d��@Z̥���΄L��i�Qx��^LG[��-x~P�=��R���U��D#������#iF�2v�<��Ǉ%.�C�CMS���N��r�i�۩u��X���<�4ڱ��4�f%��su�V"�1-5
R��X�'��PR��7�+"4.Y��b��i ^@�hT~��鯱Sd�˦`k��_rA�����
�H/n&���[a�wܭ=��p�{�=����������Z��d������dsŭSs���PH"�=g��BJ���N�4��ǕF��Mp�e�ȥR���KXM���YKñf�ז����)���P���������ɹr� 	�J!�:���,���Ѐ�n��H�e�h�VE����Yhn��nq5Dls����M<.�U�8��+V���v�U��B�Kg�SFP��\1B�g�\��&�e�ea���r�iFM#9!�V��Xee��.ko�Kl��+GrQ^�� 3~v��2��5^: �55�ں���Z��L�@*�B�X5v�Ƴ�>�C&(ȑA��.���L���<.��V0�%��L�2���:>P'Kp����+4~��q�b.�R�+J�|�D�N ~�w��]2.&5M漽y,������>�ESR��b�ؾ�,6������M�+��9�OK3���L�	0t�5s>z��nVʆ��g����ހO��(�������>�R����K�K�J,31	 1>��5	���<��^|p�����c����8��T�ix�I����#�2�JP���F �͊�4C�Pp����X�t���Ӛ�'����N�d�gv�V���-����l�}�G:M-*n]q�0�\���E�3,�����ز%����Bkp��ߦ�C�����_�k~RŦ׶�ج0��Ĵ){ހja����o(s���!��1���[��8׎��X5�,���A��5��$N<�f=M��m]R�oŔ��������)+�_�����J8F�R;׋׶�	_j��<HF�8-g��E��^�9��12�H�0>��6%��J=^x�u�u�N�B���C���)S��+,�e�cR�$�I%0�1�hJE�cXݏ�޽#�+�g�n^�I�4�`X���B+b�9��T +D�1r�7���]�ȏ�Mƒ�n��?zl�%�0]��LDv�b?N��U������Gw#{���g�y�3��Pg�jƟ~�Z���b�.�rH�:��!�Խ�ԭס�g>���O��"�r-�v�/]���&��=�:g�y��d���ڊ��dӱ��kH��WX���q=== %}�u�9�KЍ�DZv^�7N�����cuҴ��ñb�R�f�rY�p��9��F/�/����z|�k�X~�X��A�����Y�R��#P��C>�&ڦ�^���y�����7N˜R�>}:���,"�U����\����
�b&Ʒ���N��N���իW�g��N���C��E�\f�,'�akjV�9�)��L�D�R�,]4�|�Xϟ�a.����&��`F��d�
�FW�%��D}j�5���߈5�Ǭ�Uu��f��x�힨�ܒ?NK��\��u�~k4䪹�e
匏.�S�����²����� ҩ��)nrh��,� U�"'�.��Њ5I�{V.���(73��yz��k1/_&�׎�wЭ�9�\E�D�� .j�ǊS\>�)e�0��ɳ~'�$V	-������#���BM�����բy��&��׌�l��w�@�U�y�}��-�c��v���&�n�Ѵ�.O�T�M��~��s9[�%�B��FC��PQY���>��������Cբfv��*s�;�f������Ck�؏p�knzi��(�LZ��ێ9A�R�"p������'�X�N���PLc����bH)�J��70�#ǎy�UT.���+�7C�N��`I9�NB��@+�c��
LT
.OH��L8)���J
���M8�� 9{�.ӘD0�a�$�v��a�����i��}	Q�!	�����f��j6�	�	N"�+A��U&�@���:�OمM�����������>,yaZ�L�ce���%����̷��G&�]0h��z20��2-�K�����$'��VbB�9�c���>��ӯ�$,*�4����ə���le��z��Z���@v�EQ�r�K��	�ќ�T�5HT\G̭�f�2o�l\0`Q��ed�)���@t5w8��� �B%h�ӡ�f��n{�خk��T;_�>���W��|##&�9B�<��;�skELa3��}P�-��G�u�`� Em�ʕ���Z���^}s�]hh�}(3��d�Md��Ǡ�X�>C%�ߋ��U���gj�v���C���	y0C,�˦`�'}n�uKn�׷m�}#i�Q7�p�S�y ��I������'Y��(Q�T�o)%c#t���t�VQ���H:�=t��a�]j��'Π���h�V!�ڹ�����P��{v"��;��X�5h�29�
���5)�(G{�Y�x|>�����؋}�f��^��Ⱦ��YĶ�W�*v���'N��uH�T��.F�lv0{��PdU_��D�<�=���.Z��H1��},
�PBԷ\�9y!�y�C������q��!5b������Fh�C�|�Y�F����� kG'�:�k�ܳ�t1�,B?I�/���Y�`i�[D`�����3�A
U��,j�:+^ڊ��.V��ϧ`+�3���l<��+�M/�Uu2�Hm-�2���m��Z�+��zL� 5+Q��\QBY�3w����ݥw�9h��-)��&�fZ@�٭�q��U���d�O����Y�m3�*�����GDY1�0SԔ��48q=�i����>����WZJ�k��y؀>�Ye�"i�b%٪����be���8K�%�x�C�����`Me��E�ӤP�$��S{������W�lt��B�c�ΰ����r���`9B*�(����$��-�����F 5:�=��=W��|�v�o�f0��yh���-�����纱��]�C��擜�4�|/&*?�,�����_���|�&L�L�b`�o���{���`˖WE�TQe��x��4$n�Q��L�{Ih�bG��06���T�~������$<!C+Ty���h&��M`�w%n�Vus�����xP��o�n�7)�rc%D�S�H��D�y��������_�7��d�y��I�'?�o��5l�,�.�ӷ˧E���Y:�aF1�:������z֭�%J5�!��4��p�[�/�==��Ь�:��-�F�t!�"�+MGt����8Ve���{�џ��FQ_W�Vϟ��]3	O��E��cʩw���r�Wv��΃��u_��_����x|[���et>kT}!֘T�а,��|�����̙�cy�˃PRPU��"��
�{��%oʦ�`iWo��=���K%��`!�C����_�k[�(++Cmm���cl�u$�&ɗnUڱ�;%�$4��yG�Q�hfi2�2!ͬt5�X��Xmg��\U3��1F�Q��實� ��`�p��b��)�R����8C�}��/��r����&5�O˳����-c��YTaH�att�q\�k��
�m夦1���S��d4�S��r�����8u��JV���fj��IM� ��0�U�'��,�6�+�w�(E��D��X�Wl�5enw�7r��N��gM�t靝9�3\=-,v�KqZ�Ͳ@K��1��.��'�g2�z�٩f³8Kv��x�\/]&5�_i��A��y�4��P	�b�tkey	B�
+��DӲo�x<U�Β(]�XWԶ�l	D��W��B$F]M%[�4�ɔ�qby��4y�?W�iHڳ���^�gN� �,vqQ����Q_�7�2�8j�N���
�,ڝ�����lq���9U�&;4,���KSq���p�b�U����꯺i2���8x�W���ʕ����nkE `�6N��@K�L�5�N�LCwh�����������a�hcY6>[a d�3&d�y����M���$����Qr����):Kr�-�w��k�YB6h��6�i��$Z����,S�L�s��3<Y������+� �����6�Ȕ�U�(E��$��_S���
7˃>�Pb����2�N��T�S������W�ȘA��W���3g����Q;ˇM��9B�A��ǹ/K����&��`P}+��!��Hըy����pփ��EXX�a�Jt�<h"���0P�NfV!ռR����^W/������ZD��9��KU����)�@��~h�q��M�ӄ����M4^�����k�3/y��@NT-�Q���f:�E�x!���<d�`�-�-Y�	D�ª�|_猄�W`ړ�A�Q)��~D��L�=3�����r$D�g�[a���F�}�ȧg.ת<*E�<� G<,�Z��s�'�d���䢦�d׶|=6A��e�X#�������8M@��J1��@C;�&�3X���>j
5�tsvL��yH0�Nu �a�,����(hp��!N�q��}*:yǴd�]XF���ٿx�k\������7�0���;䁥�gٸ�I�j9
��w2���c��Ogei)j���|M�Ҏs:0Y2�J�D��=�����";ޟ�����%�E���խ�##{8����۽{���(j8�3�������	X�*� ��e�"������ Q��i�C� �V̖͈���*���L������X�q�	�iH��S*��<'��y��M��=��O�ຼ��.t6T���?�Y(jh�O;Β�o����9�Y�a���B!n�I&.�8��\�&/j�?���)y=����3�f�\,nΪD4�����C�H)^z��?Ƣ`u����\B�K��n5&d��4DӒ5�E�kg}��݀�->{h9_dtK�FYsA��#��3���T��ͪ��9>�ndY_�d��|�R^ȵ��3�w�}��5&ٷ_��8畲�����elҔrl9`� �$|r��B�0�G��)uX�`2n�q)*�c���l��Ʊu��8ԋ�����3���;P��j�NtN�LM+�q����j<x�4�*=�p�4�1ʠ�[�.��6b������z<��f3�Bt=�T�f΍�	��`N}�w�Q��zB�i�̛u3n�Qg�5�iL{�P�C@]#vg_��.��KZ����0�1�:�Ā��ȅ�gb�h]l���UX?d9����^"և��o�ZQ]�F�
V#Q�����;q���~f�K�D,�!�w�/�IakX7^5�:�U]�/r�I?ז���:_\��N��/n���D=��R*9�xN =3�wgNw	׬\�?]'�J�y�?�/��@=��U��m��/~k�Ph��,�Kh`Ա�Qy��9��,�Q�8g:�Www��{���jK0��=�Y��X�\��_܆T��?v֟{��ɣ��:��Jv����,�%�J��KF2S�5$�&��C]��wX�{`����yv���N����X�+ L��"�9���8-j����E����u����Q��UL� ��V��rP��ď�$�%�S���fG�."�%ˇUZZ����*T�����5�.M+�P'cE/h۪�|��UP����o~Zz��pux�� #)��Z�
`��R{|�F͂�8E�����T�����my�����E)ʥ.'�����P=:���k;�B$�� 	�&+���i�m�{x�����ݵ��ﵷ+�W�CpmQ�0U��@T��ǯoB��Mx���ab9��
Ӷ�����w�\6����䕐Q�@:���Ǡ��`��ѝ���{q�H+����S5���C��ʝ���RL�5��6C!̶NǞ1�@Q�r����k@��3}ƅ(6��S��oZ$Z�u�
&'^��S���� 0u-1�x��Tۋ��+lA����A|x݃ؼuQ�pQ4-��"r���76��&�J����yvg#5��00���h=�E�!��,��@+�}��m1�-�LQ+��E�+V`�Ţ�s�����6
��)JQ��w��|�}�E>դ�%�>3�T��ٰ�Q�b&�K������h����Ոm�;h���i3����λ���Ȅ��s��;pt����ҎX��y�����ME��?������EH����JJJ�	7��ޘ�_)C�Yq%Vxe�`�v]6Ǻ� ���VQ�w"�`p�f��=��9�� ���ByD�<
D�S��R��w_��D}���-���AS�Z�߅�3��e_�����7��P�=y�*�_��Fmm-��8hy���0�5��!
{��<Z�+�Kޚ�tP��cEy��R�/��L|#�e�i���QY�G����<��z����2yE�x�@�U����ܹ�0Q)8I��n
�?%A�ٱ��q|1������C�-��ᒈ���i�l���뽉���b��)���o*�����0<Ư��"���f�$9�NN8ы3]��"R�|��Wggz���(�)�ҹh�͝�t��yo�垂K�L����m���غ׮�4����s��׿yO��<sj��=)gʇ�q�ik�ir���mҪ�m�ڭ�RW�U��lC"���r5��4�U�SP	�l�孳�]i�_KZ��S�m/�i�+Ls���%�#g���[�1�~�5�%�KbZ��CC�b���,s�	�kU4BRC'
�a�m��0J�����"����[ј�%���;8�=Gx0l%y!�e>fN��چ����h�
n��k5fmC��g��@�кճ�v�t�_l8h��x�q�L�.��?����H>�2��\��J@�?|$w����Qh͛^����x�	���5��:o����6&hM�)�g�ZB>J�?�O��G�e8~	��I��Qd|���Ƃ����A�N����;�sͧr�D�`M�tw�y2Jŵ$�����)M��)N}���S{�`�z{M���I��u��J}^�6�J�f��,��`�z8�<����"���sֳ���ЧE%	����	��~ŝ|H�M��F����J��`��l4�C�V�6�9� kCS��q�B���6?�����ymh�t�y3�m�o�{%[����	L�M�}E��m�عۤT�l�";�x�h�5sd�&B4a��*�藀fb%������۴���_�1��k$E���e� �w��ڊ����k���6���Z�~����B%�2�`��c�8�b%��� }��GAh�]�K��ڻ��?��ǃ�љ����&,���א\��|{г��TtD�R�AiN�wZ�Eb�A�^%M�d�g��6��Hۨ�0h\�
R4��Øeǉ)��1j��K�B*���ݮ61�w�d���r4ٻ��4z���d�^W�盷%mN��܈��N��&=N�c���dHe����D×F��6�:�f&����f��L��q6vF�4H����0em��|�H�#��9y$4H��l��";ޥy'r�K{���%������P'��+5��ڏ����'�<�sk�p�}8�.B%&е���� ����ؖ̻�1^|5y�P{l�R���i�����
5�r6r;^��Of�=�5&5��8�uV�5��#����a_RY0G��dyļ��#�����E�w�*]��k�j��$yy1��MI+Բ��e��Eh-��Mt��Ֆ��ڤNqΥ,���t��N�&Z�X�6uH�둪��M^�P�,��M�jow�	�6��Mg�6Okn�T��:FP�E(Վ\�� ��뭃��y:O�[P���(��	2v��\�`����#���w�Euj����Q�j��Ă#9mS3����f�]��:���`���߃� �)ײ}��6���W�ǄJ*4����w�[�s&yA�qg�d��m����CszPؗV;�����:/d��z|�{�ch��Td��ɮ�v�e�$����/�zˊQ���
�q��>.��`S)�h\ESc����]�'�D�65(AO����eu���@5>��/a�y3�2��:�F7�6��6�~D��p�ݟ@�*���gԏ�6���C-��hC֏ŉ�6�[n�(��< ڤ�R;�ڤ�3�-�;N�(Im�7� ����"go�!m�CM�J纮W�~���)���� CAsz�0i�J��ۆ���~mctce��I��I����&ϱ6��H��i�n(O���s�mc$�XM�<��[�9sn}Y����d���~�^PR��g����NU���ɤo��eWq�]�F�[&}��|��_ m�]����gb����k��,�۞qW<ul'��Ch���ݝ���Ob��y��(�4���[���}	㍞���O�'�r�-�C�L9ʲ������pW�i��bfP��"��(ڱ���Tj�"6=������5�8$����� ��eW��y91����e��̸/�@?q?���`��@��3x��C�������G���,����%����AsM#*�6�O��hФNw���η����k0��5#� m�n�J��Wb�3lYQ(Y3��h������A[���Z9�(�M}� }�-غ�Mކf�/����8�G�M�&�6㍤�Nkݪ��^B�F�l�m�Zp��^���N�օ0�Le�=��9���2'��Gw/N2w�\̪$���p����/Ʊ3g�%�ZѪ5u�K1):������.��Ӽ|{ue&]]�)�A�����<��=e8~j;
�dr	{mw�3�D�#�G��̈́��l��I ����⭷v��	�g���J��Գ �#-� 1��%���_��c��/\���IR��]�3����ctxt�؍��>�.J´S��H���C3���k8��	7/��Eӂ,�<���!�Ez���|8���ݏ���`�2*�X�ga>Ns�m]���r���*"<ߊ3!�8rp7���B �榈YA��P����˧�%��Mb�7V�)�ME#�4�l�z����z3�z)v옎^�=;gӴ�if'i�7k�lZ`��I�O�*++�Ս��=_Q��kk�/��ӯJJ�X:�Z���=qn����y��C$������e��e��b���Fk�*����z����f4���g+z��}���Tb�&��^��1Lγݽ��]��gF�DY$��y^�@kќ)x`v-���U����ص[Ŏ�>������>��ě�5���nP�@�l�Y� ��:��?ƂME��9k��l�$��`E�c��l���\V��">��1�>=L�1��������o���]��P�������G�>[�*�����'�Ǚ�dgy�(x�ڂh[45��v!��]^}�KL�����͙�������8|��u ���$��ֲL���M��NQ�.�~*\�x�]�{��tf*B
Z9W�L~z�,�T!�j���Ia���B��y�����(��S&VWq�4�44���/u��J^7	�o��&i ;)��0�t�Q�k1,�77x�\�s:����a�FF��B�W<_�o;�`�6�2Ւ�B�����%/ņ(*Br��9KW�8%��E�c�d�c�����R4,��'���DT�U�Lm�}�9Փ�`y�C��	�x�O�>�����56aQK=f4ٮ�����t���1)i.�|��wZ�E{���@g�����ۇ�џ�>�n,�e��/��	�UvX`�0��z��c�MV��I��Y�[����/!�B�����x�:���ټ>��d�F�m���4u�)���f� ��Ib��:<2����<W�Q����M���d�5T���'��"�H$�9�
���b׿����)��xJ�Z��F�I>{̧��}��=��.����%:HCA�}�$y���I�������� �q2�e�*,��Ì�
�{ wsx|�����H��6e�2��Y��Ӱ]���2�p��S��]�̠�qmDN1YJ�^q�+>>��?鏿���2
��K~�:�;��������-��
����TZ��҇��ŒC���R��s�Bmm=�]�/�u�>簢�
?�=�}��1&Ԉ�r�&^͂��-�ԺF�������ts�5M��	:�j�Ґ� 1#���u��ڏ�7��ї�qS�*�ħbu@EPqMX�����)�8��������q��I����L�_r��L<��A�_�X<��g���F��yW�Xr%xb�^���m��_U�� ��s���<�p#~�m���Dg��I��L�z�(�h�3Y�L���+03D��z2ڨ�z���6�?d�c:�1�D	
����t�h�3]It1v���p����&!�f�M'�v�;��mFЎ.j]$�k+�f�~��yU8_�m;~$V�V������{+�Y9� F�[#�y��I�T�D��_�_~Z�Š��Ǻ"G⳯_?�fU�����*�8ζ��VtB��4G1UW;�Ͱcɰf\�T0�NÔ�W߄{>�I�W�32N?2�װ~e:-~z���?�, c�s�T*����Gx}��L3'_�Ǟ܀�'/k�㇠���R�FtK�td;N�<i����/�݆�Ǫp��⋬2S�~ zcx��8A�`��}z�սj����ܤ�N^��$���a�69~�wX����o"927��%���MJ���������#�0�}Ǻ��gܼ���)��g��Gf�7^���IW�cG�[O��ګ����q<8�������k�O�j��~��]���V7�ts"$�s�Q<���B3���s�߿.Ǉn��P��k�f�r�:�JH����?�>s�;�B��?��� ����Rxv�뙡�DR�c[tD'��4�e����3�s[�8�x �i�ޤe]<K���6��M�3�б�q��a��F�~e��+����Y�%����65����s���K6��QBLg�������6� I ����qr�a���j��0��5�`R��,��j!����s׽cŪ�q)Kw�9��g��`�yu�����͔�R˃�����XT�������g�[��a�d��4�I1f�A�/2�X,��m?�-��6���j�6���������g��A��!�󨤍7EB��ꦝ'��P���<���N��~��8���&�:p^ߘF���a�L&�ؾc�<��fo�Zm*%>h������q��d�p-��C�6����3m��{I����U�;�&�x�`�H ���a�sZ�o>v�4�wZ��i��Xg>������6����h�;#�i�/4IK�Y]3�_ժt�QqJ�3vQ�i�}q�M���B�n�d��F��\괭�3�ƴh�c�bW�6OoӁ��&fJt�׆�(D���9�_� I�0��=�C�߷�_��K�F51�W<A�]����x���x�ás��e���G�X�t�-Y�R%���[&�ص��W ^�'O��@�i<�a��~ܺ�D=W��oNZHĄ���J(�̕-�2�>o�9����1G����˽�Z��	�Ng�Sؒ0q�Ɍ�e2����㛶5}f�����6�A40F����>���>�b�p
�zt%�:����'��W���m�q�0�ØyN��ƒ���g�����X�4�ŵ��Kqm� >�%;*����5:�}��)6��sɨ|��3��VX�}���d���MM����S6쓾K.g<�Z�R�Xϙ���v���{��������<p�9p9�;U\��*x/���a�$�'�I�:�iX;G��_K��U��vE'�z{z�+�2TV ��øP��5\EF�iP\�����Ms�q�hg�P-⃎k�"���<Y3�e�4����gln��9�K��.��I�k�Ů#i�%�9�d���B�$͛s�)�|�+�&*�]����78E.���,��6��p1�9�M���G�ղ��^��������t�yM����/�n��tUqf��i�u���pYq����J�x+�;!f'>I��5&d�d��s���~O���5N����c�#��q���_n��y_  +�${����8-����ߋ�:xΟ�BYc3uL���h����������>}n(�I��0�V��2-܅O�X�#�-A�q�c� �;}�K��}��x�R�kjY�>bב,\
m����Vt�bI�(��VpI^J��:<,M'�Kb����;W���/����L������A��ƒ���Y����)�y�l&i�k"��q]�s�����2�$w�/��>��u�w���Fa��qܳB�B�io�]X#��@��#��϶�hZݡ�)l:�G�z�7�xȂjE�su9ȵ(�p�/?,�E��4�O���\�,iF��QdϦ{�<|e�Z�� 9�o�uV�h�7#�'�4w�r�Rpq?!�١�޻>Fv\I,�����!�ևj��7R�"�%:9�ND�6��#�X�@��#J\��K��)�5y�6ç���)����c����4,QRˌ�s�Ժ�8�K2������1u�y������/q��H���r+����b��Q=���f��#t�=o��&����ζ��Kl��kXia�揃ˮi��6�,��=n�0���\B���f�̓9��d�\TL�Y�4APJ�=�!I҄����s�L a��i�?��D%!��&�1�E�ۦ+�d�_�*��y_$��iS8�ӧa�EQ�N�8ʸ��0-����8�IJ�E����'��Y���%3���ls��2}Q�f�d���mc�NWҽ�tk�Ӻ OS��<(6��ÙIa_��l�������>\�w��	J�,�����uo�� P�.?4��Š�Ɉ��ql��Xi=f^s����o�Lq�<I9b=�4�m޼�hljB u�1 P6��gϲ:��a(���fI�t,�sq�ô0�υ�I��8�����\vR<�A+����:�+��t~U�/k��P򌧫K����Y�A�����	f:�5�c)$:�ÒD@#< �i���Y��Ǖ�����������L����{OsT[e�,M�tv/��5����<�(�*�r���,S��Q]q�@-�I����F�Q,�߂�� ����Ӎ��A���&�0��9w�)9B�l�k�ʚ5W�w/Gcz;*��"�:�8*0������߷�u�S��\-6�C,��S���X�]�eXT�/���T1u혢� ����l��s��VG���k~�m!����t��(�\���S-A��S�̚�A�1���7��Qj�����
��B��.���+[[2f���@h8���,��ͭ�Pi�ert��r*���A��|(lkXa��O���8w�Vrhp^w�_B�b��e�3���,���Z�����/]]�,��'K�^v�����^���x+�!�y�9+
�n7/Ŕ�fԇ{�G-�J�f���x��$�2h��ǐ�֚���K���~ KAYY>|��ز!ԥ����°l�@V&�$�vg�\{���/���O̢zdQ"�:���95�Tv����A\*�&S��!g~<����F
�6�~C$�FE>d��s��>�x�	�, �aR���1� Ә0��!+�Mr�S�f.&є�L����Y�uW���jg?��&�GJLO� �)V��4�4}���5Z~�L�r9��?�c}�e:�q�������}6n�G>�oZ�Ih���d�&����]��5.�F�t�ssJLp���z���Tȃ�Ht P��!���=x��'�>S�,�a�����Y�pǘfh� /D��)`���|���� ���2L.���~K%V�u�� ��T�5�cf\�b�8�{��V���s��rs=���kk⫟��~t::αA��U̌���C`癢͑o�^����f7��!^K)l%lSn2{���YY������� ��X�A� /���a�s2ZG\��z�@��0w��!02�{}�֠�K��7��OY )��Y&&\�Vv��������O��q9}N��m�5+�EgPݳ����i`���(0��3K�0v��~o�}օ����f�s/��Z|��
4�<���#��+j��� �������.�l�9R�3�g
k"�4s�S�߂�,hϋT�\Q����=���P�pe$/h��k�t�2ܳ��t��9��e4��j�j��ah�G؃Ju�z�������A᳃���bf�0\��P�3̇,��2�n��$�2ڻ���w��籶z��1�F��f_d�}�W"-W�m}U����qv�*ȧҊ`����X�0ODL���5(
�ϩB��ƈF��5��4V�"uQ�-���_�=mF&�
6\-��\H>��f^�^�$�nM�3�T�;$�ΨŴJbƥt��#��Zۢj*ӇX^e�(�lw8ޭp�0�,�x.�5�cFfݚ|h.�S�f�r6�Sl�^�p����5G�~i9~�zb".B&hZ���~�C-hJ�l7����?�R�b�\�&�=��៰}(�ʚX�h1�/fl����,2��y���e��\p�wML�H�3�ɞ����i�87�nNf0?�u���ͭ�44Ku6��5�%1�,fQc&�����=��D����89Wo�F$d����P��#�uX��.��uA>;���X��Yg���m֤O�X�̧���<�YA����P���M���1В��U��s�|�N�4#�KQ1掱b���0u}�Vօ�Y�0���ۈ�����c�f�Gl6���vZ�#��&��q��j1?U��aq�Ѐ��7����D���k��E�f�<��Gɲ?#��u�Yw#y�Q�N?˞����?��{��q�kb��Sa{��k05�!^,��@���l��m�<�R�c��q
7,��C�B�qCM�C�3��M �A���f:N�[���r��mr�ø�q�ڦ5	)͏ �S\~,1��V����z��Db��a	߉�ha��$��x��� P4h�>i!����b~8ɡ�����C�W&m�d�9�}B�&��y��--��LZ~��� f(��%��D�(���}N�l;�#���59�c�Zc��8����Dĺ��ԕRkW�Pl&]�͑����.&�ψ%�"	4�d��'�K�T�Y(9��`奦����j�ê)��Ǹk'0y�K�L����#�NAt��C��}�'�G�2/������Gu��yZ=ʍ��rx��r�M��SO�b����gӠ�cc� !�U5����,�z���u6�Is�1d�:)� Πza��|6e��fԕ�����;
8#1���^�ײ
����:��>�4vfp��j��]��`z@eS8~�k#�r:�m���a<�Ea���1�p���VAQG,����9����}H&n�<s��hߣ��cX���!EC�2�qO�/��
��Z��A����,\����cwQ�	�u�i�8|����۱�p#�_����������� ���D����s� �� D�Q�H%ˊ��$�~k��Z���>۟d��~ϒ�u�,+K�(�")J�� �yf09���U��nUW�(����JCtw����{ι��gfz
c�0�C��8�E�*6S(��fk�UI�;��r���AӨq.����^��P�7sUQ����H��)��{�u^<�}\�*�ii���.­xe�Jj�D��Y�	k�<�^]]�x<ΉV���єn��z&��_�WN�,�~N*N�o��
޲�:|���M����S^��lt3��kt��B\Qއ�d/y ��9ppG1�����X�s55హ��4�t�T��TV�gR�`ڕ����I�$��];��܈�"�dZ��YN��C��+�Ɓ#��@�ھ�nz��10#�g��mE�
_^�h)�0�3��ֹm�z��{�cMŐ㓩�������ëo�׿�CoS�8�&%oγR!�k��.�����!~�Hm�uU[�� )�H"��u���t��P
�F���J6�}��p�ʎ��G�n�~�T۶ךJ�=�-�o�H-�a�}��ҎK3�D"���B��7�2��O+Ud�Z�_�Tx:�o�OQA2����BT�21Yo'z��Y�.���=Xi=R����\I�G�J�I.?�ES�B��X�
�*d2)T��\�t	|��>��A"`D��5�J�vn�z�y�*����$x�}^�%���`�l�'��Ѿ��Z6�yF?P^N�ߌ�r��GoX�Κ�*\Wqa� -r�X�iܹa�������f{��?n�'aH��:�&��O�Ө���i#2���B$L�Rh�Ü������Tk���oS��[�By�Y�x�F�f�ִl�v2#�]���n�R�}";�l�aQ�ɧ�{����{��{R�\W�{�o��ot@L7Y�j������3W������&������ -z�R�/��ʚL�"o�a1Ϋ,���������I�(oK�)�Na/,�M\۴�L�΢:�B��P�5e��-jW���9��0:����� �\$�j����c��Ɍ0�e(���"#u��-�G��v��y�O=W��b/�C-V��X�B���B�Τ0��|2���0�,�����0��<=e��ڴb��}��您�N?'��ޢ�"t�V>��7%4�m�E�yd$ib�/�L�J1��f�I�p[c��,�^htj��A�}�ȧ��E}3.ք{�l�x�^���b~����{�ؓ�՚>�麢�n�����M�\�DK)C8~��۪�h&xײ}O"��n�*�s��Úl#��W�CH$V����x�i|��돚�ç�at����7�ۢ۠�S�x��I<��V�NE"C>Ǘ����#`s.��z
�/����v��E�T�~��?!2��6]U]B���U/�p?>qd/����������J/g���ጛk�ٟ6�0���5?7͈�">��靈v|���l���be�ϲ-�_��|��741�<���s*ҳ�Fq��Y���UFGȦ�Ma!Cs��^g$ݱ� ���׉)"Jr"_�޺?�c����?��ܸS���j�����C#���)��O��.g�t#g�j}��>HZ��m���%�㓚�@:����2�%t��M��a6[����C/ ��^�-�Z�)$����=U���ZSi�������AcJX��z�|���	��w{�/?�ԙ�8��b7�ЙK��[`��C4�fǢ&��=��?���.&vF&���~̀H��s���\kڰa#6�Y��$?�?ǒ�i8�/�w����]�3qWpH��[R7c�`����v|,�$��9G�b��6�*\.�>'S�N$��P8�U��"^V"�5���_Arq�ϟb'��Ѧ��V�M[ ��Փ�ܱ��}�����i��ZQ_�'q�T��w!�b�F�d{x����*T5o���>W��fw;��[��H��j�:�������;Ԧ���p��b��|������̢7�
5BR�O�G��wQ��?y޳2sHu��#�oW`��-�=-i��}
ن��竏w�߾	U�|C[��K�;N���Ͱ����.��+�S�]láC�ʿs����q/���\Ou8� |�c�����i�<���U�'�u��:��*��e_x�dF�Ik8��6ĢQGߦFC�U\�кk~o� V��B���\N��_��u�DB�L�2��>e2I,.�)[*F-�)�)&V�����e(TD���%�TF�9��e"O~1��-?[l]Řx��*�U��׽��F㦔s2�Ȓ	i�!�A�\�es��$VT]�����j�a���M?Q��M�#u��Dő�Q�x�Ķ�� !l�2d�y�a�6��
�٦�|�ы~��e����lm/�K���Rh��S��+�}{����=��]�ѐ;ǟY�+Ȱ��*s�:t'�����,4���z�y;#N\��>�4v�܍���W,��������~�dG*9Yҋ'eic0|$w��C(3��<1��-�#��%�
��ңX�4@����l~�w��I�N�P2~��vwRj`�1�'Ϝ��#""�K���M�W�4�|e蠊�w��KQ|�:�x�{� �G��@�!:����o�
�C<)����$|���7��=u:߆�t��O�4ҧ�9��d�O�/��&����
�ħ��C?�1�fn���ލ������NS�|^�ڄ/?�2z.]����tmb�*5l(a;C�����Wq��	Paz�9�>m�2������՞��,
���U#�������CƲ�.`��3�i�>l��_��Q�%��ΐ(�}a�h�����)��q�ݧ����0���v�Yp*g��qu��o�^�����,ۃ��qI��W��9mO�䉗�o%��<�!��M���H$��o� ���Ո%/E!]��{{[���\"x�-�JC�8*/l��r�U<��$�{�[���P;��׹cߝġl�����o��"�����R�b���
B)A+��j8�]����%��5s
%҉?��m�׭��fy]�WSkc���<�fH<�8aj1g%<L^+O���Tb\e�(`4�Gv�RV�Z_R�'05�����P�7]���m�?�M%8߳�i_`{,�.�o��$� �R2��SϽ�]��T4��TW���|�5�F'~oKtT+�]?h�X\�^֧��A<�y3��/�-�9TO?�:Ws.-�������+.:
�X��iIh]9Ρv��#"�<��x�g�e�V46����k�|z��)��g�0P�BO%�d���#P��bS�L�VL��raNM̴=��02��'p�͎s������u҄sW���4+D{���%X�P�n:
�T��d%r����.?1��Hyjz����T�m�k%�Ǽ7&_CC#���x.�����v~QH��Q��H�{�.fzz��[��v�sv��#8���)ivv�?�D�T���W�1�,� ��
���:�h��UUU5����Q]�x�LN߄�Du�k}��>4�vR�*+�x�� ��P�����q���"a�W-��fj.C�{P����75	�NR'l޼�����8֯���!���>w��"t��s����Z���bjj�y��߲����ի�N���4y���gM#�!11(ݧN�#tw�u((LKK�w9��}�`Oc^E�
`�[�5y ��$ #����A����uĆ
���G���ƹX��eؽ�]]�$��pv��	\Ia��]��nkič;�P]�$��"�^`��&�f�댈+ii�Í�oF}��98�t��^9~�/��Mgr��v�
c�*F�"UHVnw|˦f����cH����*yW�%|^}��v�L>��ϸ�i_C��,�GM>�I�].��ӆ������;q��qlݺ.�GEE%� ���=mn��G�!��`�mm힍"�~��q�N�<�Q�Q,�����@������O������\����i�������a&"�L.rE�1D((Fm����Gv�^-=&�B>�_��?JcIixx��;�YWW��M�MDt�~q&F�*��$N�3:x(?q8�L�ӯ¶���R�(E��l]W`-�^d���WB_u��w�f�SF! 8K��Wx�ң\EV�])ԋ�͐���x�+�[o���l�v&�Vd�|ӓ�hX��7��*���cC�6֌ �P��%����:�[��'��!_�6>����}a�7�f�L�M��ڦM��4�t�:(����qC�ylYY��с\���$ZbcX�j`f������(/�u?��ݗ�\1�����j��}��kID���r	/m����X����d3Diaa�oZ��R��qTMM-|C�ƏFc�\�6�b�i�S�SS ��o���� _N�N�YU�Q���68������]�G7��@�����5�X���z��������t�/;��%�
L4	�_���C��v�q��Q[�O�Z�K�>߉�1�E��yH�.�(/��o4�[}}����^
I���GW�H�>�M�\um۵��e-�ח�1a',�����"$���lq�v�]MI���ǰnujcC02�܀D��xiW�������ό�=�ɫN_���c�� ZV�p����*����>�����A�N������D!lo%��f���%z�(槄��o�ԇ�س�6l������G���FUh;֭fDK\(8�Xr��ÒF�RT�m�j�z#��J̋�Fш9��~I���+W.aӦ���:���.��i�;s!�&�!A����1�>��ޫ����Ss5ĭ�e(�\J%�x��l��Fg1��T�T���㫩�e"��^J�>TU��MN":�_@�W��/" �U�nd�x^�;�+¥� "566In��"�-���$��\�j�2� n�8*z��JgN�����2\��$t�K@��<���T�ˊb�����גD���gE�i���OM�N *���SrA*�J�q�t�z�J��>b�3�}�� �N��X��R�x5Jcj�3��4z!�	�b�P^���?�|���.bͺ<w�p­K�)..I��L��\����{yI���&��9F��z�oʳgO�M@�����K��6���9m
��Ο?��Cġ� �N(566sn@�D���D+�[І��k0D?�F������SO���z�(�W"�jq��J���������;�����iZP�~�v��[$���<��9"n6���O\0�#�w��@�֚��$vW955��Ǆn�hh:]G,�����x��dP5l�2�\�he|&?d�#57���Ym�)�Xi���4w⸔Έ�&�Tf��2�����Jt�.3�Y���6%g��t����I�p�D����g��<�4B��ݠB�+�Z[�}uz���85?�M�;pQ�{�ƕ��l��Rɿ�)�s���/(y7���Blk�О._�d�
qO����vI��S_��s�>
���W�Z*x��{����\��R�a$��₄�!����C����?}����'"n�ب�YO�#+Hn;*[>����(���(2�z���:���?B!��fV�~��Y-����I��P�����wĀ☤Bz�]@ >_5�Ȍ*��%�\�7�t[�e�U�Z���ny�`<�k�|p_�5��{�|"�f,��-���ol�κ�����6lo���J�;o؀U�����b�\������ç���y}�w-�~;~��Mx�ɢ9��㶏������yc����C�P�T�C�K�B���C���V���%����Cڔu�C�@o��-+*��1QѨڂf�����5�7UW�0���,,���="�i6�W��خX)���T�G�ސ�?���"�p��s�f�P#��ه߶G��c1�
jA��6��h���-[�r�%�$(@��i@��8�[�Z݇Ж��>��K���i�q;7��-�ޘ>�mp(���al����x-�i.��K���]J���%Ax	z(��՟Y��r%�"|��^1MZ����v���'�{H7��L- ���9)�?�a�x��*~���Rr�F$��cU���܏�>��,ɸ�PT$�L�e�>���j��s�Rb�"܎�����A�)I���oEU�mr�����S*����o���}U����S[�j��{���N���&����C�����!5�u��1��6>�Uz������!4�Z^�'� �'I�R�(�}�'*�m]��/����q80ۡuE��K�k6y���c ����%1���޻�|m�� @�XZ]K���C�{D����Ek/�arP<�T7�Y�.�.c���;]�&R����?��W���j�˅������:�3�H�{��%�3��k���*���p�(_����h�m�G�Z��I��}�0��噚xR�.�$4���R��[/A'b�ҫ�C�Dyp*�GCHJ�H7n�m��mmm8}���GA*��p��e���apL9��l8U�K�)�91�����;bA��V�,�vv����EF&1��]� �B,��뵍9V���\Q���(_[>���x��$p���(�)׬A����h��z*�'a��u:κ�/�N��qc�v(��an�"�"����zO���qD�i�6�ݟ�ڵ<W�z"�O"�V��X�$�.��8ϣX@YNX����՛�E�0<~��Mx�E���r�0�ᇦI���B܈�E�y�8�?���
��d-�p72�+V���ǱuM"�IY��yiT�5�\�sJ1/�C�l:u������-��瑭Ցge�e����>�����P�c7�oF2#L0���ĉ�عq"ٱ�>P��3|nI21�q���!��].d�F���vǎ���[����a������^�7��{�
�(���C��W}}=n�n=�[#�Zb�H��+����N����mo������\�:�\N�T������-d�T*�'�-t��-��Hϼ��`��VE���w��c�)D1ޱ��Qd{��6�$��lb14n�KOObxZ�(��}��vSn��������7w` s�><"`�}����0~���XU��t�7����z�ab<�G�>숼N�*�ኄ$*r�_���[�?(:��H˿�ӯ0��?���s���t�H�p\�N�k�;���06�O�=�P$��;v���&��inn
s�����u`u<��Q�5��@��f����s�?q��_?�i�b�Tg��R������t�]7�wn_@4=���[1�ɩ�5���G��#���7ใ�q����G��144��ﻭ	oY�����#X4[�{1{k����e�w���z�ܜB�˥�� �f�4�岽쌚�~���X/��U��_߀��nLFv�R�/��i��s=X��56v��I�n������Q{��ő�19���n�»��<���b!����D���#hɼ��H���q��^X7y��B����-3I����wܴ�u��G��t�m'���X|�G�\w_��㘜����6�U��24�����"���2�����ލIT�_f3��K]��r}#��z=>���=P迸�J���B��D�i�}�,>=�@Y,$o�ĕ/a_����Ft��ab�~���[����#��Sr���cd�O�Ȏ%�����X�z[�C�N�̬�+�\ ��F��#��/�8:�2�_H��z=��pLv\�PL�	��]�wp6�M�{����R>\��g�7s.��q���҅#jf�X��z򯶄�ѣ/�ؑ�"�"�,����ڼ��
J��.\�qģ��VV�8�j�Q���l���([<�b)i�s�I�..����d�z���p�t|l_��?:�w������D?��]�Ln��W�G{U��E��[��˽���cj��^�G0Lg�(T�b P��Y��8�j�:cGijr��旄����1�!oI�]OW��1�>�a#���Z�M<j�"*��G�������زu~�ޕ�u�$�����Iē���;V�D�G��+?���K��\"� Z��$�ezAM�7~om>�İ�Jƹ�6�?�V\�f���@�#� ���MU�l��z �_��R�,tO�e���6���d�ˌ�Y�r\��L�K�Y8qd��]D��MS���8F<Y�xhܗ�h�&���b��`}��Hj ��s��\��;8v�qvr?{L�/ɸT�R�d�	5��ȥ)�B��MP ����d�H�%��Crg��~��14��;7qҪ��P�z���ȇ�1�X�G��E��Km]��f��8n�j
��-WP!h#!a{��l\�o��'N����c���s��h��#�RJUlg}��d��zb@n@2+CSY3o�[�O,XZ����F(,Ƅ�qC�RW{���xW���6o�|d����\BM_�������������)n��6,��X���ލ{�Q�P� l�j�!���Phg搽�}�&O�9���H��'�����_��s6�����t��s#�x����w[��brq�	ƚ�E�:�T��g�fۂ��ok��d�Y�$'z6�ɟX.4��!�%1���3��/}���d��=���8uK#T��t�.x���˞777!F�$�1h�v�d�~%�!f���[\�KevƬ!�+$��)|�_�)��ϘX�w�����)���-e.�r�b5�z(�(oP�k����FgL�V��w���{�N��_�����Z�"�͔v���-�*������CefFB�����\H=��6����p��9������#�C����4Q��?�5��a �L���nڀ͡2�9KJ,ހȪ�x���i�����e�H"�,�T�����|���Rn����r�ihh�{o�BE�I7s�݈��]OpF�k�y�/� �񴧞Ǟ]۰���|s�30ũ�]�w�A).F'��O5;O� ��r?,�в���"���E!(��L���F?���^�S걔�8�A���R}���\<�n�-��l!:X*��,�i���J����>��R��A�Aʰ��ڎ�\~.��41MBN{�ܨ;?W���4q�*�8l��׻��X��N,@D�>�~��x��p��(�����{�((�D�x���S02N� G<�χ*�Dh���)����-m=}�@Ӹ�6��.#u�h�-�#�����#�壈��y�p�VԂ�"f.~��Yùi�]_d/�H�µ�Ƀ$Z+W�Bm�3��݈_��VSXh덈tݏ���*cׯ[���b<��7´8a8
hȵ���\�!��&&�nG���ć��rF`�]��-���a�sR\�"����\�hll��65#ls/yu�i��A[k�����,���V������;A��jK��w���1�-����S���-<�2������0d{L���熝��i�,�E��h]�k8a�|7�l��s�V~��k(�,��uGN��0c���]���=�p	�M��:�
�S�7l)�!#r{���?C������ޙ��o������R�*�=a�c)�|�g�c����;׆J�E6T�]��!���>X���{��;�������B^��NX��]��0��L��VDW�_�16���a�����*f^��o��o�Z�&� ��ҁ�����m�x �R)��m��gÚEcl���#@7%�T7oX����[�^6)QA�0fb��$��_�D*�F�Q-�����;��S�_b��)ͧ�Py=��_�._�#�����+����>_��7 �\c>����/=��6��t�o|�����v���}�FO�������5�J���&'j������+ڬ�6��D���x�C�����������s_�ʷ�3_ɾz#�r6'��0�u?��6LF{n9�壍Z^wpCc��� ���*ln�%�!���pʠH/VH�pM��ИtÃ�:Ɍbd���~x���bxl֪8�\W�}=xL�Y��I?@%�-�XN�-��8��
��T�dN�:s:p�.�䴲TlF���Vh:�ιo�!if{@*��t�E�P7Y���6�D8sF�7Z�Hǝ�Ns�F�Qbf$�"��=+��O��K�Ҝ���F�3��X0F�y�fy+�I� �;��|�"�6FMm~�ݻ��x����	e-"<��W�����:V:κ�@��{�z���q���b�uc��<���ڻ�;��2r�f$�&���s���rt����|��VF���a�\�M}�[�p����][n�bW�}�#ݨg}}�M+��G���VP1��'�G�*.���oyߣ�丄x���q�Y���q�ZQ���J��/,$�N���}� /�b�oiS3x�T�{V n�n�h�0�؟߄�8���W/H��qo�DO��7���7��յt���"�]8��OP���1����JL�ZPc��ƛt�	��s��h4�+&���r'�:L,#sx�\�Ն��*�!��/�GO�AnDRb��'�u��M�%*�r^�w1Fwb������!�Q7y�|�y�[<���w�fR� ܸ���m�/c�/�"L~2\/y+9�R�ז�&���봁H�r��0Z��Ӽ8����hn�t���β2���q�}|���I!)�����7`��} �;m;�=(k�;JQal������=?����u�3�ƻ���j��`#Z�&
]��\<T���܏��wOF�{��NK*���&W�*l
B�tw�=u��Ё۷ע��A`UI��ۜ�2��'�����2ٰ�a�ݣϝ�4#�k���]�!L�"x��y��>��$�9f\�!"-{%�y�161��>z	���31�Y{br}ܥ�I8���kw�6@d���}G0��;VwIC_w��������1+�E�bN�3řڟ"Y>7�t��׃�����r��U�Y�p��Y�:u�����N�����x��;����8Q�՘R'�3�Ł#_�m���H���b�����ifZSXle�p-��_��Ʋ���HrR�b~�c�\�};=���dQ��M-��-C����/����� ?�/�'�/.awV(�i�����O�7ҫ2����.�W}p�SD�'RM��
Z���殮��%5�m��ǚY���_g�����6@:�t��E�Efq����q<��8��Qx��aq������>�8�%�U]&�/�#e���Cy�����54������8SV��	>݌[yi<��y8T���{��?V�����(�N=)�c�l���&�&9ƻ�N:��ָy�e��,*cd二p�÷�_Yy��O�I���\�EqʕmInj)h��p���]@>ыR���Oz�_��µ�e-q�8r�]�X�Xit���l���˳��9A�ȥ�w�0��2�u��I$�B��0�ِj!�w!;�{�`�����*$���k�I"��"�\`�.��[jlQ�L���
{?
�
�IHj��Q)�O�L�s�'���K�&��Z�h$��0g!�n9\�KP��>�n��̶3oB���.Aa��.%
�H�[;�=�6{*�N���\\t>�K���[� 1޷ ��1��(q䢢���SIy�E`�Ǹ�jJ#ː7� �8��M��2�����9�|	T�BI��z琌�Ge��[��Cȯ�����D��R'���-_��ϟR/`�iي�Ŵ�ޱ�\��g��@�i��g�&��� �E�݀}�5�A]*I>FrZ�_�'a� j�YYM''~�E��Ps*g�u�:���L�����E��O��a!���i�Z�B�9�S�-BO�Dŉ�b�ʆH��U�-��'�ft�VŴ�G�}nkޞ�:������?�����)�-C��Ϩ�������T{�\W�r��S��:�<���K;ɸ��7���Ddh>����˝�Ǥ�:s�6O̬C��|E�qY�'����ya�:8��6��vq�A6Y�#�F|��`�5�a\m~�2}?淇�{�
��]x�'�����Z�)/�lL�����>ֆ�zA������֬cc#���(�D�SL�|#^89���^Q�$��6T�L���L��E��A-Q��.h)d�~0����q�p딿��P��y�(m�-�g�b�ق;�J����N��w�	d��b�
wQ�z5�*�Qی�^�Mf@{ݞ�}}�����Pt+l
l�wՉBn��jo 1+�.�Z�\��l3W����
��G�TH8��$���������P�D �M)��qUBޝ/�XY����f��Tx�/?�����S	�е)�_̏�⡫0+ZS(|��gXu��k�ހ��@]>,�@�T�aZM�$ $�\f�ַ_��'~ε�%�I�J��u���N��?X�ݛD,C"Z��ؘ�-0]��F��A`I��O	�.f	䢢��r�z0I��⺖��)���l���qŠ"��ղ����4�����g�.�W�r=�RΏ�H#�ꛈ6*d��<�R�u����xV�9J�BE$ۖ�v��A��ZԊ34dYK�vi�(�9�e��v~�Ѕ�N-�I�8�h؉�/Hxb(�?�s�z0��F���1�܋�PW�v��]��2!�3I�ʧ&���f�p�ݧ�ëI%8-�q�"]L:0���,~��X�T��F�C>\��L%�<���c"$��Xn�?#\q(*�Rҹ��A2¥7`f�j#�ezO�\r7N�m�l>/��&�WI-�V��c����&����t��ڒ[�����?jr��a�\�<�OLCn���,��!��R3�\��M��rC��r"��S��Y����\P�s��\��ǹ�F*��ܚ\�r��G��A�%���K��X��v�C����N|`�f��1Ҟ���L$�w�;'�����W�XH�<^RY�v���lSxۮ:l�j�	Okb*��i#�j�?~ǎ>��y�uE2��x�i�|!��:W��GN!1%:��~1>�ñ��$�����w+:cݨ�WND��3����j�S��W���1.�M5��*u�э�����x3.������`�f�Ǳ���\3���� �	� L�2���R�@g��7M*���<8+͈�|���⺕b����-�\,�N�7���%	'`�7C,�K"RzR���3yI�eZ�|A��q�	��tʕ���+�R�NJh���s8�`���E��@.�ዶ�1)
���>�#'���b��+���b'L8;�Ç�&+�K.�S��=4�5��d���{����y�4��P[����$f�(��	7z
�B����)a��Z�.�'\D"�	׭_�&�S��/N�R��r�ƫl�=�J-��qfd�3/%�N���/H��?��uZ�V�v�:a�����''0:�BM� ]���1�~n�т�3�d�;��+q�l/u�$���'��0V���J�HE�q���WI���?Sj�0~�*�}�4��q�괗W�F�l	�$p��ķ�q�a�C���B�)".n���-�pQ�Iu��׽)�	�a��u�#�� "P��_<"@0M�;�$��!�Hn�""�{���E7��AɅ���F!ߜx��t�K��D�r��e�2�ɍ��I������qy�Nk���sr󺍦�'��#�����罛[�;�W�bH�l}�D���_%�'?��JjyG�������G��4<��/�^/�eg����P��H%��mIE��W,��	1���o^1����(�Sqf�X��$�TV�� ���̰CִS��/r�EO>�'L\)Aa��2B��3A.Z�p{m��g"�F��E���A�������ۨdY�Q���S�����"D����eK�+9.�]�ht	3��Rq�%ou����1A�]�s�`�Sn`!�����j%Ċ�<���[i��޻'��mmI�wG3\�&��*�k���3g��u@���ٓ�sa�����iJ�b��R"K�g���j�]K� L/3����p�	H����qǾ0=���B��+���:��z��un:\�p�IR2n!�J#�Q�=����0w촔%<˛��⡄0RF˳e�K�I��Ӻ�ҡ%�{Q{4Í�͹紈���*{��X����Ӳ�ܬ1:�*8DS���-o0��*�+%S 3ʀ�f�U2*&��ԺH�}^|@���{�ċ��tm�
�i|����P冡H#/[�GY�V�>��)�{��V����hѹ���x�-��X�N����3�qxy7�:���o�� >��ڟ?}�z�3�>z�X�4N�&�^ɒw�� ˉ�ȧ��a���ya�PܴWxyy���"�2�d�6r&�� l�8	���*��,^2�m9|�=�-#qtU�d��pY�J��B$T����B��Br��FH���9oР���%�sD��_�N����J��
wjU_��J<�I|����
���]��8s��!פ�[g����h��m�o�3RC�q4[#��r[���>��NU�Q��:��Df�V������%�:�[XV����T�8,hD�v�����M�q�g���z9!ak\q�B�>�|c��$��`(�!:��0�:G��q����g9>�B�U�J!��4��#vH��Q0�<*b�Ȁ:��oƋ�b&�Y��>���W�����g�8.F�K%[����9�����[�-9%�M�����+��D�������d��!lߴ���J�ϕ�}C��+�jS}u���<��1��@�hMg��_ޮ���WKZe�";}��9'��$��`mW'Z�!�Va礡�#=��O�#>
#]S�����D�Ѩ�CU]Y����Ι��Y��ਸ���^�:�U����h�����'V�6�J�SYQ�۷I���{"1�ށ1�-��H��X7��$9�?]���q��(��q97o,����1����H��¾P�F#�s�FOh��Π��@��Y����ܴv�g�FƦq���[^�?^O$�Q7nX'%1t~�w���8Qq�"�IA�8����8s�u6�vH�|y����9�~�n^[*�E�q�Y���Htǿs�Ҟ��p	
EXc�6� �Y�J��+w�q�ΥmC��Jy�}y�}R��?�"^~ �$�S�"��Z\�V+N͹��.!E��{��7���چ���9!��q�������_|�w�qJ������� �����;Q�
:�Փ��o���	B��_�wmHr���z������ Fnل�~�j뚴���&f���7o�u�,�a�>2�
cCk���r�*�ëR��K�!ƒ��[�b!67��S��Vl�֪�֎�C7�/>�8fsN������^\�2�PV�2҈�c7���f�S��������Nܰ*�pfL[���َ?����uƈ������}�w#[��Y���o�����/���^�FMu>��[��m��5g���'�B����e!ʈ�G�q~��F�6-=��g���WӜHzɰ�w߳���D3���S���G*����ڸ���������xD�1�����'���Ӈ��bKO=q�.�P:d�p�-rMn�oxtX�P�͌K��<�j+i-G=#������֔6\�\佰QV�Ej%�K�Jpst!�˘N���'��6���s_��*pM�[����0�!fAޥ�2�Ƶ�^�y��M$�U�JL�]�_l�*�ƃ� )>)�嵸m[Z3���/m��F�6|���}||ݧ^�ڪ ���]�b�CeyL��SZ#�T�w�%D���p��"�\D�>�$gO`Sc��亵������oB�p;���'�#~��ܲk^9=�OU;/6�!�
�t J��q�l+;�XҏY�غ�ó�$�t;D|w�؂��P�,ȳ��FGk'Z�.����*Ϡjf� ���Nܲ�:<��sp���+p��iVOoA��]��=x��ASA�Z��q��� ��x�{ޅ����<�YkS��B�쁂<[�#x����/?���"�Ĉ��jP5�|���������I#Z�D/��a��j���/�����;n�È�|߳IE�����Id6�)	�$/�:݉��(��R:,^_�)g�:,�s�*�J���ֲ%�������1�CK]���^H�I���o>�×��*"^r�8kwJ��+r/��E��)W�(�%ω�P$���JÅ�����:��:46G@�A�2P^QQp��)�Cy8��;�U�("�q�{Yy�H����67a�a��QJ�|�[�)���N��*䆮�'�p������X^`�z!��PnZ�a�e1D�E��b��58s�6��`�tQnw�-ચ�o����&T���DS}L�]��j�0pm�ϣ��:�b^3�֎�����8�TQ^��nA��8۪rIS��p$�2cA7d�T�{󈲉X�.
L�x�FEL��/��V�h��������pv���Fס�(�A(��3��
�#�WZ	!+%���b��'X�����l�O��uH�-$�������^��	�R<-�h�1;js{-��H�SUUS
��LFB�0����]y��(�"�6!.������CӔjOP�f��K�b:Q@Q�WA!�!C=�V��\��(�p@ <��)�'>ȍ��f��u	����sn��b]̃Ş/�MN3��FRS�tF��Z��I���]γO�h�>^ܭ	r�H�eN��%D<����neDM�Gے����!�6y(Qe�6zޤQ��JԞum��qP�i�2F%�F���-�1F�N�d -a�i�s.�ʕ��ޜ{�w�Q�����y�VH{��P�h8"1�ԇ��l-DB׷�P$4��(7[X`�#��M��W�Wg�#x�HT06.]��24ٖ�":f1.m	����)�-�K
R���밦1���Q���4�`�g�
�^9��+W|��E����O �[��v�������@�%��|�w���y�s��c�p�(�;&<����(oQ�C�䩚2p6��<�3��|րX��/Σ�⼵i��b��7�o�Տ�xy�Y�,�>��e��\�ì>��O�u����u�R�P�y��D��tx�̳��V��R)��~)����0���E��<,ub~�je�i�j�-���>ue��S�#䠲�G��x�z���Z�SWw��;ڊˑw�=�D�,�(]�O}H ڄz� I��C �u|��b�1�{�;�`^6��Q���� ̯�f?�K�s�ա"X9�&B�$8A�br�U>5~�Qq�3�w禕�q�N�؃��08�t*��\��#g�'�x���Е�K�DK�!�㹜AWW~��o�͕/�2�q�^y.F�r����᱃�x��ǸC��d�z�p-�l6C���cty�i-(�L�ԁ|�Dy���t"�Y�l��Om<���'!u�M�.������@���yZ�6E�ay��fW�|�|�f����r�L��eo�4�9W��'/�l"d\�;�:����y�[))f)CfB%��� ���X��¦QϦ�&I���q�I�\*�)_T���xN��^!���]�� �E��8�
\�����:o	�������U�J����.$X�&8��s^1i�S�P��������[��y��g�J�t����q{���;ނ����W^ \eu�e�-���hoǟ����`?*D��'���v�
6ܱ��n<��\���4s��Mzy�8q:��7�Ə-���,��d��4J������EN���~�I�P�)y�,
�.G/�LJp��j�ѹ�9�R*�đS1���^Q���듔�v&���3�0�(�ey8���,KQLQm��E�Љ���hYM$l�//�ӧ��Ҝ���2�_5�2o�J:q5A}8���$\=el�~��tȭ�̙�87��)��>�ZUpY�Pz�ѱa쿲�����<��i��+�  ��IDAT�g�"U@e|�u!�+�܈�D��(�SHH%�AlJ�+\1���4I$eS�tB�U�`�BՕ���~�J�j��*	������~4�~C<�.Ą�:�ứ�?p�gj')��G�/u�A�hi�DKdjmm�o?p�3�C��$PD�X-�j�&!�v|�<���w!Ʉ�g�Ϲ�iށ��n�h,!$d�l� X�Kz���q-�l���g�YC��VJ%��Oo.�$uYM���l]�W�"fzqq��tcjA�!Ӓ��]�R�����x�s��IL̋>%󸫫^>��+�c}$�u�t7F��«-�q��*	���>l9v�,g\IN��<�qw7'e��/�����}ⶲ��77�M��:�`�(Ԕ����}�%Z�bi��ެ��8qz����~�3��ޢN�`}(�>�:�������s�_��v8�$^�`1Iee;:��QF׶�
����ܕQ���}C��)���J�]�ĈfH�~��u�3����_s�i���cI3.�g�`��"�aE�����%��c�u�����K>ȥb���>����3��wo�_$f��7PLuU4-aZk��>�q�U�B*����u�C�q�2��ZA��W`�^�߫���۶�hw5	Zp!ǍAu�_�2��ɛ�Y�K#�BN+��7(�i�E3>1��zp�fD��/����IV��{l�@�b�DܶX~��J)~ʷU�1nD"W�6JCAy�l.���|��9�	]6'�L�#L1[�"��r�<��o
�D:)�1"�F�		�a�\]��5��nP�b1�'��z��ԫ�&NI�'CY.���Zw�u�R��!�<��VV�?,�i�=�3E,C��S�"OL�C��
OS�j$�"�9�d(�\��q�)E("�07hU�����%X��RQn��#����Y�qP�LL��nU�b���y[���ۂ=�2젩���*
h�L:���.�Y��i�gWq�d�K�͛6���1�[��e1NhڢW�����J���a\ey����ǒ~���W�I�6�;J~/����D��R�뮝h�^p��� ��W`VPH>!��F^B��9�1�aK����-�̿@_�œ;_��n݆ݭ��̻��эFl�/1�O��5���s�K��l�����[�'�?&8��p)>\BS��!\�f����0i���a�>w���o�	�@�n�����bl�/{ê�u���걐1��F��f�~���N���r�Ѽ�X77�~'�^���>���(Wf��Z�pl|��q��VDP�~�t?��4�߄3������P�q�$�
)Ű:�F���\�����o)��Z�3��u�wE���H�q+Q������l�m�Y���!X����tu�Am:��*g\I�b�ѭ��݄$B��X��2qI�"#F�$��u�QcEH�,Ϭ���,OE�̒~�L���}�Ǥ�+���t��`k[օX;C��~��`J�YH�;���k׮3d��� R����^�҆�sDɁ��q��{�k�n� ���=��↶I&��:B�a���:̎�o�����cS�n̬����X�[oG�ʍ�,�c~�����jl޸�-a;vtM���
}?���Pva���KPs�bE'n]È^B02f�&���CF6x�լC�i7�����|��M	|o�\��%�s�2��X�r�O�
�-����o���$*F7|�#�ᛊ���wn��#W�NU��Ʊ�'��Ǳ~m��̹�c����aQ���<�o<<�^����H�18'���gu�x�~��b��Iͺ�¥>޶��~��g�?i������P��(aDL$ٜ_��sR�F����GR$���l�s�H�b�q��Ϊ�Eun(�c۶]H���j���	g�|��]Vg�8�M�vb>_)8(,��a�3��b}^�#(Զ��DuDY����
�`��Uka���y�F5�Y�PW�'9�j�����A�1��QݼOrAz�U+Y=9�$�|k�%���hlu�)TMͭ���&>$�v�>f�	MߢqR��"r���ÿB��(�ÆT��a����G&�G+V{�����P��Xr�Enf�&s�{���\3��
��S��yM|�A󢧺x���K�H����k�vD;�D�������%|��������m-���im_ߊ�8[�2�b�������X�ɹ-�k ᰚ�@�(�mϥ^G4�CƸKH�.d�٤�ĀW�	DH�O:_��'����9\�8WP��l��6�����%����ܢ_����UY� N¶Fp��CxĻ���Nu�
EP_݌Ji�P��N3��[���j��E�'�Hm�J�-h��џ��3�*�q#���(7���5�HN��x��v�иU3��
��5�h2ƍ��bږ46�Q���NN�H,��b��8�IrNԇ�4�[��<U��|}�(n�����F���"]��9�HsM����T���V�/a:5�F�m��qu��#��Fe%�t]�E���Hz����N䡽\5�!�S�?k[4uE���R�J�����ȹєA dP�כv�d��i�%����%���KѢ����e��2���%���hD�%B1��
)�.:郤�4�﹛S�6yab��[(k:uCBv5�?Kk9��@b
etDpңݰ!O������0.�kk	G�Չ�RlS�p�m��&Qd;,��6J�$���)GyBB"b�9�A�=T�HH�8�-� ��H�h\���y�q[� 
K4�����ϋ�B����#0����;�EE���t��&�����f�O���u��;&[�J����1b��}�*�V�N��Ύ����?0���.�<R&m+|��͓���:�8���(ִc,�ӵ2�l��w_c�#V�R)T�.���q��U�W��D� ԫ�(Mc#hq�I ��y�a����������T����
x�K�6�{;�ϓm����H��$�Oa�����E�i1n.��WK%Bt=ܓ`�&���S�(CQkÌ+�����XY���0�3ˈ\�ד5�<s��M�z*���+�����طrZ�s��F"*�
���ZʗڦC׌�M���8{ce�0+�2ɸtzq''��Ȱn���8|�3eg���܈��a\��cy��o&��p��8+��dy�be��1��\�ec �&lLz�l�e1���T��t?Ǔ�Y��+3�r��#��4SC�]J�R+Qه�S���p��[]�c^����K|/��cݩ�C�F��2��${�ڈP6ֆkM�&Z�#�Hm�@��e��#T������3�Ov��D�&���0(�S�3���K�8��y$S�'����W�P��#��0�n���t켧�`�Sf�z��4$݃{�:|�\���xƑC��Ր��)�qFd|K����}{����rrYvb�?�/<��;������?�����s�� ��R��_[V���y��T�o.+٨���5���o�<����2 p���!���c��L��_����w��ɣ'�1��6!1)L6������X�
CP�Y��T�F���GK�Ẏ.�ד	R���N:�L�ZƉ^T��F��~�N�1.Ɯg(��} �rۜ?s
�Z��n�JN��F(�/9y�oܒ1}��,�5-�h][�dŭ����^y�n������1��|��N���W�E(1_r��hnnŇ�h���:$�&fS|���N\�O�?�OMW|���d�=[�q��Y4��([3��>�_NoÁ/r��c��7����8��B�HAm@��xD괨�>�ʍ	,&�+����@,Qe�ò�J��F��R�/� �Y�����W��\~[~�F�2����H�-M�e
tQ��lij@���� H�k�����Kx���甫Hq8,�]"B��^=�y�O$�J�X�+���{��+H�W��,��G�ʣ0˛�zG�������=�|O�o��O�H��JlDK��ӧO���[��Ўhf�1�H�B�;���<������,s�{���U�{<�|��E���U���܊\?�D�����
3~���q&RLbͺ-Pquw ��qh������"F"B�,քAU,��}3Ν;���q�"L$%7(�#�*;���iI]�Bg�U�&C�%CO]�E�X�]�����3$� ��MM-hmm]w噝ג���:V�7�>5���;l�9�	����.8��*��6�ꌩy�i5t�枀)�<�H!�>�Ri8���-�b�"�=
A�XM\�9�'&���[YG$�� 3� ��`���d'�Rx�&!�ѾO��G�m��������H��
k�k���q\�tK�w���R�_�4(����b�'ޅ�̃|کI��b~`o`	t*MT܁��䲊SSN�@�E�a���U���e7J��v�4� +�DM�(/�Bj��Ѵ��^�^�=������z�DB6�*e���1�����c�`�e��ѐ�`�,���7�^[�Y����7��^�z\ǘ~��� ��k�	w�@,5�P`�K\���<{	���Ǝ�
��Ɗ����+Xy߳�7���>��P��Ͻ�~�ڛI��y`T^����oĕ�N����_��&F4K5���;�6�;=��7��`cGUr�d�:��E� �0Y�&|㱃��sY��)�/_��O������Ć�Y�7E̭���3�j�J������d���*6��h��:��R(�<���d�n(9����zȠ��0�ù�2 ��2l��X�+Z�C�HH]���>��O�U�K���r��un��M�����+����r�e'z��`qP�	���o\�&W	2==�?�ۧ�� b�d\�&ǟ���/�)��c�3�g���m
c籱��>�Ғvri8������H{�:����b�p�r���>t[-���c�Q"ćIc��� �G'�����p{(
>u�2��Y��M���&� �s,�FZ��Hzq�����.�aʅ�H���T�sA��+a�QV��pBuA*�E�~�e�4���WL�-O*nE�91ܗ�pY�BT�q�U�J���3OE�d�Uz����ڧ[n�����3Oi��u�����G�w�ii���I�P�a~��DB������t#�`P�������"��	�O�Ni��Hv8,�F�[�Π�J��S?8�@�D���F�i-�AF�ɪ�qi�?sO��-o���X�,	M��Y.)�>�R�r� ��x9>���pˎT����C�h�=�"{�LN*�K�.��r v��\.,8�6E�:UD�T��FdJ�K�|��Jx�C���.���\��㱣�w!�u�k#�?[�����o)�p|=um?mjnnq��J�������,!��� W�d�x�k�x��)|�� ���:,I�q"���K�Y���������?��7Ԣi�N��vW��3���(��u�cY�V�'���i�u�,Ϲ�o*�����wEs)Ⳝ������5#�,j���	�� �Xy+��:�82%}W�^�.~+�O��dy�ڲ>�S��y���Mˑ���������2="��*+	C
���:�����+\sDWA�b޼����"�<�C�		��]�x�%�^z���˾r���]C*��w!c�:⾇���O�59��,�H�"^K^�K�콫�f�q�(@>�W��b.ʔ�
&�+`57[@�$�	a��FgIKqR�/D�'[@�ƿ_�֫I�Foۻ�I�m)�522�K�.:�m��5��?�:���F8Q^�,�%����b�$�{�G9RR_S�m��R���������mO�:��VB��:_��?F�S����LW�%8-��/%�УT݆�_C�!�C�e�=3_�ҥ;�Ǚec�P���`�y�gq�$�����B�)1�l��<&]{�	�MfVUe�G�B��I���YEY�d<�%���Iz���K�z��/~�Vu���OL(�#�Qq�Bʂ_k=\1���������m�=׷@�0����f�K����䙋��厛��7u�����ܗ�8�ҡW���"aX,u��T肶��¨��¤�|�V���K�{�XZ�x���*(����R��b|r�,��0��/ 4���ueN!�8<Gw�i��
'��� ֚'�?��L��:��'o�9�H$	&��(�I�,Y�mɾ��%���ڟﻖ���}��g˖%K�m%�%�b3E� A�� ��l�.6���ݯbwuO��, ���NwWuuuթsN��4M�ָ���NԔQ�� &�t�eȹ�*��\���wE���a*���R�G�ò��D���QQC�{�A�TX�{k\�(��CJIM�����_?��0�5�}&yA������ڌO�GGy&�l��8�՘���7�C"aa�܅�:���D��Wތ��y�bWW<��� .��Db�����*��&
��<�R^�r��5��j<�S��]�si1y˿����=�G��t:�'��J4i�����9m�ݡ�غ��l��)�ؿ/�׶a�d�8�~����٭B�����]�JAV,���M���i����a�f�9J�م��Gd
���]Ҏ��9��"�H3�{�frA�T*�NT���;�š����\GD���p-��|ב�}�#/�B).]���@j�,ݯ�9m1[s�p�S݌r�W���,�Q��gW�V5��y��3R	�x���)Ͱ����<e-�_Ǫ��{�`:Ӊۈ&�Z�)�zMl��*^��m��@��j`W)h<ǜ�2Bgi�qQ�,�)m��zDµh�;*���°�Ge��~?�q����~�@��7Kg��T�.�m�ORua�3��*�8gy�k�nwI$w�E(�2���c���]�2o{�(�s�.��)�d��Qr�-F^�������*D�e�+�ǋS�Q��|��;h�0,M�+��"ʫ%2Y��yGQ����bp0F� �O�*�Z@쒄\}i�NK\�+6ex��5n��@2պpH�Ȱ.(]X�%�g�WB����I�&�4N�#��(�)�k�1�	>���@c`s4�����1��ڸ�j����˃��AW&ei�L~��}�J�cV�-�$/�����tU
�+�`�Jٶ(�XX�,8�k�$����,�Æ�v&Lw���f�>\\B���8���遭�R%�����\��ŸJy�,��yR0;��ӢcA���8�#eye3u睵�u�aL~�E��	�rp�`;� �O��/��\$w=���Y�������\�HW��Y��8s�-��Z��dzo)%�\壔�P�e�^�+n��jY����T?5�����"@�Q|m�ڠ/���n��"�Wt!��E�;�_�*�"�_���L'�8�[M����S�/��*4�����ӖV�U��=�����#�|KGX���M���$�����]^^���:֮��F=zD���J��y�����ݹyڣ�:���L5��gΟ��d4I��/��a4cN��N��=Yq̩Ӝa|��+L�J�a�$�0�9LQ�`�R��r��}J�b��6�f�����XNE�A�c�1��Z�҈��֥	�-[�\Pc����3��~B�#��h7��y��K���Tu�)Ǔ]��Ƹ�M�Is��Y�����466bxx��RP�G�G�H�F�aJ�ν0���#q��ӟµk������ �`%2��x`[}�x�W����۳4�_�%�u����M݈�<)��%u����R
r�(��u��g�����xZN�0��fA��K����q)�W�;�%�P�/l���p�}��'{ �ng�(v���{<�'�r8�O�{Q��Q�./�|�p4��%;��m�ȣBs|N�LHF���5��3��ZZ�oMӋ+:v9M�
�{���U�}n�QQ^�2;��������u�(�ڃp�,�?�D��!��G��(�c5K���PRK�=�\��_��
��=��̯ �&��+�P܈m;c|bB���At�)�b~�(¹QnOR���H@E�_���a�';���Y���3����7��_\��� ��r�qU(������+�b��ҥ�)�$)/����5�hοʣ�T�tG2�K�K�*y��:wi��n��]�ocu����Ӎh��R(�x�H^ը�Lbe�4^�;���3l&aa�%K��=�V�Cl���4**B���o��S��&�ϱ�f�cXa�?��.��X,��k�1�0?�$��y�>B��G��B���Q<�u�,覰���
#�T�i��tWo����F̋?mc	��c'����b�����U�����2�s��l'^�;��gj�:g�*U����� v;\�)���;vp���KSI�
��2ݼ%.QilP����z`f=�"�?�+�r������W��Ši��G���/�c՜Fq��cM��!zxx �DK�]�N��9<���1�]���e���Y��啘�9;C��ak>�	���g���b
��KE!�(}���6��BU6t^LK��y��ټ_�D:r��q����6���8c�m~�L�h�8n���_�z� �n�.�e�C�7��>
tM4�������4F��!��x��.ӭKe���ag�%1�e �� ���C��"A͖ e��"�z_�\��z��e/*f3��h���_{oĢy��
0X�&�Ï�L!�1hs�� ��߳���aI�\������e����'Q6ݯ�
��ZE�ʕ�z�>U�q���<��ˇҘm���6-)eQ�_���1w�ϝvEj[��l�`��@r���J3&P�\ӈ��������#E1d۰�F\~�,�Y�E�>�#��)d%h*q�\"�5,��T�i܁�4��3.����6dR10x��������b��m|T	�~F#LF�$Y~������U��L�Tg���syT�x�����f|�+��*n���e���J�cٯ!��a���q}�#ux��0O[3Ւ3L�Z�mSN�E*]E�~�ŰX�-W��_ ��ϐ�{�k����W৏��$[�i��$N�"Ǣe��ۉmWZûM�C�pFI���Bn����r��|wћJLOW�"q�>8����w�p(4ץ�q1�P�6R뤯�U�\�)����E��6�__]���^[%�	��6�5�[�@�k���o���1�K�"���<�klV/���Åu�����ߊP�U�/���=@f!���7A<�ͻ��&��z�����o�*��QM�줖�����?�������G]���Kf��z�B���(�<M���* ��4���Ez���8�Z�J$��'�L2�B�0�й��]m�����^Wl��E�u��&<��D�f�m3�X���ڥ�,�,����>v�M�z�ل*�i�ה!D���Y6
�^�A�������P�����0-���4��R�d�̝L-�sJP0E�M��pb�ݥ;����B�(243&C_n�.#UB;S�('s6ej'W9�T|R4���.�=��4ƕ��YІ�wN=_
LL�z�o�\!;�J~�T��W��sN�4V!�� Z�����w�`B�nq1�H�j����S�i-Z-T1�U.u6+61Y���1�k�?�ibb�1��g�ett��i��)���+Iݧ���T�Ib��F�A)���0HƄl�wz�#5r��0˪��>\bG�͊��Q�O	��(h}�43�Ҕ�V��J��ɗ�����c�rϡ��j���t����j[U㻖wȿ&�6�#�j���ҳ�HM�d�Ř�irϢ�(�x�
^oѐ�\\���h�d���]�ɤ�����6bqC��>�$:�j��˯���f�u:*�c|bk�ݏE�4��Q)�ë��	s���t2���۩R��L�L�qk��"/Gm\�-B�N�)4,���yqI�hCn,���؇��bC.��Qj�ٞ4k�L�Ғ���m�A+�#輦����p�t,#Mx�0�Qnԝ=��l�d�5�"lC8{�߬�)��^S��l��0���<��Nar"+H(G�����w�u���O"ՌOG2����;�rN�?��C���,����0��k͜��P�eː�4n��	5��p�R���C��JL��L��qɬ'�;u��ji�8m
m�b�3N3?�"��Mť-)i�7���N�B�5���8V�\���ϵ�oy�WMs�>~�(Nu�N��p^D��R��V*꞉a��9���B420�O�$��T���p�޶�fK%g�޵� �o�	��L�8��#"L��ͩ9��t[3���&S��we��.p@p8����%��=W8-R;Y�~�=;�A�9��#,x:-~��4_���Cs#~�+�:?8Ћ���O=|�>�+���I2E�a��m�)3N�+�IC�H�
3.e���²��aɐ�m��.��?�����s�W�Ϝ�ß�������E��)�d*�tmRU�B~Z�F'qv�Bs�UϜ|�� ��En�yh6�l�6���c��a�����ŧ�E:e O���_/�@8ͷ,ӄ1'l\�z!��r�;��r\#r�zJ����v'?�\ee�%�]�s's�Qb,�A2:u%3p�������h������T�}���h�r$<��ꮦ��S���"�_4�}˕O�7�٣4e�:�.�-�uhmi@4�C�ۘ�5�P�ұ���Q�pMM-y�c���>,m�`N�|�d1��˲1�"V,����26vV)c�0âu�e�ʁ8� �}�H$��Ϲ�p�;F5/���7��@9xm'N�li�4�~�)��6Wg�Ҽ��z^b-�@�'�`d%ц�o�?<�,N�>���<c�뾘�W������# v�B�&0�d���~�.��I���V�.	�u&�sHs$MB夎�|��d��� �,��F��M��;O�H�q/up�:�M�X�F �\$U���*ǟ~a���jqĭwp�jDJ�C"1�ݻw24�b��~�UhmmG�ً��O�����i��߂o>�g�;Ӳ��)�)�t�����Ź�sd�T�8�c�t��¥s#�7���S[��y�ްSm]Ԟ{$�o��'�*�nȩ(4�{FY,e��~�"_�����Y��f���&����bX�9�vy�G��3�S��e;��bqT�m	H%ԕ<(�L+H�u��\`~���� �iŁ���Ĭ,�s�~ZlgR�ͻ�H��K[�~�s������d"�<t�J�b�\�iK!��&�z�D��;�ϟS[/�<@&p���<囚��p������)PX�pPC�io)�TXJ�*Yʃ�q-�U�q�n<�?}` �{>vY�s�HU�����d����c��dW��i�U�h�[��z�������r��f�N��(]l(|y�Y3��l��������I�Q*���q���mo�g�׭����/���ToǏ~� ��t���G ��|5~��՘�Zǲ�З
Xزc ��:�=��s�r�6ዟ���[�d2BjN���W�f���Cbj<lG`�WTV�w|7o����g�ʬ����ތ�G�x�q�R讧&`�Y�W��h��L�CG�q�MX|R� �L����Y:�0Ș�����/��Hy�A�A���KHW��G&o��qIQc!��ik��q
�D�PP ��p6��p3Վ%��֤)����#`d���?9����e�E#��&�l�9{X[�mC���>���n�*�)�i���Y�J��9w�+/����+�T7K�5�ה#���9��{H���Q��
��:n�8�hz��	��+qF��IG��'1�?���6�rY�Z.��*�4���;��P؀p$�p�����&ֶ��ｻq5�����Z���/�cv%&v�X1�+��e�S�9�
k%aZq#�G^ێHk��[1'�º��pKk�lX̙�`��;Ip���E��}+c���ڙ�L��#�\�6�×���7�&�;E�Q\oGo�4�A>�i��Bi�敨
b��i���9�xR�7~1A���/����TTT`<[��m��N���?�9�%�  )�F�5��;m7:��%�ݻw���%���J�?έ�;��.Z���`51��S��r5ʚ�c;�g_D��shnn�{��7Nj�X�P���*�ډ�ث�M�M���h���r���X���@nf��.����?^�ӓm��-�~�tT�:K;~-��:�ϯ!�
�~�9�6Vq���ci��A5'���ɘ�.�.�?|�ĳSd�u0�=�Yp'r58����6)�~K�d2�L5�Z�����!δ���.�Fm�T���+�s�Q�1��?�����<-e4�!�F���qL:����� �Nr���l���\��Bj��
���m�S�c@�PQvP��LMMyjp�zjW���e�2s�bc��迃��ٿ��k�URy8�lU�bQ���e�D�uoX�ò-�q݌�:�s�Sc����ۃ%�M۫����ێx�>x
�O!�(&Z��X@Hn@H�������d_9:>���^�tF���3o�S�޽�����Ÿ�����s��Rd#t|���֖kL5���1�E[i$�%2GA����,5µCW�J���z�'�5��&���M�vc�E�Uռ.��~�(���Y`���r)D'HVRӵ�(���^��ͮ�N�T�*/��)��x��դh�k&:Z���9r1n�=�"е��Ea����s���Gȳ�J�c̴�_dj���@gk�y��dX��^ ���
1:��#��y:�xiM���Y��Ib�ϖ�PpG�&�J7b"���f�x�1	@���^�����>9��wă|w�5w�v&��%,��R[��OM̋���ظ��s+B�](�"��Nu���u)�s��b
�������`Vn>T�)��xg��Э��B2>�f��k�|T
Z�7Q���!���x*�,�7�ZyΆ�����C�/e��yм}����� �?x|^m0&u��:�:
�[�2��'�N ����$�jvq5��1���ȝp:�e������`���ɗ~�J(��;ֹ�E9�gW�(�bU1�f�e�ɻaQK
���^.y�T-��.QT��۲���Jf��vV����+�.��JAKVf�VY6#c�X0�y��AhY�śד��s��'���Y|\}u�t�q��H�"DLLe=��<i�����M���EUM��νM�l]��D�}{u�jL����a��}/�R�n��r�Hl,7�Y2,�Z�wis���%D7j,v��E
�i�S������ F �d�%�S���M�ei�lZJ�E�4M�m]�SC|n��`M�!���S8AFҮ%�Js���0�i�n'�QA�cy�>��i�gq��]�\ �ȸ��c��t2�K�B҂2�uԋ�37/��.EU$�q}���EV�d��o��uVΥ�@SE5�!�I<��?�eLM�:��
p$,>�u���^!E������ku���0,��W�d�J�O3{����z�V�
]A�����m����{��#PE>��S��S�pB�R��d1�9����2UG��2H�zFx]�T'�h�P
&��m->��Y�pWR+.|����Hט�貣�T�i��ހ߸��8������7�` ���6?��C�S�gy�x#�#lS�3���0l	�2]����VN&��j~.��w�TD+�fN!fY�չ�2~�,����K%f�f�9�Dxj��P����8ԇܥ�x��H��>w�p��W�)҃�����(K��,d ����:��%ð��w���E�y~����?�\.�;*�HT�cD_�g_�j���b0�� �*+�i�2T�GPS1��=�@�AsHC6҆�������lh#�O9�Ջ��	��Yv?�R=^����-L磢�g��JQCTI@c��)ߡ�s�LK�&���4�`��Hǂ��8X;�!om�ױ��8*�	�ҟL�a�!���9j1s[X�;�8^8ͽ��bKa��Lu:T�i���|VT|���w����d)�h�4���;ș��\�/���i��1l}��tw�	��L@҃����|�)�`%�F��;���;�m��H�R�+���=�޻nFk�2*��@����^|�	���̇��i�)�
�a��9XL!8:�x�/�{�܍�ߦ�L�,mX�9�<�W��V���(���\}'�a낋M����JI#㇜ο��}bY�&�����!���v����>f�{H)�U#�5����Q5N��E�o ȬT^F��+UB6v���>V�?�*6Nl����e�6S�J�{�T��RǱښj�ooDyY��\����TR���{@!��B�P?�ǟ}M���j;�3����)�ӿ?��ѹ/��"�ͪ!�J�?~�����Uz�h��Y3�7w�e������0���{2{U���v]d�I@��Yf�_Z�d!�\>��,FbW!�s Ĉ1�
R���8z���p��y��,C�^�L��գ.�����Ç\Ђysp��$�!��M�L��L�鷱�+���d�lmDJ�}C����nD*�j��K���S�[�ߵ{�2����ve+�Ҷ+��b��M����l��GR���	�]5����0F�:	j2����x�5B�(n�z!�U�a4���<�lU�]d�����-��z �j!V7#h�p�����co�{?�f�Â�Fo9���s���0.|�8���5L;(�2��N�����
�1��;�5�"CE~����F�=�۩���f�^]+e{��j�d��"0��P����p��	L�LLNN�E�'D��ųd0'uBSf�ri�[U��V�ACdRH!e�F�`��^��oo�s������9���{W�ِ�.a��0�J<x������B�mf'�Le���Ev� �܅���d���L@�˗7㞍	d��묾	Y�3��l'�2���}�.ɒ��%�^���<@�d9N�2� $e��h�ıs(e?��󲥋p�U�8QC�4��As�q��p��m�|���ބ{.K�:Z��U�0�T����ɓ�f���wȵ�m멭��-�U`n$F�\���V&@V�S��`baZ{�~�Q]U���Vbi$�ӕk0��~޶�8�L5���>Y[{+��<��F�MʌE��e��:��x[�"VQ�u�u���8�#��Wy�]�1���1�+�>n1�7i��Ǫk]����$z�ڱ��;}�c�9��;����k�8Q�v�T��
�YT��P�0��]��&a�ڴGm������Q0�a��b�b�u�M�믹߼M8��*�9�t>�X�Cõ�}:��w�A���|����RILKeX�������í�Ϡ%2 =�E��l�%���&�[�������L���F�M#[iy���u�:Ϝf3pL�z��*%[)�G;��SR�
����M�_�%����ę�.�f��I`E��J2�̩D(;�򻩹��K�e?������g�������!Z.Wt��u����<�JbM����*�ٙ��v��>ET����7��+����#T�]sc��;~y��4��8J{ٗߤSm���9�ك?��1�nI�,la���A�$���'�L���[���GE,����������2�L�%G2,[��Ԕ/}�>ܺ�����5�75W����ر�*|�!���0�Y�'$��%�������~me��ޢ�Ra����~T����M����d%���k��T�ґ6����d���AJ�{������:�����'���,�uN���P*���P�T0�2���1;�G�-2"+o��_>Yu�}���Ðd9]����dR��C��J�NM���V͹���L�ߚ���\�*]�"ɔ;��Yd������	�)����� ]�5ӄ��]@fP�w�\��!�O�0Լ�ȹ��*�g���L�ڥ��^��c�D�(:O�wRUĢed)�}�4#���H?��<�r��'V1xe���q���J�\�d��.�������يH�
���X$����A�>���{�`��0m3�����߁ϬD4~ԾB+kA��rh�j"��a��9~�n��ȋ��?�
����t:��]<C��1�<E�IIt��̊�h`���ZN,�<؄�*�刍K�1gcc�s�r�9�J%<��L1�� �-�a��"�Ό�A��	�59y���dx�8��$#�&HZ\j01E��,�⩅��Q,5�0>1��P���j%t0m�I�S������ʢ�_Δ̆1I�3g�CH���1��]P$[��4Q�SL�u�2��c�Q���i�Xr�=}�*�0��\^���͎sG`�¾�2�v1?AMm�w�K{OW,����I6�&�
�9�tL�~t��%��-!�Vǎw�D�(Q5�p�7�/�8c�9H[
S�sE�9�<0����7_��6o#�Ӷ�K�W�A�5�����0���H'�867���7n�C����zԗl�j���ƥ���r
�]��O�.�E\s����#s�a�;�=����j�*�޵��A)��\�ͳ&Z= c�C�) >7�G'3�'}*W�>U�\%/�y�Fs�I�^v�J�-̴�}��`'��16��bØ�ᵩ�S&�AWO'&3e��)Bʴ�2j����;��s<�}�AV�,�Ĝ*zb��Sf�?Ї�g�@s
 ��q�g�ѝ�2�דE$b�կ��jPW�Q���F	��i��.<0x'��PY;Lt��|;�������5�D}���J�W�>iQ��2���Vaa��H�����}��2�䝧10p��v�&ʨh2�X�A���s���n����r�ɿ�ÉSg�=�V���\ch�*�6ጯ�������:n�_��گ��`_Z�qdNmA��Ϙ�����y�Z��z#���0
�*�455���}N���[�G���\�zE;"��� ����c5� V-Y�d��|��R�<��L�
��� c��߬K��79#b��NIY�R`b �M{ZƤ.�t7j%�$'R�q�O]����T(㒎�U�g�!�Aw[��o
�C=�'3�yT)�A ��&K�ɷ������N��l�'`�0l�Le��.^fc����PF3ݖyX3y&#-�E$�I�L���3�Vg�k���i��t�����8/f��$*s`
�&䷔M�2ãgYm�}�XR��X���i0N���|�2�B�!���QMI�R�<��p�a�E��,�9���h��Q�FuA��d1Z#{w��C%1�y����$�9������Q�3�oN^)V!M�'Őt%;��o���MU:V4L@�qƧ�,C��/�kwE��?s�(�#A�M;�O~�|����l<��N��Xi�"�l�D/k�cX���u܈��`%ϲݢ�C�D�lh˲�kq
U��rj��1�}�R��8�b��x΄�ٝլ<*J��>���On����ǂ<��}��	h6j��Em�w�m��� ��39�vMX#��P�g����L��L�
H��9��P�Z���a���E�i�#C�����:��J���:"�53�PʑU���ى�5'zA�o
�2���XY'y���q'Sx]m=Z­v���z0���W�S��m[s���`(/D��ѕ���$��q(�TQI%��*�w~h�_Z8YH�A�VTb�͟aw��l��R�J���6���s��� Y,�2��(5��^�$�APp��>r"�d�KbY|U�|���#+�l3�H���ҥ�t5YM���J!�i��A��͵��(++�cZ�<gX��iR��ꊵ[��t)�	�E�� �FY���2]�H�ý�=��_Ź!�S���d6j
�l���-OJԥd��5�	����	�2}>�A+�F�X�r%�A�eO!����#�[g�h���Ȇ�݁B��';�t��g�e)�[�x	�#+�os
���&��)�X�h1"kE�iTM����$�Xl&�g�����^a_�<݃ѩ|�!u����e�kl��sJ��c�	MZ[[�n�,c�11����d-j����PȊ�b�:�&���>�����͗Z|]z4;��}�ol��CTS	����&"���h���ˉ�S+��,X��%�M�܍�^b���:��`e�%Ru�m�0���Hm�L�j�Aښ���$8K�?�3�AWY���	+'w��g���`��3Loۥ����B��u�a��@��J}�JKː�Z�q���Ǥ&K�Y�e,!�I�+���"�m�R�(X�/�� \?�9} ~�u���%�Yey�0�v�P�n��G��-:ɝ��#0��n������	n9���D��˽�2�K�ɊU�D#�y�o$��@j9MTǉ�sy�s%�tGZ?*�O�ٲK�6l+�k�[Q�]�8̤]	�ȅ]iC�,x3��s1��+�a��6�[�*�m\��KE`��vUeK�y@0-�"����4��nob(�F�VAx�a�?Dh��V=�X.��Vu������Q�bs����g0+����L�g�S��z�L���jRo;e���,���%Yp"�������nDs<��:�Fs�0����i�|���^Dr�L�,�Ĳ��N-���oT���gw���L��H^�3����Sɳ;�Pe2N���bF�x�!H�o�~��]�9�<������˃`V��J˹��!��s����Cy���p6����U�F�������&���.tv�Q������i�����s(*e��N���e�����mN���8*�i����,F4{������n�3�Q�+���`%x\���}�(Ξ=�|�b*GU�*auu5�|�f�[����{xS)gߩ4���7q��	��C?UU5����cc�(D��� M���
|��8r�S�s���*��������&Zk�=�ұ�Q|��X?�"+P��(��+��7�As�|�f*=�� evb��^� ��ͤ*��%7�P���LK�N9���Z��r�E��$U7���&BȜ�/j�mg�2���(HT��2DU��<R���v�DB�ڔ;P�n��mЅ�����\�ʖd,տN<aMjj�J-��_\"vO����QI3�+�Sڢ��}�9ҏJV���%�<�Rޡ0�QD:�Ï�ه��1�U5cX�LG(\�s)�Y~����tæ��8��}�&�]�&�+|�+M����u|��H�$��Ũ���d��Y��M렗��Kfff���M�W{���E���[�g�.��v\].�N� ��oY�*�:K�#}�?�;�}lL��wz�X&��ՔO��,̟��V|r�I�+2�dsu9��y����"�!o�v=�[~
Ѥ0
҇ˍ`C����m��_>�v���u�5��K�M�]����p9�������K]]�b	��*�d�u&b-h������chd�͂۫Z�mW�=3'�>�漩����:����𨻈���&L���D^ /�4�4j��ߞ����w�H$��>C>����14��d2E&w��P����8�Ϯ1?�T�H��e��U㙳D�"��߄'C(�]�٭<��C ��e�kˣ!,l�!�BeQ�3�7���f�i�I��ޞL�J{���m�� /�'�F�p䌆5!&���#���Yz?��쫍�S�t=�ܡ$u�Ǳc"�Ӻ�LK�{zz�t
�}�2�Ms,���[0�{��.#`9W	'��GR&܊G�֒ƽm7Ν�D �R5#kiG����ݍ�>���&��t�o��f°^�/CT���Y�����N(�Kr��C��4���5.��5�Aͼ�;����Ux�)��vZ,`�;���a�
K�`��^L^�u�}�z����
���3��dv��I�|-:/�����Ʌر�Em��8~C�*ӽ�21t%��_=����m�<����AS��S&�D�z����#��������X������e���k��������a��Y���8�eBHU���/��.c�Eb�ά��yu(�vKY��b�=:��m��t�]�p-*�\e���ۛqS��q)����?�2��h���9�v�4˖sz���1��9Q�0���V�9Q�氻{.��ѝ�I��?����E�ž���5d<�c:.�fOGH�ő���1�B/�<���a&� �q��y�y"��ǎ9��H�����;w����߇ϭY���a�"M"q�O^�1� �?|��v=��F�D���k�nFo�	��]��o,T��J�������;�nJ�MQ�'�A��f�:�U���K�cS�v�"� �����
���Z�r�&̝�a;�>ч��}�!Rh2䅢C��p��i��ކ��Ă����]�x|�cH�E3,Ӕptv������S�a�9B���ET�'�z��6"��FFb������o��%K�:H�2�����??���~�m�ώ�#Kԗ�������X��J��C�r�]8����݈!u��|h;��`Ų�D��Tk����ѮAq�c=g��C�ad�f"	�û�A#gpx�I<�ګ\ue}�eN�&���F�oż��J����ȯ�qޣ4��M,�
����OQUbC��u�;KSj����u����u<`���C�4K���F�<�	c�C��`�Ҧ5����E�4=�@�=�������!�?���[0��N�;?D�1O�b%�Kz��uf��x�o����Ž0+*Ѧ尔�>��֍���P��D(3�[b:���������xB"�C�̬��9�䈿֬�Z)W$��b�^;E�vrw: ��EaD���P �0{ Y�u9ޅ�ǻ�:�]�7�M:�m�>�L�8a\�Ov�W��d��[�1�<�X����W�%��68:	� �6'�+৏=cۓ���SǛb���.<����"�B)dJ��6&p��G�x�|?�<����س�"��i�I��=�{��B����mc��D3��,�)�j�Z�s�p;���T��q�4U]��RZ��]��Ta�5� �U�?�}�v���r�Z444�y�D�N78�
�����S�Ei(���K9Wp�@Jszz'�o��Xև��)e�I����H�ۺ���Ooe05����TӲ�p;��Omá�U�i�Z�l�Fc�������{,�-�O�7��]G	y�r(Һ��şF�t�;1`�Q3xQ$�N�����"&*��c���-3B"�_Ne��G4�2J�x�x�y��:�>𵂨�$����,�ۡ���
(��t��I�Ǧ$�Lf�)C�	L�A.��mT2�U�!;��%�\G\7Q�+�]��-M�2�8>VDHq�'=o����)��N��1F�/(�R~��]�#rJ?� [8��)Њ�Q׵��*'�F�F"mZ�����cq�z�g��E�������4g��g\4�'?���+q�%�q��3g$<!���Y����⥽#8x|��'u�bf�{�0.�A�l��:v�ލH8@&k+�+��d<sv�Gy�\�"4�N�3y��!~�l�v��V��p�\��Ѝ�C�߮Ť����%�O�Q�p�%CL�'��)3��eYS���<� Vsv��K�251_npd��5�d�dD<͒b�<s!\!GdgRe g\�\��.9f����?�LV�(���:��Z�b�|�hK���cY���r�m��4�qO�_�yPZp��'�[S�l񞼈���!$17�+�6a�Ta���x�b�(73��"�434��w�s���MC����o�	��O��E�sTmS�}D8�TJ�o�T�iI�('Ԃ���sSiv|���]4���	���WCg/�Qid.9jH�F���|k�Dnxfe�
E�-Y���;U&����äet����`�z��-��2�����ƆS݈M���O��8�%������@��xxK�K"K��,I�nN��_��Uk��4{�;�s�a�Fp�s�d�j�Q�����Q[-;�}޹��Yt{�Ug����,��!�jy����^���uqi�9�ت����ew�mJe��
:�~��-��<B�dPɒZ�ӱA�k�]�Dh�9�sy����_�8�2ɂ�J%�����s���_%�j��}QB6]x��U���p�ʹq�m�P��#��r�/g |g͟L���>j��x�a��P>@�5#�D$�eo$R�d6�M-���|W<Ɏ5�kt��iL�b��1�vI�#�r���j�[	MyN&�t�rf*�o�������6����{�{b��)��5��3K\1�y�ۅ��I����˜�nwSv]UgW� H�c�G�U�,�g5��m�0�MJX�����w��^e��+����zu�JhV�c����z������j\��e� Rf:�M�2H��mx7�Y�Ͻ�:�����S������ƽ� |��T�g��r�,�q��.�x,Ϸ�=/Ӳ��'�=aƪY�$0~�J��1h8ؚY��7;fG)��؇���]C��<[����h�S�H����b;c��V�S�i����-���(� �e��\z���,�L���
��$:�M�wɮS�7��	,[�Z�u��t.�/V�\�CwabbN�=����VH0v�o�fF�g2���[����4�ca|�O����a���U��+6�ض<2������t_q���������$���X's�����Y��h��3�LE���jw.j_1��"L���݀$�Ͳ1R%tq�u�ӟܮ��)��j[�2q��wvO�V��VE�m��XL��c&C�a��۲��VV���_*�:���N��i ����KT�Y��1UL�1iܜ�y{�6�|8��e��0F�b��f�I'�*,��,!��s���bs��k2�~O��1,}�����}��<}��^�v���baY��/:��P_Ǡ�%���nC�w�Y"��D"1|���0���Q���I�M�����xϩ���D�V�s�Й.��μ�8r�4��`�<⬪�x�Dm�`y&��T��E6hǆ�먭��e�,g i�h��~'������sU�a͊e�d`D���.�%����,Ś�K1��/��a�=�v�<��i�=�^���)�yy �p�o=�x]�)����[_nÜ��M^�7���S7�S��
�UEz]0.݆�lJ�/Gml2�۷"<��J6�a��lF�U�Át��������z��H�8h���gA���(��E��p*N6������5�I��_�����n�a>qc�.܇FG�8d15��T��0%���{NکJ��񪚅B�f"Yo)�>��rC�iciQ�*��y��sk�1�d�,3n�R�4�2&ig|z���P1=�N�d�E��'�@"!�8Q�3��d�ir�T&�q�*�@����M�6�޸�bF�E�f�)Ĵ����@ ����2�`8謠Hp�%�NU��.�� nI�Js1�C±=	L0{�4�)�m��z��9΍Νqi���%8�y$OY��ǧ��9�9���J4+NcB�)SԆ���9�#E���>-�Ffۑ�s^@�xΰ�JH'����w���
���y���!{Ƭ8��1�R,e��Q�Bn;�r�PB?�}��/]��Q�]:y��r��w�o9^��\�L۔��&	��F�Sd�� �&�0�X�E�R�����j,�P��QJ\�L�I�J�´윋!;-�]��3|'��T��O�AM��n��Da�x:O��`L��B�	GN��c<��W��3���*?�$�� ��4��:QrP������9p���K�aR�<���4E�'kS�$��ٗ-�n��)KHXQA]#�l�9�F�t�w�0'1�Y���~b��X����U��1�NK^�����UTI��`c�Z��Cho�@"�w�j"g��i8�yZ�3/7eTb*����Z;�r[Qmd)���r=)�S'�`�����Ҏ�,�~)�'n�a��T�%��΂������*��.��6g�_#�ɸz��F��%� ���3RF�?ē�����Tt	��R��ڿdBY����P:�f�3�&���Q��۰�ၫ�i�[f�=��� {�XY�S�Ƴ������FH]����G��S���Pb�;��T��W��B+u�{������3nx�W�e9g>�����&{�@��%PA��AB����L�V^�&W��+��av�v��mYT�GP�pV,[ų�ullj���_���A����I���/���~�-kļy�W�2�S����Á���{�2�<�rڝظ�s�.G0R��LM��;�<�4L��t�z�~|��FlZ�s��XDZ&�N�������S�%�m�K�k��A6�۹����0Қ�aN�^����*i�:���[�e�k�ð�����b*���d2)����ڰƽ�qY1�����}��f��ה�#�:p��K���p�a�1���7P7�{�����ʸȰ��?}aZ�ȅ��-a撈1��x{�����a:�������k8/�*R*M#��=��E��}�G���dy>Wf��j�/��������K�TD�6Ƥ���&F���[�aw�e��w��&�M6���	���q�q[��n.KaN��[ؽ�m�R��X�ML��|�؈���_�Ү}cؽ�c%񐖔(��6�?�$z�^����mh��g��܋������v�3�'�}]ݫ�|�n4642s��� �{Hy =O�6���Hp�L����L�]���)��Α��lEpW%�Kc�8�8|t1;�,��UaJ�n�G2��κ�������Pf��@�����_C^��Û�D�l'�:��ƦR��3Y(�!��D�
��������ᶶ����;'!�F-�d�S	u���='E�3B���#��y�}O�IHN}4	�7\�y�Ar�0Bu�H���A���%�ԺfG>L�qV�IJ�y����������JB8w��З��9�D��e>����8~��]��q�J�عʒ�0��	��~���_�r��ף�����]�{i^}�fP��rDU�xKvG�F��H[^�Ջض}���M}eR��PJB��׶mŎ�w�оԶE�Ȭ9Ȱ��i��p��1$���#/��ـm���~5U&1�/ ��M�6�ߟ�Cvt�t�v*jr�"]���HLUL0�V��D�2�ʛ;��	q�(�<*�:Q�=��aMNN���!3=~#��'�d�2���,_��e��d��l�d�\�\Z��wN���r�H��/��Rz1��,����'�
uSI)}]�U�����~j��s�)�i,A�>};�\�Bm��JK_=����e���s?�7�ڍӧO)��<���fZ�p*CF���ŰH�:�Z�[�l�-/#8=�*N��~h�|u�J|��5��c�9��;O�S\��Fl}cY���|������h8L�ePׇ�:�2�2ŉڄh�T�nC!�;H%)��#�NriP���Cx|�\�2�I�,��ѿ��y��û|l�:4���2���~�*,2��#=j31��I�>�Q��պ�@U�C*x�<]o�)<ݝsq�G�����SX+x�$ӧ������P��С,+�ҥ+
���u��x�2���p�y���a(�,/L�t��G��u>��P�԰׳x����A��I�f0�ׯ|�Fܺ��'m�Hi����>|}5p����w����]�a�m�P��D��N"����k��� �ّ�%��W��7~�J�_�F$����/o�p���\}�G��,����C�3�~h��<baLi�b@$�H=�*n����ַ<G%$�9@E�&i��;���C�$�rR�Q���-�a�vR{sε�R�κM���/g�c�������w���@?��O�t=enG���E��0I؏·q�b�H;��h�Gx4 [$�IA�� �F8L���3<�l3�b�4jK�zڸd}~��%M������s�"��L�a��n^�P�9�����iF����j6T�B +|K�$F�Ɇ�}�!�R2� ���V:�R_`��������#���*��r=���9����*"�����qsf⫾��y蓝ŧ��J�]�J�Q�"��v�I@<D�����V�t�mNrؓ�)z.��G�t��O1��R����2�/#ұ�"r>�+�R�I���ҡq��e?�{o�(��\�B�#�F7m����9���K
�]��⻡��b4��1�Vf�I������w݊����fYЀ�G%HZ�q��m��O�#�}&��+�,��]a��a��[�����ظq#�l�Ǹ-�L���*%#�����&����=�u���=��`�!J���6ݑ���2?�Ť�p���D�Jg�o���k���MqN��=A���_8:}�kVK����&��i�m����)���;���IV��-�uw���=�oWME�͚��p�b���£#z�"���K)_Ȟy��� ���ܸ`]q	~��d�O%3-��!������%�aI�,�stL��R�̞Ģ��0r�a�����I�C; ���nx�N���	��D�������t�	�u�26'$�9 ��df!0���qIU3�s:���*U���2G���,�8��I��g�Ζ(J/΅(����`�1�s��t��f��x�a��>�ʊ
p�k���N��{��5�!.]6eD3,7z�LKSI��*���ܳh����ʹg�
���J\���mW#D�/?
�nd�,}���w4~��|gZ�X�J��X�Q�Hx�~�ȥ�Y���M,�<�&���,���16:���#����(��teI��%�O��f��P��<tr�ip�E.m�c�6�)������%��d00cX���o��%LQ�q�U��C'uԅ"*-��0k�t.��/3���dҀ߾{�h�GUM�s�H��H�	���/Y�kTR��:<<�d|_����Tju0��^��!h��wl>���Ø���+�?��9i��cH��jn�d�b�<E�H��0���#��/��ʹh�K�9��KfZ��(�����^���9����m�
߮X��%�af\t����aɉ�!�'�Ɖs}>K�v$Q,�$ΙZ7sy�Dh{�]-V6�a���Y�34�tC�p� M��!��Q|؈��XօC��J���sp��!Ĳ��L�a��6��H����CXZ�@Φ�l^}UV��]{:�t�=�o_�\f
��cX;�e�p�j���L�'옚w�R��L�O��m�V�!�WUE��ah�F#=Z�j�����͖JfZ4��ؿ-#��ȍ�^�y�1t3ah,�af\���&��C�Q8ή����"�L8Ȣ���K�^����l�O�5�����@�p�Π�Bգe�m���b�L9�U-q%&50����a�F�ep��=��W�~�+GI$ߛ�^��4�j2�L� Q�J�^�3�ꀕ?��AQu&�j�*��mԧ~�ᰈC�G�_X�zN���-m\޲��E�ǶnZa���+��P�Lk:e2�~�z��� ظ�����0�Dj1�L��� �p3.���`�"|�+��4��?���k��I���?�V�|�*����E��j��0�Ԍ3L�c�A�F�)	��*J���ڒ�iK�j��J&j����d!uэ��BD��&΅ ����׃s� ��{`O�0�x��h�_U�� ̆���i\*W#
���x�4GU�5�K;�*y�6,��y�g�Lc=gF`��"~���8��C6]^е'{f���ɞ�S~T2��u�8�WנI������u9B�F�l����_g�K:x:����~�Gr��x�u�o����;����D6,�b���Λ�Ѹ����DԴ�cLT�Pf�2���Pf�s
R��t�eB�!��m��i�p3p��V)�Ũ���=aZ��-���d@(�M�eǐc�b�qa�W�	Ӄ��'��~�Aک,�F�������;��d�/�!۷ṷ@�h˻67�.�G~b�N�����R{��~Z��ر�x������[� �䮿&�B�:�D��n�|ư�%y��Zt���{K.�e� Q�Nn
5�O�,{j�?�Oy��)H�Đ��y�SS�grly�T"��d�r�$�9@��n��ͳS�<��V����a�����:`
g��g7�:�R�>�3�\h�L�T�<߁��%�"����5�	9��m�\I�UN*�mޜ+4����E���`OWnY�]ỉH���k��`�*�j�h]ɽ߄9�,\Mwa�3_�]@��7���S���+�1�Q�P��Ɵ C$.���,�q�s�:8��p�Ǿ}{ye~X����b\�T[�\sy��O�i��J�(ה2��򜃷�2�E!�o1C���$�G���؉+x؎���9]�c6�,L�`*����F}	���%�-8r6D�q���8t� �M����1#�l%���[ܞ$�PS���p+�@�C���4�	i�T���
4@������@A#��^�?����4MA�1��y�x4�+��'�gH��Q�_�*�	_h�1~�03g1���``%~�ӧ��e*�P�L}}���cu���.Œ�{6����)]��;���G.*���w�ẏ�qY�^`�j���!#���ZzbV=U�|h�I���sdS3m3,/浱p�Ҷa1�]��.
l��k��%])�6Z)�����zeB�LTҚ7o>�pw���_��.+�{C~ñ���ҟ)�� p3,�l᣶�@���R�.�����*R��A�P�/�����޽{�P�G𛛪Q6�K�2��_
�ď_�a��N��mũh�C��W����=��_���ވy�K��V���'_�*�MOu^�-��q������*_��>��g�2uPOk7�lXy��Cs�HM�C���)�qy�Ġi4OY67���h���~�����S$���2,j_|��B�4G��IK$uu�&�h $�����dP�SY��0��,���\�m�,���d�B����M#M9a��B���=�<��oǗ>�	���c/�����(~��	<��V��YKY��g��cp%�25ż�c��w�=�{s�҇��T\�����I���o���Q�P�
�KC*�ē��	.}��K2-Mx�<z
S7�Fmp�P	6�{��B�gvy�~x�v?�Dؔ�@�8�'��cR4R�V���@�!X�5�D�(������8���f�� �JM�c�~x�MF��>��?��gzzʆ��X(Z{{��|�����Eğ�F
��{���^���.rl��Ύ�ii��9���&0�r?-Za������~�q=9�|��_�g,M"c0�� �2yD�b��
s�[��<r^.�&��L:��;�\��r��;���D�a���P��V���دԥޣ�P�����L�Iw�8h��_<�(��R�ŋ�l9�d��-8s��4����M쓝'���5� �K�	�N;��}��W,B4�lV/�t��O��]*�c�*ԃ�������@���ƕ�L:*�>�\$������p�;g0Ow�D��YH���KA2%��i�x[rDm�s|׷�3Ĉ��::�����^�EA �[�S.Ԃ�8u���
�ŉ�n����PU3-5��P��j���ރ���Ǯ����
���+QWӈ���>�E$���;O�oDbl\�sɵ�9����9m&f��R�<��6Y �@!��z��J��ȓ�=,�����Y��eN���S��}��L$��b_"�4{)~=�ke�K��Es&����&^��kDB�q1-�:�QN�زY/�T1�e[8\r,g!9B����2%&�{�"՗��	8H��S�״��e�E�FQS�F�0��{�W-��6�A�*�e5<�"5��M�A��x�/�Bk·��E1��罠9�h���'s��N��m�ɉ��֋-o���s-@t�ڵ9���5u�"����.H#(
}';ߖ6#��bQ�3�@���앒q)6.˹�C�< ��������=��������S�7�JZ�U��e˒m�d�ml06�&�!��	/�	i�H%�@�1�t0.���ؒջVҪ�vW��Sg�綹3O�]a�{�[�>���6��{ι��ϸ��UE=�a�9R�b��ɭ�I1-���<v#��:veL���!Wj��O�;~��ׇ~}����+e�� WZ��K��}ʹ\,�@��(N�tH���p4M���9>0�(7o��"��ޓ�.I[���P"��q�p?���8.�8���#�A��\�xEcZ���t:�O�k��my���7�
�;b��?+�.HƉ��s77R�*�?�Mp�^E5�w��6��%2ܮ�]����oy�]�~6	#�t���	��w��_'��u۷̖x��Y+]�g��9v�py'��dF:��234�7�L=\�t�ߐH��*�}�d9���27�%m������$lS'	e��s{g�gC�
H"˘�6ەɐ<���D�<<:�����U�3?!w�/xg��|�����%������Z���S|>��&)GdY��(�tqz�Qd�6MS��xA��֗zv"�n<�m�ʟ� Aʸ+2��dܚ�,�V�S:�wqݭ�~��U0�_=�"��$�TQyB�Ӧ��(��'�`�i�B���T�4��Ғ��D��g`ذ"���2J��f2V�#�j5��iAg�Q�|�ɢ%���ł���=��OP�����lA,�'!�|��x�D�%�=����k�'�	%|)8����	�Ae5�m�p3Ay�W�\�G���p Un���2uN�q�����O�ǭY���-a4FZ��#���7j�y�8��C������e:�����N���Bб�y_�}�#�c(/��1�ٖ�4)��t<�Bs����-&���	U� y=
�FKuʇKnn������xb�� ��F�XpBR
��)"}�m7��˦#��9#��8���}�'b�Iv�*.j�M`qk�]߂)���Dk����o�Ɩ�_�m�"|�M�i[�T1̘��׋]�s�p�q�J15��)O�d�rX��D�1}�mND�."�xPK����J.A
���?�ӧ��ү�q���F����&�{�}+�\S/�2fO �����o�ǖ��''/�*��2:�G�3.��@G�3�>;kK�ZR����T":T��@IU�����:(l&\K�����	��	�k�e�a��7�<�p�6rč���J^bɢ6���<�&�Co���V!gW#�cf�8~�ޛa���c�:��At��`8�Dˌ|�\�؍�}Xrw>�Z���4vb�E𺒸��Xa0�bk�\�O����0�R��u�O��iuY�Q�	���u�iT�41p!��i��+�_���1~�/���F兗������~� �{b��N&4�������m�O���cl4�N%�e�<����39u��qE���h�,yc�Q����u���%�2�@��5���k#�^pN�9��7�}J��	�tN-fT9��kA��7�b��It�����Q��4LŨS�Y��F���ȥ��?ɮ������������W2�T�q�SE��'���4�O�r�Cر�8���l0��\%R�n�!O���Hgڻ~���_��$1����1�R��
�;�I��9�Q)����<��V�NEN�����H�Z�q�;O����J_+n�����I����R�2�
�0��:�v5�>��T��2<f�hÆ��j�5�&��gˬA�מq�I��ZM�h�?.^��v�@2Ԣ�����G9�h�~�-|;�l�BEsK�F$_����l��͊p̸C�Y�$����	2a��)��3�WQ��Im$��YЁRqr4��>R��򰐌��26G���o��e_�U0.��rdS/�ɖöD�X(�����X�i�E�z�b��q���hx� ~2�W�I%�ӽ<�k$a) ZO�LMh	���Rv�5�%��zϞ�8xD�
c����>F�"��w�$o�D��}���Y��@+9�S�;ú�0�q�俄�Qn�c;g�1꘾Om5~�W����5O�7�w��F�y�x��
��TB���.�Y�Jڣ&2Ne���EIkeT�	и��ϔ�S��WTT`��b�F\;�$.k�B_��-ƶ�غ� �-)�]���7�^{�ezb�>s�&�D*�k��`����a�������$�"�o�Rm~��9
�U�_�cpx�+��a��Ո9�XD�ʕv��*de#�ά>mVהs%�}�rE�si������c��W$�h�Z&�����fI��I�~G&��8�*ӈ��0���%� j� W�h��һ��ʣ�v�X,r��Pr{���x��{��}��$(�݇�&w�*��GC��
e�*f�O2�u?*+��l�L��������S����{�8س�����t�Ȕs�HZR[�'��$��m�t���ܨ\9�]G6F�p��͸s�R���Jl=�Ó^F6�Q�/���ۉ7<�����DRg�������D0r�'�t�d�ivĒ6KC�b/�"�|w�R�R��E􁆉�I*�z!�ぷ�T��Q\12�(����e$~�h���'�>�DTf��`��%�%��άd�*�paFLi���wߏʤ�*�S����f���=�Sg�;��6��39t�֭��jw��S����-��N�8����1~U�����? � �Z��l,�h=�(TWq��6'�&�Jm�R����@E���0�r�b�m�<\3����. �41mx��d/���gW���u�!��Te'�U���@v�C6?+���K�Go����H�_�;��gİl�
6l��gOm�����Hb#h�)R�$=�C���׆^'�e��wl�)Ƽ���5�jE�T�-��yj�0\���W�Mšib�&dXR�Wj��q���J@�4��wl�c)����?%�4��Ň���4��c���6�p8t���k�O3��WSS�[n�':s�I�[�v?v�x_��g8ék���}ࣘ?1����{|����W_�O}�㨭�G=�Gѵ�ބcG���(s���n
��i
f��)!����pk�J�'��G��i�4�T�3.S-��������ƴG��q�+�3.nH��\�q��}ɧ
O�p���b��5���ڰ ��|a(	6�{���<.�t|��Z<���e��<quqIK5����GnEK�����D;y��|�l�n�SO=��d���`?z{���:��u\�@SS~��D��/��u����s�m�?�LjD2*�aq�˞��y)�u�
��!6r�CӈF��A8l'�m���FtX\��P!yݳ
�+`�|PCH���o|��q�l�������_���xõ����c�7�7�t;~������3�0u������!\��x��s��[1&��W\q�|�������{@T�.a�e���B2�b�>Q�bQ�b.�S��]���� !���#K����|��j�J����^"���(F��ȉ�`\(��>��Y��R|��e��~�mx��w,׃F���a�+U8ߓ�^���.̝��o��-hxZo���q=b�oA�yܱ.�w {��p�O��ꇞ��n�G�e?�m�T�55ՌaU�����]P�1E�l�kC����H�=yWͥIQ<(��@�x�='| ����S��*�4�q��'I�u(h�1/ȝC!$���p�^CӨE&mX�ߜ�)�	�qv�@�p�:�3r�k�x/�I���Η�4&B�k;�����oۈde-��=;0<�φ~�{�<�O?�cT&�t'�2e��j�Lq���ņd�_ҟ,d����$Ҳ��5qPp�s=�5����� �;ˤ�
4D:�|V�;�H�]_�̌bV���1%чX�$���.��G�:�<u60+�	pN2&Σm\.�(-�`J\�p�-�+��b1ܺ2�ٙg}��lD|Λ��ʩ����o!w�I�������.���>�?�����0�h�==;�ͱ�޼"��K_K^����\�?S�so�]3�]���/��Z3��z�"δ�p�'��r$��u	<?G~bZ��cZ�A���]c�:�]k����Z�ޖ�i��#\=�wPUJ�A�'�ϼ|h�b��~9M#�3�&��B�qG@�(c;�ӰR�<m��I�׸����͂�j�Te��<����e�Ӯ&UPb�\�wE����e:ڏ�ϧ��1m�t�^�
�]gp��~.�|鋟Au%SQ	��c{Y�r���W`��|0(�ȵb�I{�h���:r���9Xw�r����=�Iahd��p��6-/38Џڪ8����$��|L�P�m�НmӇŘH�Вc���۸�<OGw(�Ked2 ��<�q֌i�jQR��P����">�����%�C�eF7�)��(�J���(V��[�l6���i�.˗/G�{���� �
ڴ�F�O�1�C2w����N]\���J���`hh��:�T��L?�|^{z������k׃*��@��T�pW����1� �	HiG��Ƚ�8�ruܩ��q͇���%lU�T'���p@5">f��9~؏���]��]<�x�*Li���|�ۼ_g;�q��	|�>�l6���_��#�����`pdL�T(�*��������r�8�Sc���Ԏ��BH�w:q�0ƕI�C�v�[�u����.&�ą��7'�x�H�S3��)�Ù��*J�.B֍�C�q��T���0]�6-��Ip��^S2CW�i)*V}�m�?W���K�2����rƻAt����*"i�D�X����%�D���TX#��ő�..��������MFbZs�.@<�zA�\<�6��K�����ț�uu����1@�W�<\3lGfԑ~Q�atןՉ����(�y���i�$T���%UR��Ǎ��h�2�	�W1o��=ܞ�Dyr�ёa����G�����g�ɏ ���.����1֭���魸��k�O�)r�\�E�I@J�6ǐ�S\��Y���9����Uׄdh��&!q��!���>�{O!;�$"$�p�2#�H=&�#��*ӂ�Ss@%%)��o�BH�ȋ��	$��gڸ���e��%f ���z&�\[2�!Q|�m�i��r�%�,MX���d�,�vE3�1�׬���IK�8�$rq����^�X��k_G��赑��M�����b�ʻ<���䤤D#mF���b��z\���oO��<�����ђ��Hɀv��#4aږ����2r!ۺ�\��u����	�Uu�ɯ\0X]�����BO7�͜����^t�?��{���mn�ܟ��<�.�d�_w;���6��>�o?�d���~� ����3s��P�Ƶ����#�w���*��nBJ��m�c�6b�S�Qɸ<i�r5�CP:
�|�Chzf#�cm+{�
��+�K\�ƕ�G�d\�����|�iBL�k��6>�9�"�K0Q�,�	�Hᓐ@~է���ғ������_թ��ua����O�B%�mX�^��G�!|�Z����-qU�Z�l7� jBd��}�4󤿑�ש�XH=�f\�NGՙ�
5!7��x0��u�;�Sg���ɳ<C�����������������w���n�ع��/�}{wb���\���kP7e��{x �pb���K���i�T�m����H���@7�d���	U�K�yh?6��v<!�QBB%�Q_�R`�9���x�=J�k�#�a�6A��p�]ʘUb��'�r}��`Dc�ydֈ����a<a���aRl��7M��:sf0�v(�0�S�g'b�n*�����'�F���*�R�m��wG��c����49�e�ڈ�(�!)nm~u��\'bZ��1̈a3�ʜ�S`{��.[@�Ddm��c0��N��B{��R �����P�(,�o��q�]^a�G�5Oڿ|�#ې*
U��y�ho?�n�/o�Ξ9�J��}	���J�(�]�:yW]{3�1�y�l+�4�ʫ�;�?��1F	6�����M�Ie�/����#];�B?kIFfy��ٚ�
~���������.��s���:8d����
�S2.�@ظ�d�B����nq{�`&�lr�#�Y�G�?��io�+�ǟ9\��_<���Ē�������U��9:w�QD��#F:l�*��;z������L�G��1��/B��ڷ����Il�<IDL���j\ږD�LJe������࣪���]�\�� �P22�P��(W_O�-(���w����i\/D
�D�!�S;�8U'?5%�_ʥ覵%lZLU�~�P�2F�"^�3
ސ$C�cJ6������S��˙EL���]��g~��~��Gg�N����F�ޱ���YYUHbt�]�3rƌ��h�}+by(�	�#OW��i�*�3���qcD������))��RUL
�Z#�*U����|&���N���;�
�Z���H���$���b��Q�>s��nݳo?�_ц6arC��8�m�,x������_���߀���o��i�{{/`k�L�ًx�4�:��s\�"�En^v�{�;���Rt2y^x�A���ѽO����d�I��t��-N��_�7�������*�x;{��mbL�\.��ɢ�UC�b`){�H-%�D�P�y�^�U�F�ueA��ZN �*n�ܞHs�G|�R۰d��H?�]���.����=?��v�0#�@l)9AB>��}h�+X������|���8~O���{߇p�嫹��gΜ���iW�t'[ر��&O��Q���3�R��%�:�����cYyG_��r���%/[!Lû�c��ˇ���y%����.!�,[����*�:[�E��qeB��	�UHbf��b��f-J f���}H��2�L�4.��y+�@��FdI���6E:�K/�(o"4AC�X~�x�,���XY��3�6��xy� j򌻏u���U_��~��V�hɖ��/�U����v�>}��!Ya�_/Q�mm-I�|����$����+�-O���g^.F���q=_���s{ux�]�܈cna�v
y���$���f��>!�mX�b�-C>D?b��ض�xr����XQiK�����Ee�ƥT,Þ��LuFq�������AQ6_|.�Ё��Cl۱Cc9�������
�0uq���3gϠ��=]g����Q<c���?8w�<Y3B������67q��Q�d��Nۛ́�$��%+K ��6�mʑ:�GD X�~n��Y�Z����C�gO�~�����$����C��w}!y\��I�o:�+/�mc����!�V�T�M�@b}>�{ջ�;0���m�(s{���^�Lںp����s}��x�VbP^������T�|gg36l�����#��ZbylRl!�jd3����]VJ"�%�I��]�@��sV�g<�%�Q�Cx��|���0St#YD�B����������(�FzPh���"z��+��F�N.u�=���ρ��ׂ6Hϒ~C\�@�����`6���Cd�:�곍t*��B�Ǥ�����*�mcxh �����{�r�!����*rM�����y]��j#}	{�P�T��"���^禭��'��F���\$,��
��8n�B�ehX �?[�g���͑�T���㒨���	<��9��;֡v���`
]�,��Vᡍ#8�~|��(*�T�1�O&�96qk��������"�0�!�f����|��Z������?1
t��U���Y�5���&�M����^�-}[38����6;q
z`Y���o�ښ��@�A<3�#�G�هv��Y�x����ˏ�a.��bzN�xfp'����~|��v���o\�Xq ъi��>�"��t���"���~l<4ʴ�4O%`2!�}S�;�ӂ��l�@*�F��,Z���_bG��D^�S�$Hh�f��I�8�U�!lK�k�BH阫���Vqr�J�ɖ;�H� ��rI�3�i"PP5�-�R�@�!?Y�W$lB~�ʵC�W��e�uR�:��	����0�h c��3'�(�=��0*Ǜ����X�ߠ�0<�h!�<�%C���)UQ�SC&H�6.�v���|�&���K��1c/�O�,#�� �p��H�Z>��z�=��{�X�p�#�Rj8Z��9�q��px�_�v��e2�*�a�Ґ·��rh����ӧ���o�a׬h�����~����7�PO���ř3��v�e�cY?-����[�����p�,�\ժ��H_/�'��KC/��u��WSw�Bδ����c���=gL1�ô6F������u��i������-U95)��M�X8=�HU�x&6E��������Ql9\�%$��;������q���J���@����Ȥb��!c�����=)�������i
�X��s�c�+�J�Y"��/H	=�Ւ���Z�p	�/W��ҼFў�X��
��cI{��[
*Ge�VP9)]�v���xZT��hU�mW�}�:�]͕��@�����L�V��d��Ү@xp��.ːx�
��hҖEX�yB���H���^���)s�R:��(j�(N&��'�={��ߝ=��+��Yә@ӊ��.0�|�k '��L�ߌ�����_��L��E"P��8<��gN��/���TEF��h�"�^�2!�wk�����j K�:��������A�~���R�8��Z�d�wH=<8/*T��ؘ�&m�г�3�pc1��XjIO�U�P
�d�-Lz&�
f�B�[��s�R`9��_�d����$�붚=,�H�$�m&|�Qa2jq	$KaOJ�q�>Q��)1���ȕ�>�	:\i�R��Uj�p�0�0���6#ǯS��٨u �P��5i�R��T����d�9
ǲ�-�Ӷ1���N1ڔ1��V�.�sԨ�B�~��GWO���9��	�Ir]�����@3=ΰT6�J	�L��w\l.X�ݘ3F��?K��>���X��VPmVg���T,n�~���x1���߱X��	S�3��Q����I�Ǥ��-˵H���c�a�����Y�ly����D�ԩ�H�E��͑�j��� D��p��Sw����8�g�z�J�d���:���Q�M{�.Y\�U�f������I9B�u�0M�;�$:�<�Յ���Hx��!�?�Y����mm÷���]kj�D�<���k�G�u^,y� o�Ld6.���h�w0��Pt*Ղ0,�`@�&�^�ӳz���:8P���P���?+��buFE�^^3I�,���O�!}M�E-�N��@� *��М�6X��V��f�p�{'w�{�	6,UI�J�*��ߺ2|I�/�S4��s�m�{��e�,��D]��J��4G�0[�X)tb}/��'��}�1�6�Cb&��ʖ�UV^����J��y��gX畸�f�b]l� �X���([1��r�3����Zr(�_�`��r��3^�a,;%9<2�=2P����垜/3���u�I\_{�/�E]e��w���3��1@���"C��B_a2"k���*�L/�R�)��.d�J(���&	�s|[�*��l!1+����t�W�t(�`6®6�w|?�YD��I��v���:!a��_ٰt�`eW�劓T��l;�5#�H�6�{��O�Q�3қ�1�r#�w=&}A��8{�q~�e,TC�	��ӾE�5���v����i�;��P$ʵu(���S�b �K��,��RV126���rϩb�t6�`�$cH e�-qO��0'̩K���HUU�ݐ^ԍ�X�TQ%, $S���%8NR�5<�a� �wĖ��+8�M���zΑ�0tXE'�N%�ԲHF�{��Ĥ��N9=�;��VB������?����'Hۚ���~كdJqQ��S�1r{R�*N�ĄCV"Ҩ��01>]\��H{�,����d{H2I�:���`d�VI�-��f�'�Vc����9�X�����f(�%�X�I߆7�G���R��Zs:]����w��{�c�R��s0|rj+TN�*��oLp�U���p�Ji�
n��ɼ��`�gƓ�T�����4)�P�2�%���PM�����1�6S�\�U1�)m!1ˍ�����]��}_1}�y��᭢<g:O㛯~�iQ�ҩ�x��w����������L�g5��=�&�V!�����뿆���<>r��[F*`M���;+����D�|��X�*|���U��X#dE��؞���	��7�WR�}雳-%	v~��#4�J�̅	�Nx�7ʷ��}Պ����'<3E˅��^3�n&p%���T{��&3��1Y�I��lK!o�x09�n �\d/Ĳ���eh��y|�0	WK����֐A2|I1D�Hц�ٍO�o֙��eT6�S�Iڴ\-��j�I�y�O�r��-X"����#ڨ���s���;�#3���	�uC��T\왼�}��ȿW����Ϩl2%��q�ܹ���4O}�8OjA|�VÂ�&xOP=��zQ*UVOF�����w�TN�6�|�kA�g�l�M%�"����3J�+����;�ȹ���g�p6�Ӕ]���0��Qȹ���(ل��P؝������qxtD{�43�87TR��\�6���	y�,j��M �|Βa=G�T��A�ɓs��P6E���5X�0���W�&����a�w�2`ՙrM��O���<�S+�s⎯�6%!IH)r\�g��l�F�����A��|�����qۍ
+�%���b�,־r�o��S�C�S&�S���3�7���Xw�(M�Y58]]�8��c�� hs7$�p����nV��$�F}�G9��$Im50��|8ךV���c�o�p��4���Ѐ�������%�|��(�VUi}�㩒�(<�[S���˓>���p��\)VK�l}A�"x�:7�D�
qi$w^�Q�EH�M�1qv�]�U��G�kE�6����1�\���<�*g˅��IB|+�&V��f{��s�~c�c^�}���<�&K$ݞ<�;������r�]�Cu�k��5�z�8�h_$�2�O5v�d�p�i�D5<\jQ'�f#UWNS�OKnR^hl=#,��6B�_��<�}<���i��"������=<��17;Tvi���%���Q4Q4ݑ�g����\�CLW�ōV�;l˯�ҝ*<}3O�"�����R��c[0��������
��=X��$h��Q�l�����xǃ��8
\�Ns�ω�5O<ł�PUI��+�9�2�4���0���ދJG�xCC�H0=|��<�����d!��FǙn�r�6�����n�E�i,*��%�Pz�y��
�"w)��E�;�gZC><dE���v�Z%<��+KH'c�K���&dP�ܢsO2v�#s��W
��ԳA���w���1-Jx���;?����U����
��	Q�7�I��8+��H��Բ��Yܹd@?^_�����a�1���h����K��IH������+̌5U�q{f4+��M8��j���gVj��'�u� F���W�g�9�1 /�����$�4�W��e��~�''`{��V�B�,Hd�Q>6.
m-f�A����j�b�|��6�~�\$�"Υ�]N9�m�� ����;��m�}�ZrP���SH��P���b���.�-�jD�d�g}��xT�݆G6�ſ�ln����i���٥����$a>SP��Y�)�3)%u�R�wQ��cQ��>dP�KX:R���uh&\�$�=���UUU��6c�L}upp�mL}�)\W���wy�G�R�Q��|	m�hnn�-W-�u�+0��M>���^�����ن�^�������u���}ȸ����
1t����Ո�}�'��|�p�=��?����]3��Xً����U���{}�[�t��\�z�M���]��]�`"���q�+�Qku���#���o� Z2�ӻ�NOL)�����}���M�`ĉ�5�"P;}Opq�l�a�T�/(���q�L��\����`M�]P{���H���M�38�qs��"�?
]D)֓�$gZ� 螮����Q���y	6���1W,_�!il�������{߼������W�X<3��Qx��v>�as��i���df�5��7ml?:��l�9����l#S��X��3�u_�������HK��!,��V�g��C��G�t�P(!�Е
�}J:��Fyv��^���~̟�l.���s6lه͛6�	1�_�i�vZ
cG��UW]�?zSf����+&*��8�U#�in6������1<��
�!"�R\���|Co�o��A��>.�e�8�^����+Z��v����s[� ��;�������KO=�ڠ�J}zf�nL�z+�}�ͨ��cs�f����{?܃!����)_��{������ǈ&3y��L6/1�yW=�U� �VWJ﯅�Y��B�>"#7�7�R5�YP�?������-a���n<�7��O'�͵�镍4a(���t�9i�Ig�_�T���TA٤.��>eJ3�(N����?j����9L��BKl:����w�˔�>~O.�W�.J��t����	J�ﻩﺶ��#��t�ś�����7,�dc<�K��<���2B%dZM�����v�*x[�V���π�LIBя+�4lM%����'n���w��^�{u�S��������X9���?l������k|�؁��%�b�%��ߚ��MB�1F�������O���;���?�,9��s�3K�_�Г���ب�/�|�A��e�ڳw�:�G�g�9�������cb�R.@�[�݄���l����~�o|בN��{6E���'2��d�������G��[?)���O!����6x�S��d9N�/�s;O��0ݸ��c�V�N������EIVj�.ƧxKR�1��ԡ�e*�;��S���K1v���U,��{���0)+���]���3X>G�դ�:e�:�췿�?��Ǟ��ޝ�k�T^�|S�"[�fQcZ�;T~�X;��]��ϒ4|�ݷ�W�jxC�;]D�Ly��r
Z���⃏ss���%:5o�<|�=ע��Q�[�l�k8�6!�za�J�������}3���'�.+� �>C��19p��#�C���`��CL��°�ݗ�d=��[��X�V� P:-��)
P~.���D�nuBL��s|
���T��ܥ��+�<,�BB4���O��V-�rJ�Bfq&�6��>:�������p�ҧP$a�-����g".������U&l�VW�/_G�5���o��?��P�y�Q�iGy��m��}��VD�䗵�0�M�|6F@�P�
ƈ
�i�D1�a;Id�R�A�r!�-G��ML|��ư��+v�t��EY����;,��(��g��敋�����g%h���h܇�����<�tt�*�7t�L(KO��gȝX�oI���mWL��;���w2puM����}%��'	R{�F��Rڷ��>H�+?���G-r?���Q�+� ��GA�W:�Z%���7k+�*��<�]���\M�Q��o+��q�rT���h�
d�
f�A�!��c��:C���ϑ:|a(�T/�U�"2�oŕV4v�)ہs�E)�zH���|
���s�|���"-�:;�`��b��<��j�\�ȟ�������q��mBrW}T���l����>K�tz*o�Pd���d�x��p�w��΢ϟ��g+I^���C<�L1A��kl�9�S˕�*P�^��
}Eؿ�	�����$�@��oX5u�W����+Q��waUM�e�9sz��P#��8���t���ٳg1,�	0-��.��r,i�A4��վ��»��<ô3�w��h`v'�Ν����	��B��P��Ua�aJFp�Z�%Oh}Caq�c���Gӎ%2��*��.��."�!*�k��^en����?+��7ʯc��g��f'iS�Yjj*��H�UzR�zE��k��z���K�(�rbt�˘�s����s<�==�8��~#�_7�qa�����7n%1g�|����9�Tf�DET~]]=Os/`N�ؾ�����x��T��nԧ3��3?��<��'&Ւ����KL�~
��D����	Ԏ3O�K%�]J���!���%>ꃓ�a,/����Zv�|��M@Ō��6�����)9�� ��������"c�(��;�}\@��P�H�$�4�55��	״���Ad�JT������x-۱f�b�_`����R��yx����&*mM8�d��VԺ�i`b����_�$�����/�D$��s�窪x��bΣ~�*"S�5�S�O�Ϧ���CI���)�)�B��	X��\�c_���Q<�Uu<�;'��/��X$�^��%��y�m;d�U�������Zxcg0��x��ᔃ��,2y��acH#5�#�	�Ch�Hj#uW�1|Q��d����?��M�<Ѯ`�9}�{dC�"���c���m#���G�O��H�r����o<��M�Ƥ�3Eǖ���|����%?B�u+f#;�+����.]
�-�4{����:dz����
�o�� ����X�	5���L��r����c�#��X�Ki~l��ㇶ��2��y }���L�%�{�&R<r`"~��Y�e%ԺInL�eP�f6+~����?��'���>��㍌KfZS+G�8Z2�N�����v�,����g�Qh�6l0&D�qG<�\R��ĩ���W'bep�����@b	��z���񖻰x�R��~d^޲�N�!-�d�R�����������}�ر}3���)T[��/[�u7ފں:~e�ٰ�iV�q�c��	�Q@���\Hx�d-Zg/���ڴ���.�Wo-�,�,�t;��g�%�C���N�
���M����J}f��^WρT�{���0�s�q�U[���3f����ʄOq�����3��X̠ý��d[|U�ڐv�ͣ}׏0&����"��H*�97��hZ0E��g��9�,��l�K>�KerXȞUӢT��}{S�?�Ǻ^�c��r�Z�f6�^��[����i �{�mV@%��3N������Kَ�Qe3���3IM$��bհ��Ŧ]�AfN���'̴Tf�	�;F}�:a��J�Dy��U9�3i��q���g\
���>ZV_�el%�5c��������lCε���u��-��o���p��a̞=�1���g�fL�7�VU��;ގ�1-�KW^����L�Į��8CZ������㓟�=Ƹ���`�#�mX��Dn	�4�V�؉�f�q�Y\��f�<*����:më�� ��1�!�����e+�")�I}@fD<���`���E�F'K�O�0-.��!���̈́�&]�x]�C��n!�߇�����B��ŋ�.��Ç2?�|�Ƀx�%��8��c�Ƌ���������f��hC&���==�nnC�gϨ�>Nس��`���J�<�$2�BpBIy���P��<D�-ZBm������X�̤˘0��S�>���}�4.)� �
����@�-z�$_0���fO��o�-��z���;[1��xt�9v��z܀芰vO,j�74b����p�8�L����ˏw ��@x�`:���7V]v>��?��'�_�t%>�O�=��C|�}|{�_e"Y��~�?�⋿����02,ܪ˯�'>�/�����������z�IûW~a*J&+x_�	��Ν;��ᡂ���z�uf0ը�;]��H� B������,�b���	��/#}>|����?��N��)����ş}��n�Q������s�'��Lb�"�xb�x�Ձ��IJ�9I�ܛ�q��9"�.��0�L'��c�e��~ �63��{���X==�rB��r�V��d���Ƃ��ˎ��c��א�yn�N\y)�Z.��κ��R�'MC!@V.M���K|1#&Ug�6����D�	`�lC>%R���.y���Zc���,M�i�;ڍ��h�Ţȟ}�Yo��b������2�pj �c����%�V]M5>|�26�7�ur8_�Ak6��C�1�e
���3-O������I۞������k܏�S�a�|��%o�W�����j*�qө��o�x\ f����]x���c^�|���֖��ﾏ/���l!��k�<��wQQ]!��pƂ=H;�ֳ�(�����0?�'�U�l4:�s��W�ļy�`͚k���½����E����p�b�z�1�"bNd,�p^�ޖ�UU���:���#����2�&��ٲ�����31�aϔ���˃�G�"u�Cn&�����XH▖$��TzØ=�����N���:'��|v޼E<7�[)Ƶ��[�DY��i�i�V�94��L֪�id��>;	-J���;8�T>���\�غ�_�.PE(E�x��H5�,�FR�&��D���ٍ��@CV�
΅=ܠ����
D��ٗ�9���[���}�8KT�'$;���ғI2��q#�����g��E�ݍYLU3�\�g2Z�֡n���s�o���!���%m� -�[�d%������N$!<hG�����]n�b���J���8���(�zD��k�=���:�t����B�P�y�Nvİ�w�.[Z�app��ʀ������&�H������B�q��vG`�Ƣ�1�X�w�1���ˡ2��(1����IتL`���q1I��<��w�	���?�	�N��g��W�
�i�$�"Lr;���{��=��XL}�L\E���@��AY��ս\�un���8���lgn�c#w�w>MW.����&~�5aI��~�����Hd��X�50��_#:�jD���߽�,k���so�/l|Yt�˔� v4�x���-K&6��g�$���oq�|�f�1	Mc�jUU��:ă�m�����Ȑ��"^<A?�C��D�w/����V�W]]��_�(��f4��h��RQq�ƿ4S�M���Q[[�$-==]e+m���
�G uy[�{a(QiR�d�~�����B�E9�
���$	�.	���8^�D^�1T�E�$q��>�]I�q�&4�r�HȖ��yO�������i~��#�����?adܑ�J��A����l<�Z�,�+t��ƫg�b��*D(�<��2���l��X�AD��czϗ���
�KW,�O������@y��IZr�=�أX��wp{�0"<�ȃӻ��#����='U:�}�_5O�DxM<s�#��Ρ���$(9ɭ���}��w�S�L:�Cbe�74!�Q�KN��Hҩd�&�둋&���W�31�'~�#���'��T�ɟ���â��z��ԥ0%څ�$��QQ!^�^D�p���H�$1~*��C0���O��+U�š�_b�Őx�v�g�!׊�`������a���<�3�&RZ��泓�B��Y}�
��mڗ� QZ�SK�e��R�(�G�7cٜ[��z�`\���3髟-ZrΪd��������m�G�����f�C?�9�;WㆶAԥ��|"���c�E��cǱ��W��22�$�N)-����e)#c�[�K��-É��i� �O��S�ʬ/DR�������>�ٿ��S��H~��3��6�<::����͝���`A�"�~J�T̚u^޼gϜ�J{ŝ�^Y�2����)\w}:���-��$��]8@� }B$vx��uح����XU\��չvXd�e�R�%�1���)g�d�d/�%�@�w|�Hy�Om������N��{� U��2�j���f��j�A��.%� 4��S�A���~�;���1�|@��.
���uU�F�F�����
\Q���锢|�����~�<Ϛ,�"���`\'N�?�=��݀w�����y��o��G1��Fl>��'�_��C���p�����L�	8RSLO�`F��h�C).7F����wv��2[faQ�&��D�^}n{������F�����	 Dc�������Xq�X��H_��?s�r�e����N��`XЎ���Ϛ��A1SZؤ��{�d)o��ؾ�Y�[�����(G����?#Ç$�0S/�S�����ok����6F��l�&+�P_7��9�9؎l�p�'߁��R��d����&�l�=���T�\��(�K	n{���T���C��ӥ�l ӧk�7F��G���K���=z����R�
M�"�xx��͈�@�m����`�F*���JT���p|5k��Pja��G��_��K[���߀�JUC��۲��8;V��8��v����nct^7�E$���������O`͚+�f�{x
.�;����q�:���K�*�G����d(R��*�5!ĝ2��ڻ�E����ȱ�����a����.�<mf̜��]F�*6-���x�׽k�˸~����[��K�����Ȟ��/<Ö�v�����T��&�Te����~�.�簾f��	ǹ���}���)x�k�f�T�#�(�;����C�������׬Y����ْ���)��rU���*�q]<�� ^�z~����t�%����=�I�jhh�pʂ97p߭�z(�1��"�U?	�榫�����h�]�6��75�Bo�|V��{����)����q}˵����<:B�~�̕��!1Rzc�F<�u�4�b��=�p�jPE����_4+���!�r�	.�r�8Ē�&�(�y��}����=��m����n�Ŵ�k۞۶m囐��aXD�+�?�`Η_��
���DB,��� Kۨ�2��Y��X�6�������q��9z��`��݊w��}��/|:t^���T�����c��w���3��]�>{�KtT~��7bp�OJ��Slj���vܲ8����l���Q�Ɵǋ.���)8����s��[\,?�5��~}�W�9�2�{P)����5�Z��w���2)"ߩ��v�1&T�``�$X�&7Ai~�1�9s�q�\j��z.J!H�'��x\"���S�p[�M"��uه�����b�f\��3{�ۯ���}��^��5˨L�܉Kf7K��l,��K]�U��+�V���hĊt�3�RcXnmQY��C�C�&N'�Z���ό��OJ��K0,��Lp%�XgB�E��*��EOŽ)�r;z�y�<�W��/͜��_�ԁ��,v��I>	���i
֭]���F�0nO�wfD�Jf�mع�O�-uv����kp�;����R�:u:^|�	lu�P[U�'�չɄ�D�_�����ş�����3�LH>TW����~gNu��#����J�y���M�-��]��U?_�uP�s���H1	e��j��t�@�9�f���X�+�0\y;�����`i�ۇ�c;x\��rE5U�X�v-���^ټ���)'��{�K��A�s��~��OoC��P��׬���.n�bze�>|�ͣA�����QMS��j�KSb,�����׈��S�QI��&4/��Ċ�g�7y����q�'7��x8�څ��Uş%	3ڷ8�	��ɧ 4��Pri�#��D\ٵL9Ӕ7���D�ă�ה-s�~Jk���6Ĵ��q���I?��$���3�ux�bhd?~�K�b�����t������=G����'.k���N�X���C�B-�6�O����������3��Y����a���q��+��e��-��ԉv�t�a��K�71��	�;{R�LlR(���������d���?�~��,��o�T�����Ӈ�� ë�����Jŗ"oW�k�M��H�
9��hLk>O'�	Ɣ�2���H�ٻb�x�I�����|�1�=�0˜�R�qm�Rn�j�XI���!���n��E�#{����#�gVU�g.����Y9��ښj��]��}��ȾN�Mx���o=߆(�XҲ�Cln��Ʀ)'p��FP=��nϒ����p�!<���5óG�i�~V<�3.z֒��,� C�n8�Pr)q�09�����"TΏwu%��� �o]�ǒ7BeX*h�]c
C�� ��Q����)�C�ф�0I�U�і_%�?/�������~P������'#����}����1e3�Q������~ܽ�v�n1�lB�Ĵ�g�	����q�غu3okT�T��`?v�،WY_DC�tɏ_������̜]��ʛ��
�����|�nm��t�ۀt "$OBA��=mZkY�<n�3��
ec��GoGll�cc��0��q���a�"���/+�Q\�:�+]Yobz+��}K1Fہ��`���kʑ]�c�ͥak.;Y�T�n\~�Ռ�5���ôԳ���m���l��/�^����p�$�I@�&x2���sԆ�	�O��7�n�/N�$!Ax��%�rNU�9Ectʨ��לØ\n ���ĺ�Qƨ*�&�)��A@$���h���R�-�ግ����p�Z����p}Z��C�s)*v��B�8�U�$�(Ҹ�w�Ǐ¹-H0F����)\o���}�|�3���׼"�z�����K�� Q}�Wr���4��h��eH�}gj'�J�q�G�l�$�tEn d�QP8��2T�PzwH �Ԫ�D���ayb#��_�,�B1�a��/A�>lJc-`���F�`4:�;���Yt��0��E�1��[�2�쾬�sLZos[��Y�>p_��iF;���g$=���Ke__W��V+���M;Wц���(GNs-� ���ȹD�&N���G`��~6W݌�Q�(��̘>o\=��H��Z�\�X �JZ{��E�i���d���>����Co߀Z���buU��E�Z��,e;�B�KS�d�*6�t�q���R�o��w+R����a�P�a���o|;�I�L��w�Q��עD(~�!po!ߒ���h��څ�l�^]��l�;1%{����������5Ԛ`UZ)�>�����*�ZTG$�
�{)O�Ip9�X�3"�����6�Ν��b1�����w�ZVl�
Ctp������`���R4[���.�uK��`j.���t�B6N'�&%�Kc(K�[�݂6��u[	M��݂K+w3��_b�V��A�2���V��9��?��߆��m*0��~<�R�gǩӠ�L�㪓쨥t\��ɨ��pD����)�5�֥�e<k� -���Mㆮz��扗�n��X��wP�+}T�p<��&��u�<���9Iu<��������q����n��"W��r�Tޑѐ^�<W_�zލ��ĩd��v�� Ϥ������8��w���AkYD���!�TlY%��:;E4�&T:-�d
�3�CҘXPED_�w�P��������/��4T�ܫ;1z�ϑlbR՗M�7��SǏ��f#A ������µ����|��NW�g��">��o��g^�ϒq<�?����~ģb��ҕ�#�!���W�����?d�L@����o��QD���#�c�Յۮ]�Ǟl��S�q�Q���k�_�J����O�.4 !Y���	h,x�8�	�J[1.u1G:���袪�m3���d�E�wg�)��d;�?��&�$���f��PQ!����7���ݼ��Qqw��s�Μ;q^���0�ʢ�������H���lvjc������^��G��f
���r"]�1�Y#�1�B�?ࢆ��}�܂�CFx�h[���"�q��|W��x��Ҫo.Yv�;����/�����Q�Έ�������\��9�]G��WG��Wͥ1�9�r���h�\�	��;�� ��-�vGL��Q���B-�bm�i�Ta����#�m�Q���H��{*�/:���Mk��C��c��T�<����<��5��}v�CصG����QYe���%l�g�k�?5*�9}Rʹ;��A6�婢��H��V�\nc6m�j����䗡�ޟ!Y��i���M���T�t���TR��Qi����P	���Ű,���	��Bg݅��.�I���5x��<е7?�����g:��]xi�Q�h/^ncC-{�
�ṃ����̬\?fT\��s9��Ks�i�V�����w���W�b��X��0S5"lrf/İeo��֓I�
�yJ#>xs-~�x-�cx���x!�Ww�G�X�-���g�c�k1/юx�x�R���ĥ:$�p��B�Ƚ{w
� ��Ҷ�q�^�zD��$z~�8�P��0Z)�� ������E�9��� �͑���]�1�&ȏ�ơ���Q�0��)���O9�~�:w7,nBks5�dcã��LesaWa{���F�����r�%`�c�(hj�\7�e�]�(j�. ��!R�)�nwN�}E��K��Qi氍�ɰ�!��0B�&���Q� ��pi�YF�]b����}��YQ��|�D�E\�Rv� �;�ӧ�b套���v�Ps���җ��9�eKi#����X5���/��)��I�Q�k�C�j5�$���1�s#X�h���?���'�q�r�c+���6��s�X�����(�WD�isޘ�ж6Fqs[7jR��Pn�)���a�_>���Nw�M	�)��!�V�!Oy��ݴ��i`h7.�ڃ��^��i	4U���F�H����_�=��Ar���A��X���!Z���%�e�����Sh�N�,\�r%w�'��B���wH�4"#��Taڹ���r�q�`�����q���_��g7%Y�*`�H�|��]6�����D'@���߄ǟ�Ʌ-��S�I�ɱ�B�g}�H�8%�g�����Z�x}^����3HA?gɄ�o�@A#���O6Bs~r�0���l��uy�7��2B�R�P��g����,�H��r�4A�0E�d�]��ym�sOw���(��]��C������Y�x~�]�`��H�@2�=83*�����܂��d'�}�E3�9���+P��@��S��m��X�d��Y� �E�yi�f��π^�P�h�Tb���
� ����P��IE����m&PQ�\��gm�KƴL���v�⥜<�c���v�ƴ�U�H�J��`�\Mv�ή|��O��gM	�����i��)l9^I�%��śF9��P��b"�"��_}j*�����/<�pưTx�Y`�e$�ri�	Զ$�c|�.�f�<�djs
Z?|�#E�8Y�I'��;}�8���!�����p�T��@x�7����^R磁��K��6j����$c�!�LF{�
WES���JX<�qC3� k���@ ���5Jx34!�o{�Q���L;v`PT�	KJ��zr��%��o݂����8�c�&9���x��<�wG���TY�ȋ��B*m���T���2����зܲ\Ǵ�� #r��Vm�?r�j\��f<���;xğC\U4�ߐ"7��l�F�LR��� o� �O��}%�i������;��X�Ԟ,]�2��J�b�"����ʫ3�L>��n�k���6>�G<�R|10�L��a"&/a�H�;�;���/dϰ�P�$�bA(��Qf��ckj,#`�E������5URc�sY��x���v�,K�<@�͋�Q��`����M|���IU�[�882Om?E}o�R���$�v�~V"��(W�c�`^T�;�]��a�eb�Qd�&�Lk6Ĝ�ߒ!�-�d�lM%��q�!M3g���o^��\���n�vKI���F��Y�PY�<��ϟ���*G%���&N4Ԅ��5x�5y���Q�5Sj������4$(g��ɒ0l��f{�;��vXR��3+�~�D<������31��>xUBr(�!AYAW�~ٙ1Dm�5���^i7�j@;�.ʲB*J��]]�F�z��!��T�-�����4�-�a�I�Csz#*�a������[���e.�A^�5p�a����Ln��N���-�>��yv=�DL(|`���Q%9�2��O�.([x��S����+�Y�'���X��Y;�0t�I>bCV���94M��(�rk� *�v>6G[27��H|2qF%�Z��:������y�D����E�u��\l��2�w]��[�#6�Sv�+F��m����z|���188�.0��2�/�)W�[n��{5�G^����h@��`W����ǑK�!JaK#��;V���\/GR6̄��'C�g!��dR��-K�c]���l�1�K3@�@���RR*��
JY���g���D�#
���������x�!�#��"��LC�s^82��W̺Fc��"���Bp��Ψ�8o�B��/�I���͐��{�%i�,�x����_B��&��(5��ɳ%��0��.�3KHx"ߎ�7k���E 7���*K����(��rr~�dg��k�=�丮3ѿ����r$@�  �(�$J�H*[�Z�l9�~��}o�����޳�g뭽kK�,K�h[�DR)1� �L$9�`��3�^�s�u��@���!������n�:����?�g���9���Ȟhcr���(�_���~JF�0rr�#��z�������<8��G;�������Ms�Q*�Bt�]$5(Dp�Ƿ�9L�⹓�uQ���>|�?�����0�ִ�fr����olE��OTb�]�����寅P#.���ɭ_#�U1޷��_�/��z�O���\h�p=2�nrN˒<ߥW�3���67En�:�s�P���Ђ��y�)�BzgW\��!؃��Ơ�-�����[܄�ٺ�j��8ߔwy�B(@ۡ��Hi�y�z����TQ�Abaf���Y����+�ؗ����A�s@'�i�xWmW����� �I�kǠY#��r�s�;��
3oW)v�����C�Pp֒]�x�ԝ����痘I�CE�dFX#%d�eK�c�̙�8r8��m�?���A[|9?��Tzx�u���y�y��HNR΄�̽���2��e�ě��qD�\?��p�*|���4�Uk��*�<�v�K.Y�f�S�B�����9����D�پ��~��7��-���%���OQ1���	��,��U�m��0	`��S�\�w����p��<�u�G��y�����;����L�&s��L��
g���c��<0P0d1F�sO\�m+ʒ�%��"�\.RIգؑ��
��|gA3��R]���)R<��t˕!G�\ ��]��\��n(��}u�r-�F頚ί��*z�QJ���a^.]�
kX	���z�z����L�raڇ�Hl�����l�\�j�=k��I]>߄�H��=Lx��Ж�8�n��<��Ó�gY�e>�W-�D��*�.��K�s'_���v����q���Fq���ϑ���Kt��f���\6G�R��4m�M�������+�'���U�(��٦l�I2�N`(�ă۷⬗�;K�g����0n�ȳ�ꆛq��3�4~���Z��Gf�V�G�&uD�'��R�Q+�f�]�1��P�;��	ĝ��=�ء��>�Z���1R=U�+/�LKTۏR�����ݻ�]���x6�G��8x|Џ~UD �����9J���;n���	����x�x�U�}lOmz�jDB+Q���ʶ���$-x
���~���!�gq�SH�T4%�+�F�g��%v�@˘��V��SX�ڇ��g
�/�i��5�ql����6}N�glY�|�\D��M��y���E׵c-�z�rZ���\&��$2�jWl��1���;��94�a��!@�Ζ:�%���p�s184B4�s�X�H�g�G����ܺ$���~���flɧ�#E(-Z�_��uh�c�{�f�EF1Y���
|oS������nτ�e����M�]��,���@�s�?�:�M���h�Ƶ9�l�r|�#��(�����a�n��+�}�^�Ru=*BZ(Ӓ^��"�0ы�L�YSfn�­Ż���X��ue0���1��K�;�M��-G+�L�(>S3zqN��Oԍ��*E�(N��s�� �|3�ݽ ߸�q/�Hs��:���t�L�����>2�����?a�p⽿������-)��(tV�wF�J�]�=D�i���i��K" t}�3%�K�2<t��z~�"�L��K��_ƈ�%U�,=��W<�ѡ�б�e��{m�}]�>�R6E��4��L޿B����lY��u⤉��'RL��޻_FO�>!��Y��h�O��0���j�F�~��t̋��s) �MUd!��տ���p9wȃ���id���ٍT2)�\O�>��S����qs�}Z�[y��bP�_:U�\ N���7Aq-�Pv�����"y��چ�,ڢN�pl��v�r��b�6Gׁ�2Q�����]�4|l���6"���$��Z���I޶��W��q�CN=�l/k�OHM+�xu��GM�Q$u�r�j�3����KP�����.�]� �}:/%˄8Z|��$�b�{��^V>�(g;w�s�f���UQ3&��ϖg�ȷp�2�G�w�]q����\N'��)��V�\�M�=�o�Q�2]�BmY?a:��z��kH�4�����Y������_l߿y,(�NC�'�˽b�˯m˫a�}r"�$v�K,�<�E�J���q__�خ��΃�tQ
a�������n9�a4׋j���������x��t0U�rEZ�|^.FX�fs�\��O�H������v�����,0:2��z��Y�>�C{[���h�e���N����[v��q�:�'���*EÖ́��>����h\��V�-��Y(}~iG)#-��ҠlҤ��y2�6�)�ջ�8*�ܪd�U"��?O��N��z��>e�TP���X'&k������=1Yך��5D��Z��=��x�� [�Nr�Dq��K0�rfEU�6��52�ml�d�T}u�T9�ZA������s2����锄RS��ܧ��R-3�&������� ��it|�wo�].o{b�ʕX*�oU)��;�����])�	e�u��E��N��i9A`# ��P��x��)F��'>v�v�w��Y������?����œ7�n,���߿ۏ7�$��oY�
R��Eoq]�{��}9��~�B���k���m��*2)$�F��`�\��G?�P�4"�SH��}��h�{]xl�ؽg����E<�57 ���%�o�T��j]����_�����v��޼�\c|5�<:tj��B�G-��݌��`'ڋ~-��_�ׂA�W��t�YE�3Fq��Q���xpx����/!q��{c7B᱈�һ��}?���a��}
Y�I$n4�jIr*��b+�B�9�'LPe ������3D�h�K3�RZt�r�\���ez@Oq��e�AS�XC�l�!V��<P�՚#�ɭ��9�S(�q�]	4Ȏ�t�6��e�z�����r��q|�W�s�*��=�v#v�
���
E���#�pW|]t͙��l��}���<Y�ؑg����g�uX��IiE�}\��u�<��D�{�xnn|�X�j5}�'��߃?��)�=BN���vAK��@J��Џ�]Y�^4JM%S=f��69|Z�eT�v�\���������vc����O��K���u�A�B^���m/et3c�O�������������}���bzh�RG�������G��`>�S>��*ƞ�O�,�V���`�;�W�;틸
o���%x����
�6ܬу	����>�I�ۊ��`4�Z��ӂ)B�u?���n��!9{;��[*:�ݿ!][�����9��Ap�Ϋm (R��?F:��7��uƧ��f7?����I�RH�ͼ��&�591۔��T����z�Z{�sX���]X�|9-�-Ac�����"�7���0'�K�Χ�!��G_{���yN'�H$���bb�2I䝛��N5����,�fl��_��@qz����vZC�Q���@kK3�U*9�-���D�4Gܠ�G���PLdWGXJ�^:,]����j��a�X���L���τьfg��1/:]{}�[��w�d�m�xvv]'BMK=GՋl�v8�>� �E����]�Z�UvZ��#�h7mz�Z7��n�T��ޮ&�������*�O�������
�F�T����f���e�mԷ��뀗����D��@o���_���[���âh�p�2�tò ����8U�N��|��2�j���!"bF%N��;���`��ᢺ�'�X�/�@9��$GgbQC��V�sXJ��^۲�p��J��s��Q����G
�CC3��ӌ�h��q`z�8,q��}���\I�A%��/���sr�N������n#{�Q466�o4���t�sn�oJ�w���9K���L�D��n���N;-�~GR'��m㙉��}3~����VO� �'��*E����~�O	����jX���2Ǧ��'���qg�q�x�{&˙ڷ�B��c��T>��rＱ�R΋�į(u*ӛ�-���:�c-�\*gATϕ�i��y�w܋]u)ZO�������.�_��Z���ä6��Aq$~ǅR�U�F!�����r}J!	'#N��d�Q;7B���]nQ�S+��[5��C`�,j�`�Z.�=�6J[E�"�P��y��&��S4a	�O�ǪjIaѢ;WAy�����e�� 5�F`�c�A."A�/�[n����E��țS|=�q����mR-i�$�ܠ�ו�T8�������,,������C�Am�����`�C4���#�������좿|����"z�*.�	p�C� ��1�M��R������s�i�,L�`��g}֜�5g|���T3z ����T��JVRhU��ݩ���w;
��g�5�o�XCT���w~칇_�g�d�U����'{���?z�(������2���	 G()�-4(��7�Ͻv%>s�5�nvВ;@�@����u��X~���{?h��.�ŉvtH�?���:N�1�~�����I���E6< �cS�z�lE۰�/��X��R���6�nB�َ!�a̑���G���-,��]��
��LNx�6;�h��`F�q$I̕�Nհ�IHh�ߞ�sp���:r�b�X6��]�wόd����=�`+F%����^*��)��@m?���7��[/Jzz��p�-��6��&� �_c���E��^Qs=5)�o7�L�i(��p̅��.Ŀ���X&Ur,�'h̺P:�2���Я[�`HF�"�H����AA#��i��6�X9��G+a��,�5=��9����*���?�Z��w��!�}�5��qi�����X�;�4�{	z�4~��)��o��U�[fʍ̀y��@���yB�7�aŊ���Ƽ�&�>��P{�n��S���ud���8�
�P.�s	�8ِו��SǼ �Ц�.�ӭzV�0���1�&����Ջ�crq��2�w�9>��8�?��	��M�>?����es:��{�ހ�;�I���f6³gN��o��׿�3L�x�����^�'�� 2�,a©	�`q&H�X:�#��FhXr�Aq�Tj�M��S3#2��Wi#]A�{�	8]	�Ǯ�/{)j_q��,-����h'�m�5��Y��h)!�>��Q���8�N���Ud�ʒ�_�O��)���|s���@���1<��il{�������F4%,���0�t���Μ9�����V��/C�����6
�Kרh�)�ڥ(jv�F�ro�I��%�SB��u�N����^�f�%��G���9�6��(N�M�Z��,cONֿ�OM3[�T�AB����=1Ʉt�a=X|e04�;^�Vw��1�*1t4�q�89-�JȾI~ziJg�e˖bM�	ԍ�,؆8�+k�5�
8-�/Y��8��y�)��$O>�Pب�����@���,FmLU�!��RÒ��+0y����xu�MG1	#�ذP��hx!��A����=!ol�_ك3��~ 3��:�uK�A�Zqo�w�V"���Gq��	�k�����w��#hV�c�`KB1I��,��Y�QP�j����q2d��,N�#@S2�.����$���NN&���py`�K�2%��3G�{TO�?R�}9����Z�u �p���ؐ����d�
԰��Q��T�J	�d�k"o
��t�pċ:;�w�P�	*�J�]V��%%��E^�#���5T�����uj�?�
#D�Nվ�;�zj�6���t�^Ӎ��bP-=��۱x�r��pOi�I�u����[<�i�N/�.	[�8��f��o׸�B2��M<dT��Y�={���d����߭�s�o���O�݋#����+���������1�̒X�����z���ג�n,�;ܩxl���s��",`����J���VU"L�!m$��ʮ�\
��D��PG�xHG�o����u��9E�!��Y���=Y�,�pr���� �m։�RrM�N��#�!�"�9s���1);���Y��	՘��e#��w�X�	__��B�S��1�]��^���ʤ�*3����^{J��,J���'z��3~�HѨt(��9��-	� Z=�dc�bݺ�K~O�vE{W2)i��ԯ�����4�z��[+���?"맥��4�֤NYe�smU9-��I�S�`<�󍋎�̿���3'���ϑ�w�獓��-k�Z�cɖ���>*k	�t#B:J/��yEBq�4x�"�����-�\�i��"��f���b��IX�q_Vly��_�E�~��2���QOe��pZ�fs*���r;{P�bQjЌ�Nu	��şSBK�x����`m9s����n&g�ڕ��D�k�m�,G���� H���P�D-��d�P��-�Nш�Hפ����]��z�j6�Iy���]G#� ���R����ټm�]]�J������d(�p\9YWs�q��4��Ķ�N��o	�,E��I�1��E'S�A��d*f�B�Ì�
��[jL�?���7t�I;7g�h�c��YC�)�H"Ҳ$5���zT�$�~+谸&+3y�v��(��TCN�ߥ @Sb��!���6�߯&��l[iwIӭ�;�Am�(�tX�j�Ťj�'	z�C�J�yP5�(���r
XEQ���%g��T��װh�+��>�������j�4&ԖCl�Y��[��)W'�9����Ij��Y���^d:��C)�V먀j8�������h���;�N��%�X�i��	���[��i�)�xU"j�������E(��q9�Z�DP%8�̭��`�7x�_cW�UߦS��
=:%���$R�ਬ���rz����u��a�Y��@�X6�Y��ޘe��Y#7g}:XqB��<��x1��(
�g�2�)W8.7��g����5��J����#�6���M�
�%^��<�@�#ϒ��u(g���S���6��3���)�vWFOy�)V`7��}�9�
'����,o��������7�N��J�T��.��H�$� �f:f�\�t����A������Qâ�I��*s,ZÂ�$۩�>O,L�!�S�f��[\/x8W�6��DA���8W���z��W�I��Ǽ�i�<��,�eI\X�8DT���v}#�t"��%d�#�s��>=/5�)[���BN:א��~��T#�F�MQo_�\ R�o�����ҟ�\���$�I��28�"k����u����#ŎV���m��2n�I�v�Q|{4k�XB��P��
椵Â�>��4X]ȿ�d���![sfqJ�8o�WE3�˒L'����-y�W�[b�g�JӂO��(:�2D%�˧�P-4�)Q������7?s+QD�سk��TJ1���V��v=�/D\]�L[�(B2U��p�Ќ#��!���uȮ�Y
)�h��Yr����ƨH��!ԵU|#�l(	+�~(��|t�C)��>  ������.��&��ޗ�K��D�����+���8�����8�;JA����Q���ڊ�v�/�ob|���y-N��KA;<Ѩ�Ws-��-�v&EuH��S?��+dO�i�Z5eSq�9TK��+��d�����
��X�H+(Ǥ�+Y��<.���0:��X�p�'�ص�z�������g����*Z�30͌����º�$�%���
i�ɽ��P41���U���32�aQ]LNP�-%��vU����O���5��	T!���3����	=@��I�ڎ�*�BT���oޥ�E���/b�ٮB(�/B� �����o	����2��Cۋ�޷H�7S~��U�i��&�A#��
^}}#	�Vk��RD�4�!Ҕ��|(�|��X����u��\ڂ��4�7� ��>��uu�&Q����Շ:;���;�ũ][0U��/�
��+*�4��=�����77L�,	cQW֭E}C�w-��s羓�u��<2mVռ%��1(�ùs��cw݊[V��"B5`{���h���W�;�������ɓ��,��\v:fm�t�������jn�v���zV�b����!���*���h��
��"g#G"�ӵ�k�oG��2��R|]�ƓG��=,���SF�Z�=��I
'cP6c�Y�:J�M����8:cC��O��{8�����ɥ��db����V�SB�F�I3�'+�Ob��N�h�3i�7l &���%mC����ѣ��ѕD��*���q�zܰ��E�(����C+;qbp.^�ߍG^��]���+Y�`k"h?��q��݈eO��䅾��X�]��΃��W�����f���kp%�98�)Fa~)��Ԍ�b�䓔�i���fm$�(M�6@�k��c�!L�Y� �$��~ӵr��T/����4��cV���&}'Z&����N��[��ΐ͙�M��CN9.y�O����tf�xӹi�@[+�d��˼�^�k*G�]���Y����k(�[�a�($�]�	�T*h}f�i	[s�{в�:��t]�������� �{z�sZ¨���Km��xEw��=��@�/�3�;K<��{��\y���,�﫮k$��8-��&<��	)��C����%����&Q*f;\���;�X�l�W��1�a*�7����v��֕�fȠ�I��:u�}�"�ss9(>,G
M��ꓣ�ը�u�h�GX=�ٴ�kG�Md��8s��{�����}:��e�j10ǹ-L��N�If�&H�ɡ��մ���bZ J���r�"W�5��!�(��?�+A��S���	����_G��n��	�.�s�^����F�L�V�+�`A�d�D�d9;(�;˶�C�d�16����H:�����8�H���vJ*!R��_�A{c�;	Kfa������&��G��|{}}�1Y�P�bG�����/��e�!6!Y=o���5$�
o�fOoE��Kp�9,l����}ػw��Ǚ* .O(,]���Y�P@1�I�>���1-�OM#�b,Nk�;��O��_z�mO�_���7�_��K��#ӝ��ۚ�4�`z2Is�=����9����U�#4k*�P�~W-/��V�q}�W��e��G�+عc�~?/�(p������.�B"�[t;�-gp�ltzq�L�E#������3d�C.��)�ӹl�o06�!��g�)��p}|�9��2�����%&(�cq��C���=���,=��V�S�,�ZS������]Sv�u�~������%ڌP�z����`���Ȟz�v�T{����ܶ����'�ϊ�j�^�d)nZE|�'�4˱5_��I��s�C��|���w���7Խ��-�s����$�nT["���,�c����*�,.$<�\�+�~uƎ//�R�ʪ�T�}�X;�i�پ��m)�v�LPg	�������ׅrA���J}"�M��t���Y�w���Ǳr�]�_P?���pv$��'ѽ`9�<�u�X02�=�M^:72|�{}�]�@G�
$��%�Ʊ�1�n��i�u(�L����8�{(�������9�N��Ҵ���n��)rN��&h{��4���ύ�N�g:-휄��,�_aA'`���������W8���	���X�?{��uH� ��H0!r�V<��'N��>+;-Y#iiiAg�E�Yd���eRu6͊x?�����?����>���p�u�a뎃Ĺ�g�"��C8��E������nNד��T�ѧ���9���+��*nJ�.,���e��u5��^��Sh��<���<�b�Pu��B�C塬�q��ts��d[�:�%S:����m����ҫ��q�
�̩����z����h���}�谢V
���V�M�<�}�y�D|_���<�çS8���3���/=�__�4���|{�x}b�w��H�c���=h�m���{q�KM�Ƽ��`QXԝ�2Y1^���jl1A G�쐉�H^�r�jj����e�P��)+����Z��?��ƅ��ZpX�?/U���rg�B��s�Y������׿�W��gّi�(W_6�A�-!�?�6$�u�����ߔ�C,����[e��x|������Ƞ�T"�˹,=������T��ɂa��
��p�tR��(�E��m���cA�e�:�fRA�Vи}���mI窿���4=<-/�T��f�k��@�QZ����[���cA�ʢ�T{۞S�C�,!x�K���g�0����%>v��\��Hλ�kF�%����ȑA�޿�\��֯Gf�j���Kq� ����a�Y���OY�Cz��S830�Q���ÿ��>̮r�r�6�J�i�k$�*30�f�u]���������?�]��g���ѥwî�St]!R���NK����'�2�V�HB��ʮ"<�kEn��MM�$[�  .�IDAT$���Ms%�)HM��(�e_k/lt��dϖȶ�=V�����*s�r�Qҍ��H��5�n�w%�/;۪3/�J�jS���L�4QB�o��`�rj�χ�5Q�t�	���I�,���Q&";�=B�El+D��2�y���z{'N�����Y�O�:�6��`U�S������u$�C,yS�d�%S޷2�K������gʫ��9-A�1d��,�d�h�Q�4���H):��`��Ar�;ə��(v�e�xyp�����^��=e�O#E4�o,�D�AJK�*f+��"�jMu#�(�ʕ�X�tA�-re����&�l���(nh���A�Gc<��l v'�4�h��x�G�"�0+�R�����abr��l�dDªvZ'N�D�ǻ� r���Z/)}0^�%�W2o���0::���+�9C�K1��e:3l���EO.��F�n	I�Vǡeh�ɩ4Ho�r�"f�윤�q';t\���<�IP�p;��]���~��t=jv˘/vL�ڪ\����%]V�ºDݝ�ې)~��7w֋�ҿ+rs#���cg�*<�,O�hS�,���x{ʅpa�-j�t�ɺ��d��G6l�~/�[��L��q�V(�!$w��~-�ŶI�,�UP�VOy�GC��A"�"-K��!�]�"Դ��{Nj����ߋ�޽G�	�@�D
�`����5	���HԱ���˕�&9�?Mjǡ�VnUWv�H<5��.%��.xDRS�{�ʏ4+��>�IC?l�0�	Ռ����?���U��31{��+���9�9��1��(�݇Hg�;p`?�ڹ��!��g���6��8~�Xu%[��'I��`��z'?tZG���rm�w2��_zq���slC�5h˼@���}��n�Ad�u�:^&T��%�Wc۶���U�0������/���}�d�᎟�ī��;�w���͜؂̑'�;�Mo㤳O��NU�A�E
�+J��i��GR�[�r�>�?���ʏ��E'�˫b��*V�5�\�8�*���R%9��2�jk"ja��-gZ zJV��A��lߡ����P	F�w �F'�8��� zz�qy�|��P���hTo�yd��7�|�����_�)������/��Qs��{{ۉF|�_6Oi�}��x�Tni���og�(�۾��y��*�	�Ce��"�947���x���>�8-��3rn�)�{�Y\�;�E۩�h���H�[�L�"��j�F�o�}O�ୖx(��9��lbj��y3d�LQӰ���]����Ige���\��P���D�+�B57��b��.�*U����F(ӎjLe�rA}<:Dbse3�[s�&�GHF�s�&a��Rs�B7<����8|�Д��Y{�@�Ě��|zL�r~/��"v��ê�uu^3�;������!�=�eASI�=��d:��g��_�S���7������X�5�ַ�bddx������
�۷��?������^8��#&!P$d7Ǡ5�z2�=���I��)s�#糕�k�h�a����N���ט��?�1�3)[��̗��/6
k�7n$=�Ɓ���j�d�5���������WѠ%�����9�Ӎ�⺸�z}���c��T$�4H�ڄʴ��o2�*ۂ�>�����P�c��1��$5	��x>����D��71&��K/����E|�Rs�C��R;WqG8^����ة�)�ja�aJ����_�c����~��X�P���pNa��i�<-����\)/ob�&*HMc�����)\;3�F�$��K�duXk�n
s�%�i\��*���*[&6���jDUu1R��}�S�f%+�H�tvX$'e_8�[�{��k�Γ�,b	��m��G��2�~��4��e�_۝<�i&�{��.��x-~��uXPߏ����r�}d�]8���Gވ��|�:�b�9-9M.�t�Ϟي��l���.�MW܊��� :ыtb>����W����8x�$��k�,oH�R~k�G�E��C*'e�)�(5�]�3.04�puat:6_F���ۑ�&���RYŨ����S]m��S��_+�I�R RB�v���W�93��9ߦe9�r{؟�:O���W�{���x��<����pX��8zo�I��-�q�h/���Z�xG&9K��^�jT�?���+��܊q��I�VS��>�j�rJkK>xY�*�%�yY�a5j��&���M���3"-�#-c��$S�<,�.��	W_?���
��������8B枘��,!GX����yTسm$B�K�Ə��@P��S�	}>�g�|Mʸ��\%".ƽS"��"Ծ)Q*8>��/��aM7"R� X�ܝ�i�MP`��G��_=G�)-!&B���@T��]�F�b^�:�nm0�?mn�ѳf�;�8�dߟ���$�j���F#�z��&A$�Ը>^_q��DX�drO!b��>�1o�6%x+�?�^����nH���������^u��BYd�8�r��P"��\��r�::6��g��Sms��*����,��ԟ��h���|6�����,_�Xm�� ��
�+�[k�?�Y�����*2&\�����ޟ�X��K9�TtDCO�)��VRb��L!�f+;{��CiYl�`���dx��9CEX��u[�&
��+8��k
%����̙��ـ�)d'1�m��}ػ��W�zE�<�I!�������٬��NK,Kɱ-��ٜ����ᕗ��ɵn�`������WS�ȳǯ]9���}2�������46�j�m��ʫ�;y��mO �ArM��e� CQǥRE�)�t�&iNPD��4E�L�ث\��r]�3XnK�QC�5%W�ZR��X�馄Iyo�L]�f���*Z��u$��w��	�.��X�5d8-��;I��C���5��w?qV��z�J�.��!�Yׅ�};��������R� G�L��E�����<~o[9�����dhx�H�Ť�"K�Z��e���e�(F�S��^x�"�Ee�Z8^�Q7�_I`�-.3lt��q��K��9����1���Qq4,�d�Q-�$�x���L��r�,�YHLs]�L���sT�q��g�J:��o���ν�P�6#�y)j>ĕ��K������0ۄ�7���i��%_�W��WԢ!�A&�I��ɳf
'$RB�(�n�H^�!8��1#��cЍ���n.6�r2!1��)l� �j�trJ!�aՠT*]�-e鴚�tщX�!ny�����R�A8w'�k���� ��]	�s\�Gab���-��u*��jD��	}ELYE���,u�B��ճ�?��=�I��,מ������w�M`�JY���h�r8h� ΟO)��_��8l<t��B\5}��"�nb�ݻ�ӷ`u�K,^��G����QlX�����l�!�9I�<y�%S9L���ċr�Ps��j����-q�Š��J:
Y��&��؄��p�퉗��)�&�_?W;]U��k�nҐL�/ QeE��T�����N�v��XR��|��~�����SQ�ZP:�b��0�h(�`�^K0�;֋�'�#�f=�J{������ɟ���`㤫h�ɔp�l���j)����;��:u�c��D��y�y�5=Y�JS�
kH����Y�{O`|"Y�>f�LPwtv�k��2����(�� H�<5�?����H�SNKmO���0�G_F!�$� ���R=Q�/H���n~0�Y�"�*��/�6�"�,��#���JP�	"�'�����N�a�$(ۑ����US&f�|�Q�޽�׳S?��=\rY����b�[�>�qn����BRЬ��RpΙڅҩ��g�(����.CbtG�*MGtz:L�iI5���x<�ի�A;lK�SI/24�}�����s..����liR<��q�k>L,����+$i��1�tB�����F�&J3��D ,uo4�#Jw���a�kT�6��C���Gb�EjX3�䌮
�ktt�vmǅ`Eݦv(ԋ�"�J�q!r��f�ҒB&��`s��9+8�x��l�IJ*�Q�0j��j�Ƣ��s�^������&4�'04<��<{C5{f�I����_|�FE������l�flR���x��-�JX+�}E#-T_,��QP��L	�o�auF5�8��Nq�.���9������%��ְ2��0>f.rYg��c�����Y�28�(=���7GH>�ʕ$j40�S�ɨeʋ����҅eS5������D.��T����~db� ��Cy�qr$������x:U?&U05�/�Hu}�LMQI������%����DB���pn�7/*Q����$J�9.�*
@�ޔ��VzhU�"S��k&3\����X���P�*��"���s1,�Oh���2S5ڼQ-���q!���N��������¡
�Գ����NE�ꤩ�qM��i��"rI�-��T!DiY%��S��Z�A��k�K�ټS��츬R�� ���������a�lJ��X,gX�w��tZ�0������Հ ����&CKUMH�N�0�(���˘�f��7�S�]������g�c��P��U4�7�����Sߑ��iUKjG�Wbz��������_���C�);�)�����'B��"n�HT�r�=�Y:�b����i��G�)b���ƶ/�C)#�_.UT���":	BJ�t�
�(�/.�{%+zE鴋�r��:%$�z_i���8���4��=@�E9���I���eJ�����If�m�ѧ_Fs�rܶ�˻���09�\�	�����w�����(a���8*AV^r)�����p�ʇ#�fo�یLv�/o)������:Fq�����$�E465y�[�,����������I|�/�(����
s�D�2����;��u��)��x�w�H6�̴gm!�ԇpb��h�D��.�b���Ihnn&Aa�\� �v����©�,NCwsL�)
&W�hj+�JGZ���lt�3^f� $F�L���vm���d�d{�-5��b�����
S>/
�"2H&S��Ƕc�����=ג���hF��	���(^ݾ	�O	e�F!k�j����m��%������2qs#:�:P�)w[~��t�,Ĭ������������OM�U&Z,�;⭷�T+#�Ђ�~�����%�/ş������.�]�G��9��Í�ۧ\?����ո�g�^?s��|�i�/�d>}����"i�����K/�Dˮ]Q���Z�9�a����w�wX"ҽ�ʫ���`޼Ҋ����������xn�#�B5�U̪���̖��LA�f�h�F>�����,����7������#����|��j%Z[ҩ$���9X2ͬمek._�?���X�<��^��.J�.�a���b#����Q7��z:��kT�������Oc�ʕ��G�¥�����yY��e����U\�n=>��4�B��-����8x� >��O�Ά�r����m��_×�#�����B,�cт�(���w����A}����ޕ�Hd�!���^���)o<w�k o���՞S���=�?�E��Åw_G�w�e� Ւ�EQ�)RE1�lkKN�g��QH�/��4��9�4����6�	>ˢ�������t~H;1�+�U��2bV�C��|/����+�-�{�{��~���>zM/�X�m;�#&:j����E��bq�N���ѶpêF��Ű��K�!'�K����ݟ�7�����l'�]G�"�⮱M^��B�ǆ�f�p}����&,^�����e}�Qą�'��K؉�@�8o���m%`g͂V���D�tO6��f{�Rp�Ӿ4-�k\2%����Ţe(��F�9���"#�ϬtbA�Ґ;�e�j�>D���Lt�7�)�-�iJc�jv�-�êU���}�-����v��5���V~S@g>���X��� G{�q<v��^���w�'�h���>xy<ۄ�}�Ә;	�y�9Y��ލ�|�H�[�c�\��`���#��>��������N����F�ܹ8��K+��K�j"[H&'0������� �9�Tj�
;�V�Z�Nٕ�N���:#epZ!9C������,I��к��+a"���A=#��s����L)LЇ(�����% 5%��� �@�}�^>u�d 5;&R�ŋWb��UD/4j@(ʨ�B��f���Y�;�|���/�G埿y���>zy�p>º��6_n�;pL��[J���5?��Y��_��jL9�l6��� ��1�<���V���O�i}�w㦛nû��JOO��)ĳ�A�G���M�\
�d��м���%57Џ��,Ň��©��,�t�� ���	7�_��MZ��CMt�i���z���Ʊj��뗀N�Jo���Q��3A��H$�dN�� (y ��㓍�͒��ҡ`1�S0%L�����$bŤy�zE��JiEW	THP(��)�����EkF�D����Ϭ����y�f���~��X^��:��ʹ���\���8���k\�p��TaM�f�����u�Ǖ�����*_��v��Ƈ��%�'"���U|t˃l%�mF��pZ5;6S��Su��qUm��"jV%�!��l)gU3�J�׸H R���il�>l�ځ-��L>#��W��H(�ڎ�bÁ�XO���	�'�f����M8�hg&�̬_�rV�)?,Y��a�"�n����U�S̔�*ע����pV=�I��wI�Q��Q�Y��.C0���|ڐ`q�ޭ6��V�;�u\>Qu�2ŕV�B+CM��4\�f��m԰�����`"P��Bg��mq;Ј��l�ZTJ���>ӺӝK�tհrv	�{%u]�r����%�9֜���s}#N��Ul�D-�}+yS-�!
]e	���X��
=����TT�E��\����z��;j��*�|t:)kX�Q��WZ�{*+��J�L�s5�l�l����m�t�5�E˪e�X�4!n~6�3�D��Y1��y��(�*�ۣ��sJ��MI�CJ���秖n�6�oV1���k�U��P���L
Q�
�[j��($}.�8C:_�(�
���	/0Z�3���ĉK��btd�t
�U'�9<'$�QI�4P�ѧ���U{��:2EU�A��2p�S�	X��Ù��Y0.zU�S�p�\���P�"V��&Mhv�����K�-ÍW�EOs��v��:����P+������ǁ�~lym>$g]	a0T�)�t�|҄<H�ԘV��eA:R��4z�p!��B3�*Nw��C-�*nUS�(ǡ���Ð���.���K�b��l-�� \����BN&��v����sH~w~�����#���a�@�)�U�G�{r�����G3X&��>X-N9��ù�w@my�����^�'�<YU8-"���Ş#1�����?�����\:Ꮅ��e�%�)��������t���=��o�����Y�ޮ�3��@�6mC8O*���Sb�P�rp�j5VA#u�fܦ��r����?���2ˎ�w(gepZ��K=M��J&����?{'��2�.� ;Q�]1kh�Gln#~�#���q�mz�f�M������d�1�%N�a�<E�`k2@��f��9���f�>�ʁ�,j޴�o����iIV�Q�BnX���Ư~�&|x���Y?-��,�}5.�o�:�楏߽�~J?�n�R�qB1�0�L��P��Fa���/j���.�;x�W)s����L���2ꍍ���/~wm\��ײ��LLC7�m� ~c������,� �P3t�s�Kl1GH*��G1٬]��o�`F6����VaJX+l�2���L���:�R�����"�uhZ|�99 ;C��+��/�A:5�g�{ދ�"p�(�{T�ruE@U�K%��2
�dz�οa.h�tp���H��>���F�䡸��<�N�
Jُ�FԷ�{儞E���+�{�~�<y���\��p):��l���ci�f��E.պ��H���;`6qz6Y���?!�n ,.��X���X=/�P�s`M��~�z�_���|�J�\qtI:���k\,�ai���xf�ZMk��]�N�q�r_�� ����fK ֭[�Ko��-�l�e��:g!���y�s�!���D��	IqS�Ò����j�����̥nԬ��uZ�����(��[1��)�I7�j]�˯��m��駞dn,�@�n5T��91��8�|&0e]s:Q��1˶��щ9�M�������nﴻt*�>�o�76oN�̭��4�{r CCC$�w�Z�HK"�[ZZ�za=�M�1������/#�ŀQn���B~��l���+�Zο��Q�-U�k6v�5W�7u�y@�@�hϞx7r��\q�X<p�u���:�v��V��wO�~�e��*.u��uu	�ש��8f�f\��s�v˂� ���1F�a��x�AZ�dk���Xa릛nƗ�������L�I6x�e9jVڊe1���&XcQL%��ƪ�W�ȉxs�۸�L��ӽt�簰����f���9/�G靰 ��ZG)ћ�s�}�S%������� �.�j�Uj��-��Y�I���}����?��p1ZU��-E�i�I'c�p���ǡC�n�׊pߡ�=�mF��L"S�XRy�f]j��smk�\�a��&�em���)7�41}��5^�3����,jk'�ұ�Q\lV>Ғ��gB��/�w�DG�QyXR�B�j��A�r!^QE[���@���k��9��+.E��K_pE��!wi���>1��z1.��O���Z�6ۀ#M7.�mm5�0�744���;ފ����	8
��0�5�Z��y��P���)͆�pZŭ������p��M�8�;�G�7ґ�x��� �:"��;�.���� _sX����r��sǵ�sϟH�M�B"e1Yˑ��R�W�1� r��f5��-��ǩ9�V&���񓧐?W8{��6�ã��;%��7J'e��RB[���Z��2pZV�i]�V�9kV��O�X����N�M�e��׉=s&�b��=�A��������r�Y�ٳ�4��+�<�f%�Lô�3q��=;���k�e�Vz�8��O�ڎ�*jX�\�4�H3�%o�h�6΅�k!�sWiQҝV��V���(լ6f�Y�H���u�vp���B}�R̦��=���~~C��j�.T��3fi#�s���B�Q��f�l���&c0#Y�R�z-|��X���S,����M����=��e������8���k�i�]f��O�~Cב�L ��!�iω�PsZ3iԷȒ���l��4Y+i�?!��9�Ç�[�W����{�:�\��M�����O~&?ȱ5$�*d#��Ev�$�.���},]����f���7n�Ʉ����[��` ~5ޭ6o�G��h��fMk��\׽�7�&��p���{��MԶ�A<\�%f�r�!x�����[���: ڶ�df�6n���ay��)q����3�c���Ā��,�&5MH
�&�c�f���R�%�Y����Mwxc���!Y��ss]�~Fo�p�N�b�T*���A46.*��Cr\9(�z!.q�t�����t,Ų�������؛��G��F�4a uI�����s��.BM���>ڬ՘���y6�{sCQ���9�� i�ηԣT潏t��LMƭs#k�#w�C気qd�Q�r�4��ٸ�)
��uۛx��g�B�hZ��? g�$��?����i���V�����I��(�F����^�U=��J=5j�sm|=���t|1�u��Ɗ���^̫j��+�n�c���l�VQ� �*s�#5�eX��PD(bfN�<;�	����o?E]�#���ԯ���̤]١�8����v���~N��)u�o�N	����C��/�_�Af�,K���=�}���S����k��\��!��4�D2��P3�J:-����Ox�L=�l�����c��S���%��%:��Xj���	����x�7�C*�'�^�Mj�Na�{��#C��i�QV5��<�zχ9㧼��vC�qR�q	���c��kB�|+)!��ȭ��u'�� ������;���̍X�b�K����1��ڃ��|���'���,a�DZ��!�N�w"����n�ս��kKS��:&f��KUZ�Y>�&�r��x�I�f�U��3��(�,r#f璄�i��/�L��s/~�#��5-+��2�Fv4Va�[�fGzqv���s�?~�U<��㞳�Ȩ(��3���j��9��>Q�'�$�x�ơ��qI�FMs>�k1��ւ5� V��h3��8a>U��,j�IPt����6/��Z��|�l�܊;�� &���k�Akd�9��[Erǻ o��$Ύ��s
xf������;rYe�r�9$a� �2A�tD�+G�ғf0i��W�fߎ9�g1�+����yѼu1;��+yg��t�/F��I]�v�׌R�D'��(�f'8E�ˎb`` ���=Z����H$��b�i�����#G0>>�LF�|����!�8��׈,��Jyb�f-�=�V*�B��H�'��&TS���g��c��ND2�ˬY�Ō�-���Tĕ�-ĳ{/�L",�iD�'i]h:�����LՓ<G�p�hO�M�KX�OB�;R�Pm���ҁI�;װ���x�C�]I�'��4]`ױ���,Kˈqu�ε}���#��{�ս�O�)X^�A,o�X2�9x��%���7\L&���e��M7݈��~�"2/s	R�p�H�L�l��(�"�cK����S�hy!���eGD �L�����]8!�qq�JI��zC1���?�%����[���X:��?|��H�øj�R��e0�]���XE=����0&&�%����Ew��G���9%���zof	�;�7�J,�Sϼ�G7�###����'��>�)z^�b9���}������~(j��͸l�&�5�KFQ����TVá�"�L�ď��c�B���R���ۏ����KҥP
�ֲ�Y���1��?�+Z[[�D��Ԃ+���*7�J��)�	NK8�r�aN�j�?~j~�y�~��0/";s�46n�Y�/_���s7����_�ҭ8GBn�j�ERsy���YU���n)�\v\V��耣,f�:ڪ�(κ�:����R�$*�����ٽ��8::����:�V(�z1{1:*�FG�b���>,DP����ǫ���m�$��@#��i�w���LU����d_����f�q�
��g~���K{��@��}}�p�Uk������������رc�o�����̎�Z�k�ΰ�<���;����ϵ7�ꪫ�կ�~��⡇~��լf��&�D}��ٳgp��>,]���-F4d�N+�k�ƥ��FSS<�-[�ǻ���^z�Y/l7D��۹�'��ݍ�M������.>o&�w[���º馫���Vt��;X�I���P�}�Yl���_�z��c�=�����П?~U�uuu�ꫯDgg"���������+�<��k7���?d<Q/���ჸ�o�����.���wy��z�����S���~##��Э���sX�r)�r��X�hQ��K�b���樂��l:&���'�z��	d2Y/ڵ<�U����_��;v��G}��)/F�;�O>��~/Γ��	���?�?����x|vU�.d��r���ǡC찄E�/����ÞS�h�V}}�f��ڈ#GN�둑	=ڇ%Kz��gUg��#D��@�C    IEND�B`�PK
     w�O\j���  �  /   images/85ff3ff6-223b-4d64-b6b1-3b6b2877ae4f.png�PNG

   IHDR   d   �   ��6o   	pHYs  �  ��+  �IDATx��}|\Օ����M�Qo�e�c�����%�gY 		����-)�J:l6d	�lH �!tӌm�{���ջ4�h4���sߌ$[vH�l���dK3��{�=�\����կ}/��24Mß3��4�?���^�b���{���0s���O<�Ph������f�����M7݄+΅������U��n�O~�d2YCe��'DO$����zD�c6b��o�@��`c=�u�LY#+۔a5q�{[[;!�f<����>�r%���L���{���Db	tv� �H��!��sxr�W�C��Ɣߥ�����ŁB�1ݽ�DMcG[Nӆ�lܸ�y" ���,�����1�u�p{�H&��߳���ּ���e�?�?g$iSϨ)�g?u=.��|���=u�5��Ͼ,�XLja�a��D2�+.:���M((������q�p6!�ߌ���I��S�����p�O��O�nީe������߅o��g4�?ϫ��f�V�߹q2&�Q�/���P�(�o�-d���<x�;�V|�k�v2&�+��$���<�c\~�����3��G>r��a����9�f\����.�g���R�u�Ϭހ��h�SAc�NX=c�i��|]yI �C��}�=&ڥ˖.�_���i3f�nF%����)8�)�j��[x]�t{
����78���c|�[�}p�ڜ�A�XM!,\�C��A���FC����q�`Mjhh�u]��G�Cy��!a��*ؖ-[p�W��mظ	C!�lo�c+L�w��S�4���6m���>a�٬i�徴ڬxj�˸��͘��'|��p?�{�x[�O=x�nظ�W>�w}�#'�0ǯ~qFFB�ee��8�6PXH�ƛ��}��-;�#�m��wn���-��N�.��:�۰�����s�<.����]c$G��[o�ʗ6g:L�*yǞC��S���^�~���sPR�X4��6��?K6H�q~����a!�� _��w��܆�/��U�He��߇ǟx�m�E2X#�1����c�}���~��x\N��ӈDc� �F�����E���>",���)g�>cya�M���
Lh��������>Xf��j����$�����1���>�8�-������,I�����6B���!D�\.�1#�N��H�Hd�Ȟ�Bq[Y����h�?k�h�����B��c5XTm�Ń�����q��q���geS������?��t��HG�׀�9��5��g�c/}k�X�f�$��e��6�X"�+{�ܬ ��Ҙ?o!ND(9�����5�J��u3jq���,���>/̀�4�y����7��F`Ѳ�jv���Y!i�INz�8�ޢ#��ِ�3X�1�&�4pXSH800���O6{[[]�`+�X��[��[�o��BeV��J��SO=���zԔ��
r/��tD��/��0#7!��@����`=<�'���񷮴�*��o8-�%4+�VbS�����9�����[�q�%�'���C�&�`��hh�	�K_�V>Q��Ԏ_:�|q
�4��F�,��P ��e��aMY�=��{��l��W����
����0{v�df;&:EI�ԉ7���jޯ(s��&?�8�sC�����:��[��<���O����M�N���U����8���P���p��s����H���t;�/��x�����IZ�n$a�Z�8�н�H���Y�)�1���."���T��(/� �?�H,���yx��/�D|�\��a����s٠[�z%Q�㰐Z[Y�E�߁i��h$ᝎ�a�ϡ�L �u[6%���q��a)�����ain:��&K�@/:֪��o[�`�Ť�g�e-.�p�t�ȳ�\@�`,�e���/`��f�t�v0��n ���Tsc$�2*����b/~��K�+��ϟՀ�;p��{`ג0t�lx��#�d9[��i��߶�"�t�q�N~�ّFd�@/�C�k���<�d6e1��6�={&/!��:�]�4�@��Y�2��r�L�a��I�v7��)%1a[��T��&�#m�Grv���}�}�!����e�V�mQķ�Hr�Kr VG�nF�3�h^2�D�"�$�0�ƈDm�d��A^��'.��4��դ9j�v���D��a{ר�A)d�ˌ<vuR���h�7	�N����ޛG��b��#�)V�"¤Qx����\�Q#�P��y���}��',9�ݝ��opv�e�E���oR��1q-,?��|��U��˱i�Z[�����c��a��X�w}��-���K�� �N�k�ʶ�Y446�����d}z�N�GtFkV̮`~Z�u���DMm��x��]�u�G��S�����U^�s�83gW���2<�6�Wwt�&����Ꚙ�YCs�Z�&?�`Wmn}�QY'~i��`#��`��Y���5X`���I�[\i��� \Z�/��ۏ���-�M���</�e��+P��6�ٞ%���{�X��N٦��ɞ��!���u�!��|�������d�	о2���~��ݍ!��v�!�Z]Y����������d�t���>-�MM1�pa7��G�J��>�@ǯ�ft��7q�ؼ�Q�s�T�cKcoK��CǉTY'��6�;�?6�_�I4�xp�c^jh�	��@/p���Y�;�,���-���X��u(����7�F�[��C�8��C=NYdG�!+��j�U��˙��=N�7^;\j!��q�/�o<�D}s� �8�0If�EK+q�r;lg|�����1>7�_j�*�0B�Bt�[��J��8ҝ��$����F���H�,Ԣ�kK_?�2�����ڇ�S��j�K?����r�g~������]{�/w�&y&�N,�+�a-�N��"�i�(�l���0��,-���hRK�O�/�w�5p,�w�\��64�E"s��!FYQ��O��b8
g�S������{�����]v4)G���%vX}����c�.ƴ�p��S!D����p]kȪ�t>���Dc=�0Ŵ?�7	�����c%)�Q�-#����WE��
u�`�N=�i�q�4��A�N6t��z�F�>h{�zuI�8F�U�e�jX���^[�En%9��4���2�Q�BU��B�9*�%�&2��vU��F(�#O�����*��ء�AOȂ�0C�x�(k�}�c�������b(2l7�ĽJqu��b����������$�G�f.,��8����P��	�!���v�9t��
3ņ��l���|�4ޱ��m�04����C�_�LI*$��sd^|黰as��;��]���2��N'�����x�4v�"<�X��1ٗE�/���m�����a۬�T."S��jʧ��ZQSY�/_Y�@u��j���Vl���'�� :U�����kr��h�䞉�}��8��9��k�Č�\1�Ol�y��rH��^���{��[��t��F'�q;�n�9h8ɮ�� O�C���2dt�I�Y�/O��}����������'C#I��9Ơ��g�h8%;�G2id4% s�,���a�xlsY��9��Lfզ���t?ߓ$C��g��{F��J�xE�v�!zOq�ڕ�{���X8����{�4�xn��-��RT�B=�d8�g���v�B�ܡ�S�l�L�եItp�G8!R�Kr!M��\vj9
�vl?2���8Lɺ��Lt{^o�r�P܆��[x���?���]�/�	B����a��l�nd�4<���o �T�����Jvp�cJɀf���B#r,�A��Y@�H��XZ@�t;��]�k<n
	��0F�î��R���),���ABn�D�X蹰�����,E�8ga
�];�"D-=,&Aj���4&OAn�~&.Yh���߂o�އ��{2,,K"�"E�����|��6�����>�>�';�^��p�^�������! ��j��u9������V�}�	A����Jv�&�4=����e��tF(��,���V��r�%8����	���7��H���f,Y��~o��u�����!�����),��f��yĉ,6�A���C6l��9���;�I���%~X���S������sWcW�Ü`��r��&NG����){=��;�D�6�'E�YL���ǻ�K;�K��Od�����9 '�W
c���٘aFR��3Y#�S�U��Y��=�Yi���g��P#i��U��o��k0U[��J��\]C���r���}��Z�����#h�
T�7\�;�'0�!e>z���w���x	���i�X��7k��\P��?J )	�ax
�u�sh�9�bx!���`B �t��v�:� RN<Ų�߼�-��*@�;_�cd�$�ziyA�>ެ���ue�ݙ;�M��
FB)м9F�B����'�Вb7���a�ע`�kx��_�k���J4�ٻ��w{hC��e�J�D��5���0�hi�n� 2�oӃ@�hm@c۠����[
`$D�$:[��?7�)�4�e�3p������Â;�I���RgrTf��P����<r��'����),wo
3!�������h��[�ʋ!��0E.�A��kK 2�
_�#��Z�c�ڢ�2�?!*@�i_n{)���>�%�CGpǪA�7/7��ȲXmk��3*Q9s��Z��13����/��f��<U(/GN�����'ޱ���K&O~��D"�m�c(��a�͏'vE$h�8�s����涅�[W�������԰����Q�5��~w��}+�cՖ"⻤��OZ�q$'�0��Pt����R8��Owg+��� ���K�bZ�P(���~_���-�hm�M��C�V��s%�$��V7ṭ>�Cc$�Ro3��˪�aq��8�:�-c���:�=��:�V��.����!0�d�k!n{`-�lk�뉩���,��e7~�O���;��n�ý���*���r)7�����5���x����	�:c1C��i�!�,#�&E�����n&��̪B�9=�ђ2�\n�&�[�:�P�S֪�Ӧ���8�sg�p/�G�2	9��������6�����y����Zƴ�����Kpe�����]����.��"��%�.��p$���zz�g��_���騻���ì��ќ1e���i�`;���[惏d��,6�iǲ��$��+�뫰|a9G	>�߀o��`���|�x�C���o�a؃��>j�}]�ț}�,J��fp8��ܾ�ϦM�)��#���um#1)=4#���'�p�lR}��p�!����[�I<�#�Y+.]Z�3���o!d�{�.\��	����1��D0�ˁ��\�]�D�ݏ��~��9`��tT��P���>R_����/�F3#!9
aY{ᩅ8uV1��~
�����s�%�z�6�f�ӐL!C�g:������ؠ��@�yćî�����'���.�"����so�!���|�RXs��f�U�K��]73t&���3a!���d� ��瀄*�`Y�0�֜�po�	{F�l��w�q�_�|J�7�܋��OK+�?�I��VZ�{��R���OӦ�(ȵI��M�����](9�Kޙ@�Xs��M�U��][��������V�ĝ�k{����	�>�s�>j�=��7Tb֜!"� �#����q�fSɑ\	D$�����P;�=�Exb}�2MVb����~����7����,^m����]�Ʊ�!�] /l8����r�1�b���2x�G#�@ʑϽ�C��˃5h=�H��,o�~���`B��������Dcc��܊�Y�x�	�\гa�O��FF�"��F&NƵ,Swf=�(��V�]���G���8G-��b���q���p�W��Y���2^�Ҍ��`�ZSe��~�Rx��឵�p�Ӈͬ��B]��(%#a(��ǚ	y��tg֗3�:��Y6�u6v��]^��.#1��"j�uy�r���oq��P!XRq�$,�چ�d�ϴ�U�b2��_%D@�V�p�g*�`2��?Je4,�?^Q�gk����L3-t��5�WEM,*�Gh��t��&Drj�ߺ�8�P!ZU���ፇ1���`�Y�2q�]4�:/�b���F�zk����y���uu����`n]��勷��3��� n5X>(9��y���5����Bw�&���`|���{��s��^t9������,��1ӫJq�?c�,Ұ�ոd������)#��d�\�ȃ93J�0��$78���=�ދ���=�M5K��(����U��Q�H��q7�5��<x݅>��ŘI�^XX�߿¶����8�pb�y�
0sZ�e?"�:�pU��g?��;���\����Y����q�"��j�J��ka]	>q��E���J�uo3v��[u�+�/;�n,�����"-j�ȳ��H�߬Wߒ��͌�J�:6�7����C1\�Ձ��?��D��9����T��|(OQ�pqz�a��voa�a�ɡl^o�L�KA�"�烜t捾�H]]=��燄��v<�U{3�Ǧ�r��ᆣ��C\{�Vx-l��kG`��8q��B8'j� ��T!�/�&R�EKwhR��8�k&;�W��n�M��xyyz&�`����C�GZz��z����wn��VX�#ٟ�۸��z�%�-����-/�Nr�	ҝ���Y�_d�Dc�$6I"�I����`8o��U�*O��-8�V�GRh単߰6��7˖�:��]H>��-{��D=9;B���A�[:D�]�Cc}چ�敇ky���&�t*�%��p�X�k��.�w�+7�����XMK�J=��+����Ϝ��n�Ïn��
��Cl�I�$�� �LS��Ǽk����F
d�;
ŷ�G����*g�j0#!�=����C�=�Q�K*�,��xˊ���	g�>����9'�1H!�r�W�YuN�K��rBK=C� ���%��.���k����'l
+5��W��pt؃�#5�{��]��x�"BƸa8̆al]�*�l�7�l2��,��p��3�sRc��Վ{_h�D��c��
��)��p�uŨ�}iYX>�E�u�{es��"I�L)\�B���ćo��e��4��lb9�>�����;�u7>��.76m�B{[�dHN��e�Ω-�|ȍj�-|3qv�*R�k��&'�����γ������P��,��G�G���qT+&���&��(-���[���e�$*����q��-�/��8��3�����^���'���n�y���n�s�{QQQI���lf�Շ+ߍ��y圯���!l.�48�~�8L��p׏9q�/�דP_T��U�U���k��l��B��� n��,)��B�}�T^������:)�OK&�-1RaB��vL㙋zk�����̱~ ����v ��&k�L)\�@�e=d�{%xe�IN�����[�k1$�D׸��pB�L�_�a�ڡ(��`���0ܕ����;����|SGG��;>�<���돤��TX��L�K���y����=ͣ��o�X��#��������:��W��yCTU�𽻷`�:�v�?$�S�Y�;�]��m���=�X����^"��(̻�9��NT��Є�h�+7�.�����5�MiGp��a1c�Yq�If#�4�H��m5�V�>�Y֛�JG��p8�VnB��~k� n~((�|i�A��m�C�J���6X,R��-�t)�T�d��X)�7g�����}���
8�K�͟?�gz���C�o)R�P�������Y��ͨ�7���0v�p/���n'�*�H��>����#!i�On�t���J��0t_��h6��[9�w� `�c�кF���s���\!�+�ҽ��1�@�v��~�����O�?�g�ב��#�q�S��K0�eJa�łL�i8����&?J����'__}ű���њ�)�o��,Շ�N)Dc��<��٬��}+���[Q��`mC~��av�O��t�͟�߯!��}�
f���nd33p��M��)�nh���Og�(��7	2+�ձA��?���7;Rr� n;8�7�X�K/u`�� :;;L�x�ά}ɼr|�J��]�������g�>�4i�y�0cXq�\
��ϻA>��,o��>�Ye(D��G#�;ݏo|�
%�U���X�u;[��sm��)��Ҁ���y(.���R�G6X���9k=7̬w��Kf�	�ӡ/��|��<��g(�y&�"����'�aăd���b,i�&3�Z�p9p6�H<���,V�F��.�n������iD��-���0����_���bݣ1�Q��!_1��&��풒�S�!vK/����p�����}�xpS
���tGM%Z�Nx��%C1_�<��?T"� 2�0�z��N�`�jݾ�l�L�+tw9B}Gq��$��)jE:�V��{�x�Yi8;��H
��6�ew�q���zc����^2?�K�\҃��>�9���d��y���r�P_�s=�X��޽2[��m*�.�C���tlI��bC������8�/�$;�B����]O�.g�4Y�GZǝ��b�39�Kl�����(p������߉M�.ܴ�BE>Ba���u��4ۻV�̼��x˵�쐜�Y�:��l�ѪEC��_`�K5��Dq�|7n�֊x�48|K�-2[��o���lT��x�Q�w��\k�,��l���f�+��uL�z2���~��N�SG���0�h��
)G��a7rGQhf%�&�,E�V� )�#,[rS`��O9��u����7
���ݖsu���\3�8m*��Ć!$HU��a��/A:��0T72t>��E��r"G[�:���#�{�#��]>�GG}��n+�̹Azሔ#02Z[[�v��NG�x
�T���ى��}�� ����Y�|��ѣ��9b�$^�Dum7���]�Qp������V\�L\ww��bgK~�T��I�Nj��l�4|����I%���Rײ���c�@GbZ��cE`h7�ߏe���ށX,"*��߃����ɱ�s@������x�{�UߒqO)��yM��'�M����k����U%ɓ���<��c�5���S9�G��ί��wz�~}#��������Y6�_|�ޅ#�p�[s�����#S�YҚ��9�.�}�ԧ�,,�1��d������j�\�:2��עe�ɕS�i�PE�5e���?��H�f�	O��)Gچ0�� ��̳�{DdIme�����cX<�L�ʥܚ��؋�Bup[OH�?�& ���h��֕����p�}Hj�K
Uύ����1gZQ>���-x�>b�e�,��xʍ�jj��l.�u�SBFw��&l�ĩ����uOmr����2c]�F��{�C�G0�D<��*���^�Kg9�Ȗ� #+$��|��4A�9_`�H��ux�����/\�ӂ`8����n������ޅ��������v���m���/G�cE$��'��>����s����qQ��/�ԥ�{��_���>w	J�N$������5�/�{ϛ#���m@�问���� ��+��ɉ<\�da�"am��,��� ئ��n�殢ݸ�a;q��'�����v���S�xg���8����o�%���J^�<��U��ӎ�/��2N�\r�i��ovāt3��c�Q3�)x$�V]U�S���$�R� 	�~,=c���C�D�`�"zf��q�=eeI,Yrt�C�V
-5�ӗ����B�,E��ϝ;C���-�)���sa���#��ӗ�Oԑ�bWͬ���"��v��C;7�w�}�}��$�dfw�L��l*�h<9���x
a���A�=X���Md�]/�!�N����ǂ���-X����v5����[����N�#�B\6f�CM��a?ZZ�*W���h9�M؅�E�)�`��{���B	�������5��p�oby������|`71���p+M6�`k �6��g�kF0�aÆ!,����K�I�;�5���N�F��;��]��R�a$S�M�GP�v�җd�4���p?>�f��)�)��u�H'�*�9蜓���@S�U�i��|À�"����vo;ޱ�^{{Z�hj�.��x���yb22�76bC�hS�䉏ۣ.�� W_�Y��N���ǹ�{��le��6��y`עH.$����q�ݽ?����c��8�z���ij�lh�bp(��צq�� Q�-����k�ϔ�*n���]
�g�+C[Ȃ��Q<�Ɏ�Ab����{zI%��g+�&�R�9���0n[�Dm��ct����~�"n�kv�adx7?3^���	"){AuM�R�9i����b��Cє�o�H��;Ū!����&v,:�B���iY�e���fb�ԋ�d�1�W�aN�N�&�"@��-D�N�W.ꢀ�d��Pf��úW��=���)�aU��VmhB��ݒŁ�1�m�I����/˜$;�����mH&b�ه`wzp���u�E(�{�M<��a����N��X���\M��8r4e�9	�W��!y��
a����2�2�<��bs�ŝ5�3S;�0f% k&BH�L�n�q�3�RG&����I��h�!��Tk�2�Ad8r7�Y�Y4t��/T���$�&��@x,�Q�I�wQ�����Ғ(�W�ڹ��Ț�H�4��X����2�J�j��&!���p�E��X,f�V�nE�O��f��0�$Si���Z�ÔwY��n�y(#/+��	���2h�}�F��(�P��,g9N��Q����2h$-/��un�sl3~y�?����/�UK�rz���|��;:��(m�`����\=�1�\nG�R+���f�����%Xz�`(�D&f��d>�>C,cѼ��╵�s-xaw�{�Q�g�"M	��
U3���ƭ��z�)�[�D[� ~��F��.���w�T�M�ݢ"�Fɬ���p6���Z�~ϳ��n>y�P�~9�2�P��[�N|��9��3�3hnM���8�;���J�`I5���ӿ�W�e�"���z����$�Iѧ�^P]�6kg�
̂�m��3S�$��H�;�,oQ�u������x�;	ܤڕ�Tf��b��[$����l�<�Ċ�N�x?�s���c�]�k# �U�7S��!�!��!�;�V�*>i�/��S}>�� ��i��a���M��'�N%�9�z��r\��
��_؞V�_�#k��S�:�Ү�_i�#P�b����
�vɑG�q7|6�5�X4dG���5��]a���.�7�f�}�|\� #���!�|b�;��N6�	�9�6��#D�膖B"���:�S.[<_z�O�j�q/�u_	�tM�y��?Zs�0.��#Mꭑ@ڪX�����l:*}	�(��ņ��RҧҤ,�۲�(�QĲ��gR����j�c��	p ��]A��O�^~�	�waִ��z�S7�d�k��5�k�6h����GoăX���ɴ#�W춒�����P�,���ayc���-�X^h�wK���V�#MÒ�O��{��
;(��H�d/*�g���@[�6�~K���^�MT�ff |�&ww��jG�[���ҖB�G�v�)_�+��~���F�����d c+Üy��|���Ȣl��`��6��mw�w��Q;[�ʹ�c%��6W��$�`�ŢҲr��� ���e���ҟD�}p7��Y@�+h�c,:E3~	I_[��-(�ՙ�[?5�d��/� �CZ�|i�466aO㠔[|nx�X\�����mYP��~��8� �޽{%WX&',����FHY��	�=.�-��$`VRV��@�T��&�dB[*k�_��=8؇��Q���Dmľ�m��_����پ���~R(D�8�"i���I���v<�����w���le�tZ�
K3닳jO���r�f��&�������16%�boc}�Q����KʏG���s�0�	NG���� ~��a���J���i�-�㴚V�g�:[���y�6�����M+uJ3�F2t�{C�;�ӫ�M�k "41�7��2���ő�6@�u�kw�����	��lTI��ǫN>�I3�8�TR\5\l�^�֎
�I���tm�R.�r1�h�XTl%��{�3Es[B~v(Î�QSF����.����]AA����F��x<2'F���A42J�N���B�g����7�m�(pG��i�l�a�'0��K����]� IVK�8dՎ�������a���V?#��Gg/>�,�c�����R��{m�~ֵX�a:[�̨�Z�sW���ë��w��5��i��Z,�,� �z2bt�`0��j���(9�ʁ�.ڟ`�����8��<I�Rr�\o�l!���K[\�F��A�dB��׫�����|���(G!¶��	�j��v� ͢�iC'�\�J:�&�'�$��M��
I���F����@� R�I��c�#�{ISa��b��i�^X5Քy�\Ɋ ǙKPT}� ��ЊgV�)L�pqZ�]�-�n�ő�b���B,9�l�2v̚A�|�Լ�a��hDҗ��-ϗ.��g�p��_���w���u:��1R ;�"lx8hviU2"S�gd���i�k�.��3��`L����d��,ĲU$$��s��}��碉4�h�4�T�6�1�Y	L=�g%!�0$/i0�EA:
+ɥ�ᖂ�">�=�kt�ϳb {J��sWa�EAؾ�O>O�BD�["�D8ԏ��L�_���"b�j8S�'��&���/���@bĊW^&1������%:H��K@���F�L#E?m��Ӊw�5΢���j}�GH]v#�gf C�+�Q(��'��uH[�<�N3t���C�'��lQ!�E,+����є�f��;�0�9M���g÷-��Cm��X,�o��E<�v��ijG��~	O>D�P^������x�oh'�0Hr����]��ҶE�S,䭻�k�#�ٻ%��Z�vJ#���J�ג����l}�|~Y�iL+s�ל���wcA�wرߋ�o��t?z��
�q�i|�j4g�E��o�m@�(;C�������y>*,���э��aώ��q��45Z;�r�������q���y�>	�~��b��ҳ0`̆����Yy�ho�����������e�.�������L�	�#h��*��r7,K�!�E��>q�f|�ţ3�9�lu�B#�"$*�BwT#3�G��J��i�&���|[Sv���1cV3�o��>�RZ5����h������l�v[�H^qya
\��;�I���-���]��ۂHe��-��ig���g=
�N�X�PW4�l�	�����D1��g��(P 'Q��� ��PL$�h�>��'3%�.�¯��o7m,���U`�:/8��9�ֵ��м�0��$�|7���$����a�VA'��O��CE�&��B�����Q�!<��Khli�{�x����_�m����W����a�#h9zT���2�w�Rt�{��|F��@a���:I�nϊu�jw����{�I���B�t�xf���'�ɂ������"Y��lI9=m��Vm8��v4���6q����H�D��|���8�	��G�eV��U�����a8��@[XΙbmj�̮�A�م����j���*�l�E��M7�@}Vy!f�4��)#���#9���W�3�u�D㐃X�
���Ob�=Y�N���Dǉ����LI6���{9��&��=2�D��F��B�(b���'�8� �r��A�J�\�w@;���L�|χW��&S�ʊ�c��w������w��B����x��f�;T�f���<����"'��v�q��-�
�n��!{�c 7�vD<�LM�P���|Ø�m�aȇo�G:��|�ty�m���ۡ#���p뷇p��\5v|^�⎕�I�ԩ:I8I�������X{�Ͻ����dRu���U��΀,���e%��Lv؉���f�I���`�۵��L-W��)Q������$.�9cVb�ٴxi9�û���JL���j~��.Y-�1���hc���)'��>+�?�n�j2>�֜�T7����n�7��^-�5េM�C�_�0DfCb��e͑���􌟽��S���	�1DF�f�IW���#](-��$��aÉc��C�e�������Sݨ������ʊ�Y�u{����C6��rb9�+ֿ��;E3��5�	t3�C�Z��Ę��P�I{�5����5�������Ѱf�J3hn��Pn�V᪭z��T�W��0H�BjE%�K1��	GVh�u��_<Հ������a����P�X|i��W.c�j����,R�p�=��ްhP�DBt���a�6�Ql{O�������)�?4J���E���㔯��[�|�_��a��.7��
nA�,���
�
G�d��I���Eq��E���d�F���Y�s	��4M�����&�#6���|r�`llX2hTf�u<4��&H�&%G�$	.q��U�o��?nȩL��L��a��"C��Li����*I�dm�e;A,h�q�s�e��J#x�����G&ڋ�]O�ȕ�o7d��ս���g�v��ض�(>"Ϛ5s�>sZm�<X�H��hw����gc��,�ߘ�O5��g��Z��5��]GQS��O�����7�^��Y=?�6�7gq�M�����H��{�()���O�H��փ���G�p��4����>ڈ+ϫė��E׈��U#B#�4��d�Hj�P�}<[S:{'�b�X
� -K*��e��͝Ҧ����x�E�R��ʬ0OI����-*��E��fb�Σ)�>�	;��L:��l_����.�@���Gbp?�Z���aE��4!���QP>�vA���f���3QW��t��<0f!��tZ	QC`��e.Ӌi���"�Oj#����#j�Ei�z�m!�,�!�_���z|*6$K.A��v��y�0�ܓp�BE�FX�aF���%(��5��O��� .Ҽ��F�{EYx]�j�,�%YI�S��i��������*�ʕʜ!��*�ȯ���bFy��3��d����H�	i���6!�-W�G�����R������k{:��fhdm~�v"¾F��d�`�έ"T^p�vB�lYR�lu���z�J�[�fB���b-����G���J�{�Ӆ}��ؘC� b[�(v�vIG&��p���׈H� kQOl$�������G����)@���i<��������w<�m�XZ<�L�m��c�9��E̬՘^�L�֎�3�g��ԅ��Q:�g�	e����VǱF^QQ ���Z�c���'����!���L��&���K�q�B��n��AɁ��+���/�r���[W�1�҇��]h��c��W;�ok���s���V��dMckB��c-5��S9�_C�@�ǉ��硿yH�+�oϭ�ޮTQ���1�lv7Kl�K�s���v���Ke�:$�=vɮ�,+�B�|l��L��Y�p!"�Ei`���i��Է�/�!�g!�!��,Ē�?�G7õm��kΜ����1v�|�a��	��ydhy?C��9��f>���\e���|�5���NG8�BK%��T�02d.@��*"�W\��_u�'55%��PO�>��[�Ŧ��rȖlD�����J��v��GI����(l5)R�d`Ű�9�S
bȱ��#�%��3F�E�H���1-����	�o����O�5>�l�B�	!����ϖCd�ψ��sD x��dM�Q}x��bV6ne����1L�t2%G��!�#��Ȳ'!B���r�)NSc˅t�Y�Y`d����҂�s��LB�R{;uD���mz��}��YK���̮��|l|�/�s�v��E��.8c�'a��f<���d'�A�ʕpLI>���M�H�/C���%��&��A��E�qh����[E����y��.����f�^@�������Å�,Bs�@�ꝲ���:��ѵ������ܹ�b==h�jy��1кz���Z�p�"j��<I��#��Ř�[�`ddX�S[3
G�=�b$�u�}����GWs�}�fs�R��
w����s��>���S�?�B8�k�6���Nl�a���N���U��Pg�.�Nd�����ɒvQa�;Q�`]
��0c��i�i����5+��b�̘Qkn���s'�{�g��QS�3�g�:?���QRR�;��/���V2py�^�,�o{��l�����?2p;����H�����e��g�!�a��p?}�v���~lm����U��	K���!�G^m���b���-�������R���8፻	�"�D7%7Ęc@ñ�LVSѿqeP ����ƍ�S�a�Ia�
ʶ�����#�ZR�UG�XHn��>+�/�<���Wږ��^���#�'����nϥòӟ�N�����௨/�2����ۿ����9�N�Y����I�;������+O�enKJ��c����D9�z��옼�߸q�,�����=��#�]�9��^^=;��ɾ�2,9�Z<�i;��x̙}
���t�����+�d:׈5�<"TC�ʱ�c0Bʿ��͛B���RY_Ngu�ͤE=K^S�Rw>��)Т��G�~����� �]f���.{Jb�Y�C/��JiU>!Q	m�Ӝ��=>��/8��[�Nh��ٌl��3l��Ud�魀�͙�Ţ���Ű{*@_��Y�m�w	�)����X
�R8��)�� �㼽r�UQ;�W�S"j�+Rxmw{>����9XX¦�
ԏ����B(q��ĺ6<�9.�|<�U1�)8rh��4�Kf�ф�:r�f��j���;RV�YM����Ⱦ/R@������zD���sha�����w���Lue�*���%��(u�a����D��V��X�������?Y����������o���&���W̳aD��
��̛0�����"�]�xnY�6_��3g�>`���>[M��E{����8���<6��M�>�|!��{�"GS��#����Z��`z�>$�8�|�\�:e�vCN�Kj��t������CI<�kr�ܸaH�tɩ>�:+ ��_T|���g>�Ww�ƃ(f�@ j���摶�G�/G*T1�i.��Kq�d$��dȟ5��X%m����O�}[�n>|���V˱�?�G*���aQ]�I����s7���>�tdt� �.+�/6���Y'�_�/d��Lc�a���Iv�l�1�W�F��cw��M�M1�'OA!j��䬪d|LȝS���Ǧ�W�#�����cA��?k�gș�*,�R`�ESwO�����
&�!�,�5Nv�{�HBG	n/	����@Ζ�4�|lށ; �4d�����Z�I�J:�Ə�YD��-��n-�uv�A'�Y�eI���b�Y�a�5��lif���Z:���ӿ�ȵ\RAq�Z��*Ǌ���Ϩ��]�i�f
�5�圽R�����w�孭H�#R_2�Lr��w�E�cJ�)穣�1�r�0���Ĝ�/G����\�����sd��Ɏ_��4�m*����O�s^�Ӊ�GŇt��[e�������>έ�Φ6�:$�i�����(��vV�?,C���9X����bH�Hx�<�$�4Ē� �{�Y�.�f[%��&,)��g.4���E�А���(�^��l>%?L�;�Ϛ�Ζ1��P/��H�M-N��b�r��\T�P^�҄����@fT���x]9C�c7��s|-��r<+?�vѻ�S#��mŖ�q��d�,]���ͯ���z�XV��7��Z��Ԗ����QI.7w���-u�G�A_�&2��X8���踠ڋD��M3C��Y(�-˞�ךB��c�u��14�R�)!K�F�:ɦ���	r`&!�����J�Ԝd�$�̶�Ī��H;��Vi6�	$S�P�w�R�s��#:G.�.���5�u�%k�&�fm���&w�f�����qY% %��գq����r��	�Y[o؁_o��g�����δ=�[�2]GVa�rl^���qi�o��7&�t|7����.�]�2����u���~��mGr�--�BIK#�18���`	R��n�.Ʃ�
q��;�tH��<����F�6TF�o�İ�=�X=��d(CM��M��U4�|V7kNU�i�
3x��@�e�王�X�����JȘ���3N�6r�D�������5e���{{E�e������VT&#��d�΄ٷ��^S-u�1~l�=�N�,�!�c�е�����C�[��C	<��G��M�T
߻�i?%!���?��]��Պ���D�w>�
�K}�F��r�Ʌo��!����(	��L����p̼
{�>�{�܄�5g�{%�G��ӻAm����%�����㿓L��[g��8��E���z\{�4�s�/������O� ��X��ظ�_��4��^��C[p���ߝS�ˮ�
#1w��H$�f���	!�׼�qg������C k��1�JJO�&	ކd��պf8\�`��n��.��C�x�w���Ŋ'׷IcJ�p�r֌r�z}j��\�Ko��у/��i�c��r��X$)���NE��Z�)� m81)�	�ٯ����s��
'F<>��dA\�(�Ɩ��a���DM�=m��x0�5>��C;X�g�,vI�$��	�ӉW�ɀ��=���#ƣnz�_)�Ev���]����PKN�2]��h��l� ����a*#�H�#e`,�Q�}i�}Yu�(-&eԒ����
1g�\�*\޽��W��^h&�BkN��-tcFM9�e7��{������TZ_�	M�j��fel�Z�l��Zv��r\�b(�b2���rٳ!ն��YD�,��`H³R���	K	��8.��c(��)��`��K��&fI�7�*��mZ�+L�*��,A
��PѤy�������^��V�H�>�te��j�f{Z�	R8�����0_?���38�B�*$J�Fl>m��J�`�u��J_�I��R޷�~<��;U���p5S[U��\
�|� ]ZZ��$z�S����;g�/���Σqbe1,�[-��P�
���g��a����HI���9ce��<��e����g��7��x��KG1�ՁM��t_�3�wֶ����ʵ"L�3���JWbeiV`�}ؽ)#�8�X2��E��==wy� �$�p23�z4=Β|d� *g�H�E�
�u��Ӎm%�	2Ҵ�rb_����g��l����E3� �E�u"���3v��Y�t�z���`l4$^�$��;+H���q�W�&@�O�����������*ƒ�8�[_����?]0�vE-���O��ɉf�h�C��"�ip����w��GF�������[���M�Չ�� QE;�"X�o#��ܨ�q�tFːU����q��E�~�vH���197��9)|�q����uP����ӤW2 9W�Tt>Ѵw4��!aR{w��Ⅎ�'���߶�p�]���M�S�t�z�ܯK��Ɇa���l�
p�Y{pe��ق�^i�UK"�L�I;a�!��،${�2[Hs��b�2��ݯ!�R#9&��H#\.b�](�O���CmR��u^kϬk��}��#���ӷ�e��XX�������Ӄx4�5�u;�b�A���3�RE3��m9d9�]U�u�������7|qQ���	[v�$���%���Y|��X<����~tE)zmU�og�ZdW�e]{���<-xn������`bL�L^`Ðs��t�Y���z�=��S�����R{9ax��f�$�`C�'ũ���9]�������������ƆVRѳ���~L�G�!a�Ӟ�/�Y=�Zc�A�.�T)ɰ��)��	�l��XZ�Ѕ�9~*�AS���'��2Z&w0����.(�%g�PI��g�e��+\�D�3Ϊp�.1��mz�XF:I�\i�$�xz�Kϛ����f��(�ݟ����K���2�}��-f��z��QE(�D�s�l6�dj2ٙ�&S�yd9ʕa#Q��I$�V��N���}x\g��{��hF�^,ɲ-����$N����%�&,�6��r/�,��@��@�&\��e����8�d�8���Ȳ%Y}�F�H������������4�ٟ'X͜9�/_}��sʚ�[ˊ�h��m��Un!�k�{8O�ZfU�a�F��,�;��bY���x��p0̩R�Lt�8f␰L�#b�֚�KE��܊��ab����JXZk/���z�����zޟ5p�G�#8>�H{�S֡��7��݇P�/6� �Ɔ��س��ĊM͉����Iѹ�N�+�d�U���P'�� �;���fF��V�;� ����~��r%�C1����?*��	����^��H)V�X�}�_������l�!�'��$�k���r�����<r�8?m��Y;q�J��_9߱Sؔ���aV5f�T���3�(O�ʘ�E�E�3�B�[�bA5f�*���0ڻa$X���4�P�18��Z���)���1�"���if�S��Ȍ$p�����y��R���q����O�=�q,�s*���K8�-d��'�8����z*�+p�L��m��8V-�q��$���w��܈O(�I�F�u��8����+���1B�R�pff���j/rYh)h�h�|���-���Ӛ�����>����:TUU��y&�òף�3�����l�i�R��L�H��~tm��y��ee>w�%�Gz�͎_</NWr�W�Bʣ/�W��o��j�l	�h�.�ք=�.vS
s����*Ä���}͚��˄3)NӲ�y��|���0w�|~�h2�[MMƂ�w���k��
W���17���I0��N>�
���"3�&�ĭcT8���|N|:TI{��)V�t}��ʊ���G"�ܔ�9��a]Q�6;ơ�U�L3��B=Z�iN�����IdQ���٥��c^�/��o���uۿ=q�`�<u��[�xPY�m�W�5�x��:~���`�*��.v
k��_��{7Z�0�� p����Oi4���a�e$�T��nY�C�O8g���Ƒ?�i���P]]+�l*�A%�ȩ�ض�ذv��
�L�9��4�������jǏw��05r�D9����P[� m�7�:|������g2�,�d�tTVLQ�09�dƒ�+E�*�yo"�cZ�ys�`G[R�R��
�)\�4ɕ��$c�yQ�)-�\���N�������t�S�l~�.C��YXF���UQ���>�z�c�Ů0��H��3B�"ȷIGeۼ耘oc�Ek^�<;����Xa�:�[b}��a�HT����I�.Kk�ıaI<�[��*�~/�=#�A�˼�E�R�9�E����m>��0���I�s}�ŃTUU��W�$2�"7��n~j���i���72�	��B��.(��"�|ٿ�]�H�~�?��ra�\
�������ʋz��1�t��	�ɦ��l�;5�!���=N&mhk=��1!��u���75��ߜ}��)�ѥ�4���]�FQ��LB3��YZ�ŋ/B�n(�|\=��S�<��Y2�%^k� �?����%J81���պ}�8�$&�-.F�����78�/�ҍ�l��ܶ㵳V���:�3�-�Q*�L���GXICҩ��%����
���z��{�E�rZcT��~}R^�16���2��z;�.;��z���=�����یU���r�\��:�U�\X��^r&�1(�rX�ꯍ"<1�p8�5���؁Gwuq�.�
ˤ�0w��5���/N��٦�,5�b���q�c#�SEI��6CI��g�C��� ��V	בȋ�x�*.g>��}�Eaľ&��l&`c���[{�CL�dG�^:�R�%3�^�5a��}��w ��P�0�/w��5�ch`�_Ǥ�ϴ2�ճSV6	>�IX��q�7�֎~Fg6�[�d�bĉ{��n��N*"O��<u9��i�Q$�2E��-��GB:/;�˹�`X�t@*���y�Fa*u�E�fQ��|>�B��,ia���w�<�\ߨR��R��'a�6azfK�(�h�����*6��mG,2����d��S��!b������#�(�xaslr.;=_�����q��,���s�'�3N���a�%ۀ�_���� ʺ8sQ�znn���,u$ň�)�� ���Ƈ�X�[7e�wD�JG�{��p(7����h�����/��v3�	yѥ�c���xgA�]��U�R�s:����kS�5��j����yi���k�݈�k7#.�ב��b���(��E��sX�x	�r���.z8�C׵��L� @2u;�|�"@�]F�9Z`u�MÛ�m�NM����&|�r��li���}O�0hڂ� Y�jI�s��Eױ������*��G#���cc#p����������I��^?ЂJ�^�������&*L�K��ð���J8R�nX;��zFF���dͺK�+.A{�)��1�
�����No�/ʻZ�C��p�t7�cz��ٜp
�3���E�5�\�:�R���- �̪�΍[L-	`^� ��{~;-c(e�6ͷ��j.�E���)�����rm����|1�*�ۅT��-�3���HʑR�:�Hn4��R�ȏe
�q%"%�hr�-�l�(]��/1F$؊Z���c�Eذ�
�x��\�Τ������H���T�;��]�|-*��~��{a?��2��E�ٲ���Ţ�@��i򈹝ˢ�ʧ����_dۼ�C�ʶQ[7=6$k�&����$JOw;�Y;�--�-&$�I�HC33CV�ݭ����-9[��tp���i_�
��ϕ'�T�a&;�{�M�G��Z܄���F }N|�;�B]C|&�V=�u��cl4(C���(� i��8�pM��#��dB"d�E�t|I���50����R*��'�l��Nf��͜�PF#��΁�驌�@�
;�����ؔ�4W)Ƈ���]��Q.j�.��F
��������K|B�Y]\l������G4��d�Y��^�<�c������|�x ��|���Π�e�^�9O=�"��Y�_H%��\�.�����b�wow*�f��O�88z������X����5��F��E�C��-�����4�H0ߋ\Ĕ2.\��6RJ!Nt΅�vb��+�����%B�u��Wc�G'�8��C� ��V\�܃2�)��-���}�X%w-ա�5���o���o�������"[~����������s7|S��p�Ow�7��Gn�;�:�;nǈ�ުR{��`z�jH�a(uE��I�Úb�a�5��a��H+��'�B�C*#eEwg:�	�gs?�ʮ�8�!#�6%�\�:���
ң�.���I�6���5�N��q|�=�jU	�� ��%q�t�Y��GA�P6ǂ�x�%��%�Y�X"�5�Ģ]984��0-ɟ ϖ�AC��w�_�K����]L��"���q#�Z#���Dw?tMէ��?p��a�����*+I#���i;��A��LB��c���fd��w'�{����k�"Nƙ�Wd5�3��������oyC��r�,��GF���Q�ᥙ� S�`4�d�fFrd�x�]�X�n��aO�|��]HQ��o9�=ݽf4u44�g�>��(�N���/=/�r�M�����N�$9bu�T��1P�2�e<��Kߢ~�8�#�6���d�6&�'
z��P���C"�)[M�Cʲ������j,�8UMM0U�=SbV�[�E���M�2ŐUYTm�5�,�Ɗ�����U�-�R�`���á2xz�m���$��V5s��$����ڈ����lm��Q��H����3dz��5t�JiR���0p��ԥ�p�S�{�a�`���i6#��Mu��P���B`$�����)s�ΰ�m�,CmE1��$�t�C|-:��.�j2��M�m���Y��d	@��錌��'�n��z��9O]�iJ�鮯-�.m�Ó�O�6�o^�	�؊�W�.�'6dX��-�]�G����xfO ׭�Fƙ�d[
�G�SZkG�'���,�	�@�6!w+��N�o4�}�l�{�z&�l@Wի��z�=f&��p��n�a�=�=;���1���j4�8nƱ�G���A�w����t״`-V�\�˼ϣ�Dv��c[Kq��'������a��Rϯ���p�c�ض҇�l�D�V�Ӄ.���dȑP�f9��0O�!9Zlu�߸YK=�8�_�;������Bܳ[V������3��U˿#��G�y�(�|��9:i�`�ˡ!4��O�x򨱊C,��N�	��V�'΍�Hs�e7�Q�H,0at���5��R�P"��E$��زQn�"�m�=E([��t>z��~�dkʰ�(���&��J�jlI�h͊��Ju�9؇�PtYY97�]
����I���'�	P?*��Oq����*����ks�\�Y$2��N�ikA$��PV�<:'I���Ӵ���j��+4x�(��������$��M�@�ԩ/o��]>����5ވ%5�o��'���e�(�'0�sq�]c����a��$,^���l�`�G��8N��`�����՛�L���7q����vd_D���_�E^_������w��I��q{C���F:A�B�7�(BF���ɠ��OLF'�b�K�!B���u|���x(:��P$��K����?�^f �
)���q�_y�XJ���»:��k����Eؑ6��B�p�L���S�d+.���]:��k�ks������6o挡��Q!C'z��Ӱ�@�hL�ͣcGy���G�����������S��r36���]'���;q�ƭx���={��\Ͻ�-h�ph�(��Vš6U\O'�-��J�D_4Ð}�-Ŗ�X|hZ����m��Ӡ��q��i�y��9sg�[�)nÞc�##AY� �'��0��8R�rn��Ԯ�?S�����	��[����+墝^��z��!������=�c�yy`�0�L_0�t�Z�,��bn�!0nU޴�B��KG��cM9����P�}�Q��*����bh(�cp�V�{POZRz��[q�e�,"5<< �V�dŊ5(+)f?ŏ�.�����3��aT�dXõ$ɏ1��6N�#���Ӱ�	�LhyE�2f%cHB��<簊]*af�EפLf:����-`���������:����&@�ڨ�ت�s����4�����*�-�-؝E���G/��|m�H�҄}�W�x��m'q�l�6otb_���N
&Ü��9�=�SS8���Sr%��8���s�`�ڍ�|�x���������-�m����Z8���9���Dč����N���kGm�ɒ�B�gQ'N�~�x"��*q���E��T�ēIU^įH��!������ΟS��Ye,�܉q�q$����Q!�:z31�>ىe��,��h�[b�����`�>7y�1~���Ӹv��h���g��Mcߩa����,4�lG-�Sb#�K{B�;��n롋�����q���+N��@`p.�>G-��2�������kp���2#G�8��A41VZQ��;��_��Z��h�@�����6���:-��<�Gd�e.�,�w�RnS�>�v2�O_�ǒ�L�}�\G�EٲbJ�T��-\���{��x�9��=|K�U`��DB(����'��&��ۮF4m�P�az�jp�U�0�#�}
ϼzq*�'pV����L�o/A8��8q�h�d37~��}�jn5��lj
W%�.i�"K�u�	X�i�3�����}]�v��I6;=���r"�&��(��~c�p8��O'9�_g�����4UUK�uT�$�Q�G!)u��X�ƒ�U�NM���؃�#�
e[���	��i�Ӯ�3t8w����t-
%�u��V��7�]h'�m=���bg&���6�ͽ	l:�3N8�I���7�dۯ�*�f���Z��k�p��7.c>b��2��O���/_�Hp��碼�cH���	6�/���c���1n�h��>_)��c`��۟m�!��+qQe��|���ʥ;��R��8�x�F'�)�śʱh]~��(�(vJ(œ{����b��d$���)e�6!��g�'�u�b�O&q�������c���na�C�Fx1�yu��1�O8]�t��O/-DQ�W���;�!;v
�Va�u�9J���[���ҹL�eI�Ž�ص_:���1���A�t""y�4G�Ev��.GF��:9�,qs��@�z��܊���zh������C]q�8���G6ظ��l��y�)&^��(�ǰJx�C���[ދyV�{�:̩o�Ҋc�Ji��e[%�#���HG�H[��Ɏ��̢%&�Z�K��ek�����d�lhr���K�s��k8p�]��8��/ݗך���mrf3p�X���Iy�)�A�|_?z����:q�ex�MX��Ȯ�QhɏE�A2�R�!"��V�ё�+�Qs�2B�5�������"���{nX���-n��% �D��+�����\���4�|�$�F�۾�PT���٬RQ�397�2�
;*L����(K,�qd���*	�۫�	�#M��Խ�R�B\�����ոfn/jJ[��ؑ��fe��UE�Ŗ�$'q���r+&k�H��9jaD�l>��;5&x(�A	0����fi2�c���� �q!��IZУ�sA����b�����cx��Zܲ��ʿNw#ֈ��⸎���y�N��T)&C8T�*�^[�u5ˏ��1(`LX/�٣���t������=�Yev�ۅ.i+�A`ҍ��r�c�Bs��a���R��{p��,��N�VJ��"G����i��t�xy��$6[Ob2�e_�@պ�Vv�Ʃ��_��O2��Z3��V�	a���P;���M���5b�8q��hk?'.cg���&M��n�m�ynC��4�:-���/ Zc�?�)AHH���I��A���e�d�f��]/_�� T6�[�yAs�1bA*t��a���#;�܁�j��a����{H�{q��(=�L�!H~:�T=��n?*K�4U!$DF��=�ߢ�6+\�YUs��v���uV��W��Ql1���!+N�حH�#X�����uJo؇��<��0K�a}��H���V]���Im�mu�2zF򉮩������O�h���O,��dr��P�YE5��>�a�[���+�X|R�ۤ)�H�u�IN�6t Z�\ �g,��;���v��c�KpC�..=n�Oそa�q������I4A:j�S�"����M���mGs�S%m2	ꈖf�[Fj��BMQG�	D�C)�hKqu�$�=N�����э�?�Qު�vx_����t-��^2v��-E<}��Ǆ���̱t5�+b�S���� �x/wߏ���d���	)������������]��b�c�Ƕ�4~�BHlи�1WQLf:�=���S{*P,,�3�7��ȝ#��]S��5 w��̚��M�<��#����n�]E�q�����P��w|b!�Յyq���_6�2<c��b�02:O,�b��ā(B��Q6?��娨nT!�bT��
t��bsQ[p�&8<%�����K�BX^b�Fb.nS���1&�[W�>3V��Ȩ�&�p����6�P��tO��W�������	�jW���̛�/�<Sb�0s�2�-ӡL���
-�W��D�E�o~1)�{'��	u��"�_���$���g����^�����(��Fq��I/B��xK��}.'2T�<��ܖ&�&����=��<����CI�Q�qi��b	����8�?��`�V���R�Ԗ��:���I�����I��}o ����D�C	�4p��!oH޼D0:@���V�����{B�L˾T��H�T�`�����wGbB6�u'�iS�; �;�)��@:#�i]6r4�U���L�$M�h<Q��2�,�.6+Ĉe�b�̉��]ރ����ҵP�I��0j��td4�O�T�3PS�'����y{}ոtQ���>��k�ps̙����2!�6#w
e�RdΉ�2]��p�X�e�pdbbi;��1������K�7����g]��]��Tr��?Ȩ�tG��Q_7�Is�=���t���Hm(!N{MM�����kuuN��y��H[�(�:0�s�N֍ٴ�$��ڸ��<b)��!�EsX�����X�H#.��+���+�Fu�m��!L��#x������,ә�.0Ʒ�ƑS�P@���7��0��+g1Й���� ���Z�ӹ�8y���p#\-���oYd�Z��t)S	T�Wa��&>��}=X/�o��C��g������pFS'�D-�E�Q(
̯k#sK����ېp΁u�4�^Coh�\OL�u�-QF� ɬ�Pκ�oN�l�9T>OF衣C��ؘ�R�M�ǉ�����aP߀_؁c��D��V\��׮;c���eΩ�3�����+6me��q����(^�~�V��Wo�Ex������3��kK���L=��Ő�:5�!�_:��$Sq�^������{��_�k����o;#�Hy��ƪ�8��
�h ��<��d�x
^a�nذ��}��� �#	�P�M�Q*,�ɤ��&�@
���6�nŜ;\��9���XD��3 ��|�<�6�#�����k���=��;���i�`)Y$/U�U��9^%�ϧ�u�z4�2�89V6Zt˞��<+%���\/���M���P�XȚ	'��v��`w;O��E�N�p1̪��勄xKx��>�0�3L��_��S�_�8�ekː����-�2&�o@~����e�ԗ有߫�/c���ܢ�.@�R��{�)�|Kq��ۅ�jU�QW�����L�)v��qH�:��~N�u�t=����dQ��iJ]Y��5��@b����gd��3�C��ɑiL�̐mY%�L�bd�$0���hPWO~HMҺ��8pf��O802)�]|��0v�>M�)z���ɉ�������*+�u��p��dݓߥq�����v�����y��e0���Q�D���/#��Χ ���$u�ş�u�Iڤ�u��.�2��p�,8Щ��75�����R����m<�L�eW��A�k�b���=D���t�Y�(��$�gh24]���i��S�I�گ\޼�R�M
���a^%F����$~�#̧��E�eE��En��w5���1U��)x���}D7Qv��AOZ\����{l��X�������v�l�DG曽2i��Orr�oO�w��r�ap$�d4�� �D��yQ_�G(g�~�P/�8�K	�haŋ�#&�Ѥ��a���Z���l��b��^d��I!����Ǖ�-|'�N��o��C�I�����}-B���W1��9�X�'���c���[(����aȲ̩��}���p>��0x����B	��.���
�xS�$����X�v���˭�h���LX7��Ug��oZ��W����;����uڤ���L�ʩ�׏���x�����Q�+���{��*U��hp!#��tЂ�i��8�9)Y�I!�8��xTN S;չ��zMvd�i1 �pZ<j* _���� 4�7|��m��ɨ ��z�ײ�
6
�w����-���9-e���,4ɑ���'8�F�)�sf���kۺ��[W��^;O���ƥH�a�=l�t�8!f�r�L���R3��\���5�~��)G�V�܊�i���;�nI4�:C,��(B�Qx��'���kҳv�<b1,���h�Rp�l\�ә��r�(ew����"��6���:-9�Z둑a+��'�@t[�)B�S>d";��E��!�;Ig+�����i.t��aNY�p�ΰ
�j�a~��h�S��'�/�nj�$�+�-{Rb��j!H�3�7�5\BL	=�����5�n:�s� ڔ0#��DFX@���i
�XT�o7HBj�N�ۼ���E��1Y�Ou1�C�Mr1��!i�%12:����p���8',���v��3N9eW_}-֬����悈���<�Ki�S��K��MtUYf��V��pϢ��`F`��+Ӷ��~+BC���[WU�뒵%���G�x��0��R+����XR���g5|�"'�>�����S�XY9���/�h�a}����N�b�W�0wO)J�0��:hc�sn320"J�'#YL����́_?�)L�>F�3ə�b*u�KUZ&DPŴ/�4�{	_i:~���T�%�W:0ߩU�MT
�!2tT��df�֛��+�'���Dֆ��l]$6�Í�������F�j?�̋b�J7�J��[0�l�hW~��!�����K��n�w��KQ\\��DvCÜ�;F�B=��s���ĢP���V!�7��� ���oΘ�̔�䋚��<[�L��5wN�.�3t8�{���^%KR���2��Ktt�۞w�-���IǸz�K�4�7�J_�E#��%����DR�=����g��e�V��w?t��E���ɫPRLD+
#$��_.WF��%�	2������/
e��p5�i��-����ie䤛[:��D����H��Lz�"Wz�c���X)�� ���`aS��?���s����e&�p��3�y�*�{W&�ט�ӂi�L�_�&�>ޙt�O���'DZXD��A������Ɔ�[P�/fn��Ǐ�7�l����9�kĲ��i��L�}�d�����@&s8���^�(����ȝ��شi~p�?���"�Me⿆yKp�W��;��'�z���|�����Ƙ2G��x��բ�񧝂w2L�q�}5�u�,F�p�kp�?މ��N>r�a��M��)����ҶT��nu��NN
�����;�y;���n��f�Y��-?�.��'��V=~B��$;'�����fN��5���`�"�);y�E��6�˖�"��Й���1r��v'֬X�>�~�E(//g2K�����z~DcT��[�Λ<8<��d�BL��E�Z�O]Y���~��/K���Sm�P�f�NJ+k�ч����a3��:��q貽Ĝ�W��d���t���|{���a8*����!��)\�a��A��ԁ음X$�d�����S|����)�O5F��_�|��՜HiE�&��ߕk,�L�С#�r��x��?t��1�,vu:��c,��%br ��M�G�Q-��q_@��I*-����8r�]ڨ]�O>����~���~ 	�G��z�?�����Ơ]�x�Gw!�]����aUD2͍?U�;3�Hت�u�&l�c���g�вԑH�r�E�,���{p�����y�>�������c���n^r
q�����X�ְ��%;	"BbE��O�$�$�'��3�h�x�,��,��"$6YƠs��a�����'n�>����ś/���沵3�'�_<��{wsU���奧.cYy����Pa�T�&�� P���{w���kƾ�8�������.��+$��G$���l��m����]TV�X,����`�Kx��l��dbVU}=�סq.��CAlYT���Q~��Z��d�Y
�3H�]�x<�aq��R5/������K��ۍ7O�N��}����6������~:ܟ��f�hÑ�~�^�^L���������&����7�;h���;�O��$6l��?���Rp�f�1��v�A�1C�1Q��_�'��fܰJS*�����Wۗ��EN�o�	��2�����b�H��/��$C�Ch�M�!.�8�Ү'�g	�ԅ>�'�F4��ے���r����z���I�|���}����g�)�iLL�D��.G��>�\T.�r�۾��o�	����S�2� �;.`�|B{�7����ĿS�e*iGCC%�9rr�)[�z9���Z�X�R8�v��1���{���N!�{-+��t4�����O����    IEND�B`�PK
     w�O\���� � /   images/bb2d2ee4-fa83-49b1-89fe-70727f49c778.png�PNG

   IHDR     X   �v�p   	pHYs  �  ��+  ��IDATx���	�%�]�_��|g����]}MwOkFs�f4�,K�R �/����!B��h��X([��e�]�h���2�¬���>�g�g���y�ӿ�?߫zU]=���	j}?�VW�zGf�|/���     @E@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�      �A     �� �     @e@     �2      P     �     T     *�    _w>��O�*�㚣�������t����)�V�f���{���U��m�.�y�ʷ��s�� >�+�A3<s�& x]    ����?~���Co}�_("/I%7�iJZkR��reYeYN'۶u�Ss?���$���L(C���Nׯ_��������a�����χ 7�    _Μ9����L��=�udYan�9TH�>��(8xȏ��V.�"��^�9&��9MMM���������ͥ��[_��w��J pS    �u">�oq�/ٶ���[�����,KI ٺ]B���!l�o|ӎ2?�Lk�Qo��cG�n�������v��́'" �   ��8x���:q����L)�
+������,3� &t���	)B�b�w��k��
�Og)}��q����.<x��g��wC �   �Ҿ��������t`�ȷL���vӑ��3[������%5F
ʋ��R�KP!m��
���T+sm�|����+��@   �������ͷ�9�,�\7Hr�{�q����2&�Z�ov<��1J��\�3cH\���g�{V~. ��    �4�q=�qT�ui��l��Te�(G�9����j2���Dn+H���a��̖EI����l����h�	   ���ۅ�|W,�.��v,Ǵr��W㙮�Y��-�ƍ-�0Rv�*R��´�p��d�H����0V~��� �   nqS�8n^����
'Mb]��l��&����,r3 };<��������5@��^�L�*�8v�{�y�a��&@   ��&�Uq�HGe�os�*��]���,��2|L�1�
Қ�
�,�{�_��'ϵS��3�k�p    pK;w�~�]�/�������}s������JG������aȔ��-���Q�����tْ�1�f�2�'�*
�y����*YG�p�p   �-mss3:����gͦ������{��z����r��� �Ҏ֑Q���Gi%1�W�֑��!�LXj��}����{�����t	 v@   �[���R��ы�_{��j��Cۭ�i� 6vL�+���A;��.�e����Ddt��8j����Ͽ�Ö�I��;D��X @   �V�<z[Q䷿�Mo���{�#�ͥ��F!(����ؾ��(�욖wB�`viQd�x���j;v��>���9s�w��   ����}0����~�]oT���:52L�F�M���k��?�����}l�z�`������T&����6�_��#y������C    ni.\p��>ժ��ZVY��Q�.̴�H&��5@�j��y�6��M
�:~�������ˇ�f?�O��?�����n��}������	��   ����U�Y��E0�2�g{����:fT9߱�LP�� j4�R�����){�L�;y�A%-#�m� hi� EQ���w2ɲ�����<ϓ�8a�@�o�[e*�~����s���V��ޕ$K.gI��'��Y�gf��4M��`�pXJt���� N�d�l��u�{�^���W��'G�����3ٙ3g4�-�    ���i�}������<�^���xu�</�v98(��,��A�e�Τ��=jپRz�U˄>L�Q��,���}~�TF ���\nS�hڬf�i�/]��YNJ�#�o*�E�u�r���s�M�������G��ᐟ�-Dt��;��Tox������-��z|��-.�םnG���666���Y�=�{�Z���<���ֹ��"pܜ�8Β��i�;� !�Y����;ڟ��r�K?����?C   �[�4�[X��Hx����^dyn�GY�k���H�&|�;Z=��}X�1�\B���`tgk�,y=ѕ+/�ָgt?y^_/S��8��K;R��[c����_�^7�9+P��2���JƑ �]�0;��}i�Q�M5��őb�.��
z��X�R=��)Ó\En�RMI��:e�r�$u6;�w����+J��KYZ������
?��q����������������>�D���   �Ҧ�-��*��0{�'����z��Pۃз���a�E�c<��*��ǲ�[;���Ĕ��K��q%��Lh(�b��Ǎ�K���<�'��K��2y}�����b4?����$�p�eL�mK�1��=�s]��3	��}�_;"���y��u���1C�s�\�"�ır�U�Pt`����Y�q$���
m=�8�Yl~>�
<q8��o�ݬ#/k��O}*��'?�|�·}���>���Ŀ�8s�LF�u   neVө�A��WJ�K_���e'#�	
�ٯ���R�gY.����k����H��k�B�!Ǆs�C�c���[j�<涭*mbP�	 �e���!� -/�(��}ը���)I��l]��?���rQEe��`�"$��O]h�[9���2X��2�}F�	�� ��6m�֗Z��e�����T�B�8��@�?����͍���~�W^�z����?
��9iE�P�ܲ@   ��u�̣��F��u������g�Mw6;4����.FA�NR<k��cyew)��*��O��L�<�vy���dˇ���!aD�����h|�u��´t�Ͻ�j��xf/��B�t��k�x�g.��7{r�����9�*�n��J�]�Y�'x�(��:�%�PA�8Hd��s�Q���#��d�Wi�)��U��m�K��ǎ{y��w�ȑ���"
#��zm���/�z�_
�����n|��N	n    p���g�N-_�gZ1��~.j������s��ez��wrq�S<I����I�![�.�j�(�2P�J���k��؎�v�,?�5q��-3�|�XyEu�k���[c$�84R�{�`i����G	^I�(�p�	�\��.����I�����
����r%I��E�&�fx�8|���%L���y]�x�x�� 2(J�Y����j�F�%�׬�վ���S'�Y~����>��+/_�ԯ�_�e�/�����>��O	��!�   �-kaa�h-�� ~:M�Sd�'/_�2}��wQ����JesK{��Q�"��r�G>�'}���j����e\FaO�Oo�ɠ��q,e�]����[�U�-�x���3�Dg�C�ε�⸎�"e��((l��2'�<μ��1�3ӅKm/S�ܞ�k	��"4oW�bb�]�L�����+������-+�SG��hW����'�d4�t���z��'��q��+W�~����^����/��ޏ}�c��J�5	   nY+++��Ç)7�76/ۮ�v��5���ճ,��W�B�������$��˿w+�}u�s�*�r�4��8vȀ�Q�of�*����ǃ�wl��{��zF��̨���y]��3�c�J��V���P;��-��N�`#}�F]�T9F���֣�2SbI�5N6f��2�l�g���P�8����-K�yNsS�']v�*g
�1*d^[��dړ�$�9\:~�)�w�x���O�z�������K�����=�k   ܒ{�1��;���vFE����9���*Kξ�b����I�(����X��!g�q>5�w��P� �q+�Ϋ��.Xzb櫉`1:�]�&���5 }W ��a �fL�����(��Z�1�;f�����O�Q�L<q�x�x�Ʒ���bSv�R�Y�v�.�(�����ɢ��#�B̴�؞�X�rF/%�X���5͓G���˗/���������W�~zjjj`�ڀ    �.D��O?m_�^wZ�Ua�]K���|GK�+�/S��U��3(�tw��BAy�AS�k��e��5!cF
�ͺq�z��m��:�ήWzW�ZSʟe��](�+{���wV٥�<���q�(hG 2�=
�vk��7�ݏ����b�ŧ��=z��L�ՕMo?�dH�GY}f��>����2���	�.��������յ������_]�|��]�xa�o1   ��X�=��:O����=os�JENm���}
j�^�YOοr��6���c'��8XE9���e���a<ƶɖ
=�^��w���32Nv"W�-%Jo/������\k\��A7lK.�s�v��I��)~��;9���T»���[q&�k{=��g&	=����o�V�n�x�uf��k��\Ղ��C�ߚ��C:O?��Y��~�c�����pĿu@   �Va�9sƽ�wx�|�g\�Nf><ϕ�R��&��Z��&Y�������fд<�P���*�R�.���nQ�]����Pn~��o��״~�����T�f"�q��n|n	!��}'_S��Co�Pأ �ZaI�.{nĉ��}��ݳo�u�d��Q)�O�u�l��B�+/�z>kb%�9��8l��"���ܴ�P@y�-�͟V�տ�z�ʏ�o���ߟ��/>�q"� �   ������Aoss����K�����<{z~~a��Oy�(L�:����8t��%%W�:�y�WF/+�����j/	�� ;�!ɘ�bG)���&��J���(��0�vDߚk�`p���}ʰ��q{��� E7���לlA�Tn6����j�d����/r��>�na�s]
������V����9���=~���_��G?����ٟ��{��    |M��p|���f��]iu�=��[ӽ^Ϯ���ѣ�˖m����}���WVt{��s\w��r���1�A}tu�E�0.m�6��
s�� i�O\�p�E@..(3]M�>�k=Ə���s�
��m������A㻞o���轫�?b�nl1y���o|���]޶3���D���"k�:29ձ_�~t��3�c`�]ͺ�Y�w�}�@�IB�z�o1�i��i;��n��������{����/��C   ��2��w|��ZJY~ݪ���y+FӧN�9{�?�l:��`��a��쨛Y�B�EsQ��"�����յ���F����p账��s�p�~��c��W�����K��|7+�'o��b1TnS���/{�nV�Dv���kr	��a���3�<�G�)Rh���-����N�L&
vlR�T{��\���?��v��?q�ȯu:��|�����A   ���Uq��u_9s�T�����}������NǉzéC�v��OY��$�;��]�Bw�򳾲������7k\ާ������:O�<�kIlO�4ǯq� �]�F-[�'ԍ`�dK�덃�3�&�sm��}v=�����h�{ոǕt��qj������5��&�$��1�ϧv��l_�q����L����i��\KŌl)�b����$miO.hR�}Ǜ��|��o���yꩧ~�G~�G~����B���  �O5ZO?�������;o����w����bX�>�����x���֕+W��/�}�s�����1y��˗w<����֥uyي��;D�;^^NK^���S�w��g�� ���?~�<O��3�2]>p��/~�666����Eg�'�'�~�&m�F��vݫ�͇�����<
�}�����T��Od�f�8�$�xx������q����jm��������U����<���]]�N�IZo�[t�<���
Y�V���Ϻ�_����L��w���NTX��ʺw����X��۲Lg�R��pH�x�ӿ��ފI.�>y�Js~�����磊�8�66�$.,���;��"����z/����a���kz�H��xo�ʊ������;�h5�>�P�?�\�w)WA�-�v^��Q:�#t����mp���s������w���聣��K��0W�`���羻��î��Q�-o}k��Ѡ�֢��SZ�J쁓�V��Sϼ�R�ҫ��Y����s��W^͖	���I�!r������H��~��q���A�g��N�TE��y��������T�Ȇ��f:ӜK_x񅢳�Qo[���V�����^n��W6�$��3Y���X����v�����7�=�B��~o�+W�Վ�vt1��c��.9�W����Gi����6Y)�m�z�.�Y���0�/]����'�"H6/�|�ZA�UK�*�Z9��|��=��zSs��N�g疴�]��C�O�EŖ�lu��vD1���P4/;q%�]+z�K�ţ��Z�"�}��[��'���t$9R<M������?8K���?�dh�wu���������5/���b��Rq��[�/,,X��ԧ�gsci���֋�"e�f��cb�q�9ղ��++�N�M��?������i)uڶ�yR� ����]ϲ<����᫿��ems�%ǡN�d�u���;�^1�3�h�б��'?y�V�E�\-���i���r�\��/?��O}��KW�>�R}=����p%����dG>yǗ�k���ܻ�9Yxy��y���B~S��v�g��e��W��^8�&����Q��"�j׎�8�^^�;2�u{�����
|�6L�d�y奡K��u/p�����y�U�7�Wbߡ�k���W.K5on�{*�W6V�����v��-���<�=%��T��˓kM8�����u@�Y��`�qHP{哅�xڭkzL<�L�[켸�\�o�Do?�͞�Y�nv�{ �����{�%��yn�"c[���m_d��Y�&�������q-3��vL,�˒��k�|�>��C?777��������0��1!�|=���;�wokn�Gn;�8��x[/��������^����437��,��z�I�T�e������Ёe���}��5�T��/,��4W�������C����o�S�/Q�� ����6��,/9>x?��.m���{｟�aLA������t,W�%.����H�U��Q��To4ɛ���O��Ѭ+�X��� �_�/���[����/_{Z�ʓZ.�e�.��	}��k�WI���|@�/�wӝ4���s�z~G�>����o��w��� ��n-��A������¢+�Q���~�����}�a9�j^ng�p�c��9��{����dSSm��Ô�Qk�ŹZ]��.(�?�«��g��{4ט*�S^w�d^�Ν����SW9WBS��$�N��$�{Cn�ӝ�\؄�:ml����;�P�.����ﲷ�<�U���x9o���<���Y^kt�_3�N3�8�����>��/���,�
���wr�M���N%���fo�O�g�쑔�����9��YY�f��[ҷP�ޠ��hqn���y�\�l4�U�G5:�����zy���¼�BL�zp�_+���nzS��m溾��'KS��D{\��:���ZMFe���Ա���\�Y;��*�G'�ѧ��F3cL�4�'ȸ��;��VkP���}�ί���p`��	\*��xW/�Tнo<N'��B~�,w�s��RF��k/�����{=����*j����g*��t-+�������g}�n����0�r%�(	U�ׅ��v\G��>���$1����,,�)�Z��^��:��=���^]]��ŕ	:y�33�O�'��t4�N������:�3���z�>�-����ko8@ğ�o�����?���N�̅��0���t���T��5
H]�j�'I�_��<��oR���W��%Y^��x=��r�$�\���:�)ne���%j���V�Ӥ���_@}��AiK�*��G��^������Qo�9[H�s�z���#�:����'�M�(�A4Զˑ�HU���[��=t�{�����yRIj^��(�3���~���՜R��QT�^�VQ4��/Ί�N��N;o<Fo�x_��c^�3.�u��^į������ų���K���M�jd�)oS��ޞ��z=l�y�Ļ���OQ��4�&9�G�s��?�L�h���,J��1�n���2X��Go�u��Pn%:Ҽ�Q�O϶�����kۼ��ޙ��+��4�w񂫜���fo���33'��,I�k���W�bS�8K?�=1�����+��5����g���߹̴%cE�����G��ֳm���e�:��$l?�z���X�=�� �Z��l���F�}��/U��1�nJ>�;�״Ó�h�d�H
�ڮ�+��y��633���{�c����g>�\7�B �u�?��9�8�O��I�E�iߎb*�V׷m�k.t$=>�5mM�*_Z�xHs33d��x��
�d��Un0q�i5�T��g��>J� �(�b��$����&�G�wsJ�Œm��r����w\�ˡS�Q�f">h��R���O9Q�L3Xd�.�l3�����|�W�<QRx�Ŀ���=.��t�����C�\.�s| ����q��T�9��Z�57��h�r'5��DQW�IEy�Z�@�����l
)���upU�ߗ�J�x�w�5���h-pqe{y:�h51��J8$���֚������)�<��b��N��T�A"�"q#�Qw���o��G�ZyQ^�J
��BRث]~��%^��bS_���p�;N���y�,N�H�"Kq0kk98y6o?���]�����8����z��^l�?�@�5�ɟ]~B9.��|䨤rޞR��A�̬�X�/j���H�t���I���q��E��Qſ�@n�1g�$��LZ
��Z�$xd�s,5W]IU�𾣬\i&����]Zuy[�~$d0g���>!aVB/��J�?9_�����6�r�$=Rɵ,_-(��}y[�6;J^KN��m.r3	Z�XI�J�a�;�r$Le͔��C"�vˡ��W��?���.�4Kxq��[��a(*���H�8��x��ޒ�w��3'���ƀ��ʹx���7?���B��>�(RKGqȏ�y?v�$�T�G��8��u͕�K���Q��)>9DI�{Á٣9�������?c��܀$�I�h�|	&���EP�88k~_�}"_(��gV8�xfJV���ty+h���_<�
��y�"���֤
�r	P��o	�r j�gIǼ��3�y�ur�;��q]�.)���l�����?�4/S�8���q\�58��g/�{�d2=t��g��/��|oټ�Z���`�5}��2�hϫ���i�%*��W��Ʀ��\����7Ջ�%z��I�Uo/�?O�k�0,�ƟI4t�w��7�����t^��f�ߣ��r7�{�<�3�����dz_9�t�e7մ5���I��x�:�����Z�&��3n����sꦗ�]��z=iz�<���!�/{�I����GKEyE�� S^��2��SՎ�~�����55��c�jy�٨n�B�{��q����ivo�:ehQ[cm&揟g�b��-�e���������>(.--��j?��������ȗ�R���`ŷ���텙e�ѲW�ޕd�6(	".#.��T&�Ԭs����R�Ka�^���1���lհ\S���B7W]�q���Q�<K��������5g����f�Kr��rm3#��\3u ���/Fgpd؜!;�(�*JB�������>?�5�J�X�_�Z�D9ʅ���p�ů�S���rv[^/~�i₃�ۣ��R��A��5�����Q��!?oA��)�s�w��e-��쌜��F�Yk��.^����r&^�<s�������)�NM���Eo'[�JU阓�-,p���t��#9�ș�F�N/�{��e����Х��M��i��T�9.�aq�ry�sPJb.dl--<�����z��sj}}�lO���,;���}���0���ϫ�s��Фv����6��wԐ�S.Kش�ɟnS�՞�Uݗ:\4R@��Å�k�����
-�_"	a�Q�7PJe9��H~Ox��FS��jNY��5�G�y�$�4-�5=��gZ�����u��j����݌�ש�k��AU��V��އ���9f�y�� �����3.��%f�&�UāEm69{R��dߜ��~J1�/��̴��v��K�ߪњR3S��:�+o/~2�!o�2Xr�|.�%��7�w��˦x�L�"�稛�|���0�)?���\M:���g%Eu���M��z�l�8i��W>��TG�F�lp!^��c�2����M3.��}�pH����f��\�;�o�u%\��N8oi�q�x��q1l�]����?S���N��le�)�d��w�|����TQ[W�r��=ל�$�'L;���=e։�\;M#���\P��j����tʢ(U�Vr�*8X�҂��04ؓ����s�9$�9"����o�w��d?��l��(�$�|Sv���<�
-��|�%�F�28S�`�t6�&8Jr��Ȓ���������iJ�{���m{J���/~���a��� ��\Z���>�J���%|�iyR�煨�� �[~C=x�.�eu�����;�_7�;.�.Ga��W��Wo�.���Y��FK���wx�����[v�h���u�u���&LD���9��R`���l��w�����S��2I��v���
�lW��T�e�}͔�A��Ǯаu�x�a�k�݁d���a0�.�m��|p�����h���+�.��@~���Х�z!��-����ozӑa��߻����k���e�R�z���q�����V����A'����p(_�rn��R�-��\��43?'g��3��Ţ�⺢�r3s����*���C��w�|�J��[�Fn�<s���匩=�r��ǯ̵/e���R.�"5]��Lk4���ș|m�v�!d���s��3�r᪌��C^٥g�	,� �3)�(��ΥЍBS��\P���	�j�)��4q
.^�9�����-�ڵkZ��l���U'�K5��3���r0�o�7��[3���X��qX2g�S^_�4�{�kMgfj���>��-�j4מ���Y%�F���m.��繩Y�+Y��k���H�).���w�+��˸��n�2)�}."��l?'T��R�����׸M���d�t��n����Tfqyۋ��f�A͊��
�ρs=��27�x�*]�2s�b.��V@i����@���Z����8���������{R�R���:́���T�&��)ry�X�Ы�+,%�HJ<��L�jJm� Y�t'���1���۠qA,��\�У�LI �nA����i. #�i���HzA��\�T�Ҫ�x�I���5%;��ύN{����K�$p,��%��G�K�ţ5�=�8M 4��-+3]�����k
����b7#�%�9T�j��!��,�j��T����G?p�e��,�|s�?0��@�x�i��nt��3k�o��;��O�����AZ���%���S$l��)���[����R��\Nڏ���YW�y%]���P�:��S�w�Ukm}�f�W���$?�ٚ�����f�������6A�v��H�H�8�JK��R*��߱��\i�+"����)�r�n2�̉	L��j;�m�W/�.��(���uHB�t���J��:{F�,9�]�V�h�N�1*�Y��k�i9��[:�H��j(����}9(��(ż���!�͈?��/�P<4�L�UG��,�N�����ɡ4������yK����>���兮YJ_�u���}���$���N=/R'ѹ}�7['�ksS����^��f����ѹ����8]�W�m�f�
կ�
 {ؾ�u/���s_�d��W�x�V��^o��^�߫���x�^�e��n]8q����c�&��{v\eW����_�ud<&�7�ˉ�ݬ5�t��w?4j����/�}�w����+W	��A �[�{?��Z�X�s����Er5�8W��Z�[��iJ�PӔ���f��	���$�&��6� �SR����>�w���t��@r���&]>�2�K�i>�jצ$�b�.h��F�,����wL�]��k.�>�����ړ3�rpr�S��m/'˜�Bs��s�7�;�v�����\��ʊ�$}�.:�|0�˖�F�PrV3��U���<�o�
^g�p]�R�n*͏��89)rSWM��<���υ����
Kq��n<P-��Z���ӷ�R��ǨI��x)#9^P�ד���f��3�B�` �ť i�t�wj9�9==C�AWI�kN5�AC��p5�(e����KW/�%�|r���/��~��Ԍ��#g��~�����B�%�quHR$+��;��M
.��`|r�������=�^��^1T6�)o%�$�M�t-�Z5m�ޤ���\>�|?.�e萜�6~�d_��>Q1���&�e9yyRh%���v��,c4��`�������t��,��0��k進0�nd��J�C'隙b�Q�S�rc�?W�\;Z�ѹ�8<H�[p��>/�ŕ��E���n��t#R!'�,�h�ХC���?�Y�P�R�r�=�!=���3�n�G�9	8�(.4�N0=�%�K�l�y���U��p�����ʉ]���t������L���w}�JҐÑ|tR��Z����X���8���f����Z�3�iΡ����I�q�2-	�(�=�D>�$ ��fNp��v(i�HyY$�X�3�2X,�0�%���Mx�U6�����p`J��Ҫǟ��â��q�/�ff9��'�x�ZJ�}��e��N~�����I@��������8�-0i�[)�Z����	�[���d���:s�XBiA�V����I
�����7?��0���˩�>ȗ�a�Ct�%������/ӥ�~�y�q ���N���u�LZT��V�
m)�
Y�4��|���d��?��upp�L"] e���亵I�0�����t�����G\~�&�n�$���u��}�u�s����z��.^�XﾔE�K����Vsm�~1$�k�a����s�CIdƾH��qT��VL�H�r�����;���������T��~���ͺ0�,h�o�����.x�%�vN���,�S
��Ik�ӕ�*7�8 ��'�������L&�wCx�u!���cp}1Z^��9������	�L�?M�������9y�ĝS���xw?��}ꓟ�$���_	�҂���Bk)͓�(O�q,�>����Cn��β�M�+��\���`�[Jk_�!䚹��g
e�v��KO��H�!�zey��琳�\��6�R��NA�����`�V�R�r1���rԗ~߅o΄��p�a˗g&��S��*ǧd�U���˕���y|��򐗹Թ��Ԓ��i̿�).miȿ�I/+ʴ#~ʥ�dd��y5���tI�K��&rF��y�ra�E6!҅���7�fZ�������W.������Ow��5�����_��N��M���^��;U5gܕ��)��}�ՍU9������Ԛv� q)
�5.N|S�ˀ¢5�N�;<:�&�íqO�r,�!��A�\�X�),�iA�I��m٥Mou�0�r��i9�?�4�[uz�up�Z����TD�^hO�z*�"]TL`��r�fgt�+�6��銐�9�pQ�_ݐ����N�p.�_lއ�hh��,�Rˀ{�h����QǱ���ק$N2�����xi��R���`[���@�E1ʄ��2�A��kJ�`^x��b16����@&50֥�Z��@� Yfhv����+:���mZ�l9���$�J�/��/�ĊQ���U�y[�2�.O�0���J�17��0�%�ҩ���~��-C\��Aj3��+�$�<���2��cU�'��~ q�d���ҕ)���q=�;����r�ǥ���V#�k�:E�@֙����b�e�&r���ҚfVDZ�L7).�=�7cY\Z@��$ЄQ�m(�TUę	�I�S�p@�3�Q�S�CL%�,ߴZ�Sf�W�C�r&gmk5_
Ps�@Zpz����AK����L�[Z��=��]�(��Լf��ln~C$�q��P�o��>�~�ۿK��]��`�H�D�!'D�L�.��l|�����O���f>Kr%�"���ZBO��NnBo=~�%��w��oT��Ή�?�H+�tQs��ؐ0f>�2�������Ì� 0����9��ih�6�����{��Z���@�"�j:�����=���tzax pz�l[�����=Æ������~_�>�5w�kUܼ�ԍc���k=��߿^k��q��&7{��=�k��L�Oپ�h��Wa��1�����&�C��-�p��T��e۱L���z�'�_�+]ٚ#�?��$�u"_	X���e����������?�[��__'�k� �4g��,���c>�̑��|lT��Gr�鏟�����{�ȑ �r)z�`)��Kl�
j2��|I�ҍhT�B:$�\�����eZ�uh}�3c4���`���[S
�L
+�3��y�/z��~�rJ(�x��YQ�%FI;��f�+;��ֶ	��E�f�4ȏX��W�3S��?��G]�"��iϪ���E�F��W�f�%$�Y�3S��/<I���+T:tq�G�|�C���>�H�q-ڴb��A���|��>��t}�4rN��m��7���.�_���^>�n�/)��l@)��P�2 ��=%s���N����i��0'�W�ek�i!�M�#�KeT��&�edV$iUʹX����</�RJK�3ށ�L�ȥ��z%���6Ɂ4��)�b���Z.��1,��}�M��f�uˑ�l2݀�6���^V�^}N��<=���Q�ͬFu.�j�	'����P��W�9ݶ�ͪ�8ǡ!���5�CB�,�'� /L��d
w[���t���\D���<s��#�?g�@�(?��!���kG�Id� �Ǧ%��Sn����9�v��5W�0���F�\ٮ��3�2PÑ	�x�+d����&<6�K��وS�����tQ�;�2�B�rX
�i���ۮo/�{.�6~���*�mny���T�����Is�3�\�w9p�d���FSqV���/=LT�d(�)�=�GdP�4M�����M�����z���}M�J&'$8H���)cH����
)���`PV[�Z-ˑ�V����IZk$$��$�H���z�}-�^v&�$ӥ��ty�+`ǡN~��n%��|�(7](�4/S�Ll�!ctJ��>o��F���@�d\T�����T�2�E�hLˏ��WR-�����~$:��%C�MeH��k~u%����÷��N4��Ȅ	-� C�6�n�x%ݺ$4�DZ�t=��o��phS&��q ��M�*�?�YAf@��E���3�zr��+tf�ۜ�6O�f̏��ff9��1#�W��E�9�F�S���le�N9|�e�-��T��8�h��s_���+�N��3��-/�����d�\��|��;����h��q8Tvw�nɲcBh��[�a�d*���5-c{������퓏�}��S�~�r �N�A��c�K�	!j���:��J�1�|��|��l!��v�ϥy~*�@O�l�_��?7e�2A�����ڌ�ڷ�����<����G������O��O>A�^�_+��E�x*���v�<U�8̸������ڐ��lL�y2'����GM.��x��������-S����������.��4�\Dg.΁�#B9�g٦����Ƴ�ș;�����5��G����S�>���t��)���)z��2��_�������9rv;3E��̴j�ۦ���`���S���/��o8E�����z��wr��E@V�d�X��PD���St|���-�x�%ZR3\��GEYN_x�I:��S�K��!��c�E��nSc�g�i�Բ�N-Wf�,��\/y��\�\�X����T8ҕ�OS~K�R,�"�	~����U�v�U�nl��ӧF�nH�l�*�m�<�kZ2�2И�X���S�LS�Ĵp���Z�,�r43cLS�&���<9�,s�˩t�:�1�U�������]�@���tp�<��˴�����荧����o���+��:�����C��:������6	��c�ٓ��0cm���2C��ѯ�$3�[D�wM�}.,k����Դ�9��I�<ՠ���L"%3Ge}9�.g�].V��?s�����v��ya�^qmiZ2$$K�/ȫ8�����0����}Z���l�T����̦MK�lz~I.Vmu��Ғ�'�h��=��g�<%�R~�u��P�.*峦.&���C�|��̌Ņ���6�GerB@:���c9��f�3場�e����J���E���$��i=�dV����r�.p�:�U!森i���z�"�MH��Ƕd�
�8�1����Ϸ)x�bT妵Ӽ��Tߔƙ	&������@0�ǲ�����U�Y&j$ݗ�rк�f'F��5F>�.�g��o#��N��7[�{���җ����9�%��6� ��W��� ���٧��}���S�'�	���m���Ɵ݅t�l���+j�5EsS-Ns��{�,��ɜn��0Yv9 �"c�h�%&�C�GcYLg$U(�}PZ[�&�L�K��mq�Q7���3߻�[>���l��WCi54	�6-f�8�
FG�z�8YGG7{�����E+�V#Go�j�}kI�:|��*�$sk�z.���Bx<�`��o���/�]g�w�q�I1�;`����5��m{���5h�f�*���j^o9�>��c���	"��|.,g�wo�ݳ��o�٭mo{m��n]�4�j��:r0�Of�����Ϸz�C?|���ə3g�����^ pK��ꭠ�o�9)0]9��|e
]�7��)M�|�lr�E��t'rbMS�K����8XH�dS�Ll%)����̢�I��t��+�p1�(�wHH����i�$�M!����<�*���Y�P2&��/f9#�����r�`0C?��y��=rG����U��.L���.<O'��+�G��t��|�Q:h���c�~���Pȥ��p�fT�N=���&];r�<z��Sʡcs�KW_�S�����M/���w�A����lZrЗ������Fn
y���FO<�=��tms�9d�ϰ?ࢱV�-#j�5-|��3��D��;]p��X�4�)g������JW9�,�␟�hO�_x�0�X�ʾ��>���&Tn���Q|K��]�@!S��Z�A�
�OC��=*�|Z���k.u���oi����{3�G�+��V�j�hqi9��ӵ�kd�i����*�EC.e��q쓮:2��o9��֨˕�R$��d�������tz�o��YZ�_�\�ii�)�i�L����f.^wܻ��J3�sԋ�􅧾LO�~���ݯ)���Iv��!?֖��~J�Т���|@>��w�8M�W�g2�D�o��y���.Xe�왂@���2�c�b��Y!��搋O�,�-�<j��N�����(���̳6��Ȣr
�z�!mY�N	B�E����f2< \��V&y������ϔ�quMK�i��A,Һ$�a�yd\�\WEά:���2�Es�~�t%�k�ȴ�T�Z�q0fR	$\�Ǧ���kDƲH�)�T_���PM��[S �ήK�Bӽm�J��@��Q�#A��nɴ���*�(90�ʳ��j�;&�����%A�[����'��Ԣ���̈́��W�KU9ކ��Z^��uBS�?/�M����eW:���/���sO���cƮ���3L���#�=���ȓ�*2��LQΡSBt,���Z�~��2K�0��l{S�JK�w2�pͯ���}��7*�I!9#n��/ji�$�,"�/�s���X�_d��ts�s3뗗�!�d�z��>�ZS�(o��w���V����(
=9)a�g,5>K��ݗ����k��0�6�7�WO������c2$L�7k�x�nZ�����M�_�}x��j�=[��xZc=Ԏ�Ŏ듘b;����9t�Մ4`����J&C��mp��/g��3�m�Ÿ|h9���G�����~�O~�Gt�����ԑÇg�,V��$�2��}�J.&g'e��Lsi'��A�8p�4�:Դ��9I���&Mq���@f��i].f�7� :CӍYk���� �m��AX
����?
��L�̺$E��o�����B�x�S��w���>53�N����ޛ�X�^�a�]޻o�W�����{��g�g�M�BJbYJ(FaCp�؊A���0�@�%[A"KQL˒l	�`	2͐"i���3��p���}�����[�w�������[� ���fwU�z���������}gL��SB������r�^���t~��&�x��i<t߃p�H��в� Y��'�%���x5�`u����>%4�"k���~��/�64+�ګ�ǻo��ɬ_>��X�fe���'��=��?�*�x��-����sZV�h5�yz��'��C���7����Е*�׬Fb�*�}hJ�lc�Ȉ7�1%��^����x���G�'�eً�,��Y�,zB2��p=h���,Q���\	��#?Q��c�X�]�����O�@O���^o_8�w�}]�ԋ�pd�8Ν{OE�V�)�q�}e�]Ω�t��ذ;P�È���=��5����bV��SO��S����a6?�w���%�q�U�$4�vfN�]A�\��DA��Dx�|X�[���soh�q�T��qIH�t�����>� &�<J�1�}H� ڮ~^Z�K3�uN(��8J�S�e�gd���/�!����u?M��я0!����x��C2�>me��8)��M�V+h�z�K)ӎ����3��#�gՖ��rw�,_�>5y�(�g6��7��6�nv[V"� ��6=��0g�	�	Hh��彷�Ob*��"0�Aq:3ݞ���v��y�{]�t�VAC̴��!-5v4��~=�J�G��2�vaBy=^��g=-���e��Zx`�0�-_���
Xs��$�U�`��50��"���3o����ˍe�9f����E!�CG֚��Th	9,l�
�2p����}��*+�k��.�Z����t�c�T��sِ�J9x~�0!�L����k��Z��!-�IB՘�7&��\����^_�広0
�x���Z�{�I��Z�}>&i�<��IT�#yt�;i��kq+�ت�V@k��n�ޝ�m}ￊh|t�Tv�[&c�R�����fо�u��q�fBv:�����]˔��;<[�I�"�ߝ���ax�y�8kI(�Y�a[M2h�=91��c�>��g?������������C��c�������'�C�tgr��	Ds2+@�.�@�=����ǋ�845�����X�%�u(���E*"x���!�{V��y�2he3dt�����5m�9���s.��rw�i�3L62��B�ƹl�fe��'�E��nS,���}���-ѡ>��F���'?��pē�|���P�����~Z-qm��u�ȉ�x�����b<t�4�A�	��,�`�M��)l�����DT]Ƌ8��i4Y�.Dm���A3
�֬����W����þΎ�`��ǎ�H������Kb7;6��b�fG7B'%^�'���^/����M��hFa��	s9%,�Z�peT����lAg	���Ӯ٬|# �$�C��`:pL)V��F$d2}� ��_ Yա�K6l��5s�(��{W�_TA���+p�x�VZa:�ό �ZȨ���<1:�QMHMF�?�
��g�S<:qD�g9��։���sX7�}#�X�߸7&�j��*�LI��q�-d�0;?��G1/�������ڤ!,�?��Ӌ���|S��\�L��ժ�0i����X�ɛK��m�͌��rm�J��{��^�����w�6`9���8��o��?��8��Ŭ[Ҍ�6�SU���v���;�(�$��eSS��&F_^U����^�����Z��>+=y�/ǡ�*��EĦx)�c�Ro���Ϣ�+��$!J\��B4��>���
�R�Q	��r8�ȳ�}6�7]��g�̿(C���0�7M����1�0I��.V$j\Ҫ�a��=8�@mi��g-/���u���ve�ժ��4��ŷ +��I�-u�s��tW�o�-�-�����q�C���E�4�d7�/�C=o>���Y~�l �Ԙ9☐��l��8�����/�1�jC��K���ᦍ��>sT/n������X[t�~�ϔ���ݽ �������t�sN�YJ�N*�N����Ljy�th��̇m�� X�1n��da����T��s���{�����l��_o=��j��Zŏ�<�f<l˾�k�0Bv��;��Nn_���w�6�H�2"�I)[���-�l���d�q�R�	� �?���8}���y���7�w���=�w|��C�����0l��t�=��
p�S�l�)�����g��?zࣘGI��a������u�\��O��>{�Ơ�0�nS�UWV���O��ߜ��w]l颣 ��M9օ΀O%*�T!J������oi��~���, K�����ױ֮ ��fҸ�A���P.M()�)�~��
��Wd��uݘ	��~��Vu�����z�:�:b��V1���s$���ڡ:B:�}@��i���*��Chs� �ȗK��ZY�F�®�
ī��|��>���M�x���6ܾ�.;F����SJ�(xfn�g�٢�+���͍d�2!c�BNǚ�
M���Z���Vb��t�L�As/t�r�)�'����,��m �+�2r≇��4�
f1��,�'����O?l�7�.�d�K�#���=!��N��:� �MYJ�=��ܛf�	���v������������!�ے�Lső��v�$!�6>�Bh�jZ-Ga�Y #��=4s�r�8Ӻ��?�>8_��g1K�Ć�'��V�J�n��l�g��װ�fo6-Gaq�H��a~zt=��׿	� �K�L���A!Vh6��/��Ô �I,�<%Ѧ�7�+4r�N�G*�6�����!����g)�O����������NMJ?Pqh�8���M��k�J�,��B��Fs����}�M����̤�DE�|��ݐ#�+$�J�ݺ�Z����#� Om>	'I!��V�[��\�e�c�B�1��%[�\{Q����S9D5!���0�YZ0�x����k� ��Z��E���$.y�����3j^�d*"mYk��!A����W��8{T��qG��!��24� B���k`ʸtd)�,��24���TC��)K�S�]%n�m-�[���J�a7�䑑G��=/��C�9��n�o˺cg3y��ʙ�;��U0��;u���z5���J�^�r����U�w;�o�Y�(ӱi��N�n�|kt�7ݴ�d�ַ�ov�7d&�,��c׮ڔ-����QyٶS�z�8�B? N�|{nnn:�N?y�̙O��/��7��?�'{�X�c����#7����A3UHe�˞0�J� *v��B8A��S(����) �rY2�tR�mjvn֛�d�N�Ǿ�=�0^\}�� ���8e������K��PK;�&u��D6t.�v� �P�NQ\-st� o^O��Y�/<�Q�]���|�[�k�5Zh��
�h���$�̕�\w� ^���lJ7���
�g��0��2� jd�N�AQ)���iG�/�*<F+��H
Thm��؁�:�N��d`�@,�0��H%����=K_H�>:����ss�K�?�Z���'@q�-Y�F��0?@>����nw�n�}D�u��P�H��h����dC�1H\Q2O��@�LF�B��.�c��nKǟ�x�L M �3�`e�$�d2Z���ݡ��Ҭ������=�R�m�B���,L�z��*zTnt��Ss��ӟ�qLcY�kd:�6Zroi1Te��a_��Xb��8o��Pc��n�Y6㕊XH�񩇞���wpmc�2	|扏���!�Y�"ﷱ�n@ ˄d�{}-�R����~�Xic�L�L�����Y8py�������7���fMɘ'� ;�P�Dz��E��v�d�@�=� d��tz=u��	�e��H�ھ�9z�B88�8�x3�s��q^��L cM{0�'ȹE�}�̓sAݱ�&Rϵ�d]��V��1}���~D�*g���hf�ChI��)�'`��qMkf��s�2h'������"]O|S���� �	��7Bn%Κ��>;�a
�qč!�q
}�q�?y�M��=�#�PO�Cy��7.��3:^JǓZ��|�Y)�1�]�Kߕg�	�����.~ԓв8#�M/i���ǔϟ%�羯Y�P˭�60��A7z��3��"� �q&���K�Y���q����jd�B�yǉf�){zB�����@�:�щ�T*Qv�_�mqם����@�)�2h���IoW�ܯ,#H�e7��_Ž�論�� ��dF������a'Ղ��[��N�}� ߾�߶u�5��SF�	+y�3'��݈���J�v,MK�9Li��񤡉���M��Q�SSS�:��2�����h4��?���3��c��# {Ǉ��E���i����tq���Vk�)&Mg(�M�R[��FW{u�dA��oEa'7>n�^V�>�{0�O���@ B�����_���*��o��G*�T�u��i��TdJ4(,U`���G�h59�J�!L7�JXG�h�*�"��[ l��^���Z��}\�|՚��g��4&'&Q�sec��'������p������(��U�ͨyZ��OZ#Yh��#gNڈ��ȑ�����*��#d^� sG�c�����h]7�S��-#J��h�"��RrgE�j4�	�Y|v�� :�r���}3s���\�Ɇ��e��Z�z�fNx��n�a�������k��Q�Vdt9)��Fs�-��C�a��K@ecG� Ft{"5�k���[�e�ڷ��e��G:��{����$A�V��80=��Ƌ�~�vC��^�.s+��(����c(��ui�+�����[�� ������1h6�|㚖�P�@�+�f�W>WԿ�垷�m,��`va=�(���|��r��1#D�PyV���a�����Im���x&�d����6vP��u웛Ci���e�=�9��J�K=���˵7en��Y��|��`_�������{/�ҫ����ۢ���y$�m!���j�;����WʕP��`�@����i�kv`��ۨ���	�k��H��t&IJ�	��$��y#�j>B7�r�P�NJ�:�`�O���,plS�u"2�q,��� Ka*�`镂%�2�D}52`�D�,A��cF
�I��H�/�ڑT@~����������B�'�:�
�iV�.�r���:�O>�,./��̑Cx��W��o}K��T��c��}�o�����wݾ�yY}�G�jw�~G�ľS-c��2ϣ��ш@0�f�>ǁ�D�f^Δ�1q"��>�C���5�h.1�F��ɖq�3 ��QR
74�ͱ����	�	��Q�BY�"�"�i�zSi�K���D��A��W����ة�j;��Mwq7�Ý��dc�a0�k�̊�nǹ��h@p���E��L�f'�1����g��Q�?L���:���Վb�e\<�=0,3����9z���{�w>&��������W>����a=�M�r�|0�&Y-3e�R�+7��W�Db!�O_6��/���j���֨��"��c 8XoࡃǑ�@#oW����+���rP��B�X�q�����t��J��� �4=u�a��'�-?���*#-i�`�e�|�*a����&u�v�d�&1挡��v�q��d���N?�c��(����h6�h��
�
�;��ǯ�گ�B\����O~�3s��ȱ$�Ƅ-��� ���HKθ�[AR�.�e<Z�D��� jMH<�2�vO�!�0�㛨�?5��DF����L}='�SuxMi��Z�)�%wZ��\r�A5��)���R���b����t ��k�I�&y�;�"�������4̈�@ȣ�}���_DS�E����(�\Z��,�ɳA�7�X��0�B��^[.壵�P\���q�����l���7�$R���Tvxr�R��f0=#�]��|�/cffø��W>@�YGQ��cE=�ځ\kJ�Ӯ]�"�c�83��{��F��Y)�O�
�p��Dfbg�Y-���R_�Fc�O�G{^�Ͼ�ր.fF�o�,�$�x]���VW�У�`��g�::'[&J/ d<5�S����ʒ�a[�ʡ��{�˜���y��WP�%$}C�k�Y3م��ˀ��������nW��E�3Bl�b�C�u�a�G͌�+�e&�YƜ���M��t,'�&�%�s&��+Ҏ?�r�ϢYR�4ʣP=�w\�ӝ����b��V�:[�f��a�e����!B�#p5��,I�4�j� ��Pѹ�qNZ�Lq28�py �r�s0�F��)�Ա��֐A:l��c8|��rY�[���Ԓ��"C9��<g�Q	Iu��=�ϛ~E�3�N�s�Y����t2sd=�l���{f��˟elN�[�����k�M4ʭ�[�=����2�w��kt\j���ڃ�FS�(���M�9��v(kPa|,���n6[P2�b̄,�%�=�RNe��1�S�{�H������ҫ��Ý����{%9�#k�E���L��6�g�(|'�����k�>0�f&DK �,�B�igTxy�'Ӿ�h)������i6jK�������m��j�q�3�j[�qe���xBT#[���+��*�����W��;>����úv��B�x6����s�<\F���,Q1;�C7-�n܇�up�_ƍ��~�1;��O�ؓʹ��q��bv6�v"- ����c��g���q��& U 턇@�J��is���=��Ji���-�M#W*(���w��Q6u �F.��,��|L�P�*Du������T������p��1\:	W/�����4\����@���?�����s�XZ���t���O�u�Ր'�r0�>���@K%�%H,�ac�{�IVI��w��34sNOLyЅ�DA��12Kj�'Sd�q��w�sfCظ0%�����81;�󽄔�T�`��X� b���)=l��f��f�°a^*i;�RJ
#Mm��9ы��V���7�c�Gw��]M���
�!
�2W��8�Bl�8��[Ĥ @��Е�F��k��.�o|����mlT.Ñs�L�ul8�$N��g?�_3r�fx���֠�p}�����V���{B*KccJ�If��%5�����ׯ^S��H6��������������f�;,�8��Jm�n�V/"�B��%����R1����T�֕�|�BR��O�H��������fh��Jp�8�����xTz�c����r	!l3�jr}�~7��Y�t`~c�"�W�ZU�7/s��(\��B��&�k7Qϩ�}�\�K�)��Za�3vF�gd<"%��(��7�S��!��#�ϒ�.������1�3	��Tg��Q��|f4�A�4뙒�؃t�������V��Q��B�ѱX4H25<�;�YJ���0�F��@Λٯ� ��� �n¸�A�f�@?y�ڊ�}�\^��ӏ>�D0B��o|�~W�&4��6�LD�e<�x��Ouh�'9)����1K�˘.��s��B����[���R��m��z@�n�,g���?�5�D�7hw��t7����v�j�Qf�4�>:�1�����X�A���|�#��N�L*��{��6��4�����^�0�s̮�F���-���L���`TV��{�8\m=�i�N4��v�}7���zh�l<�����a �I�}۹iO�8�Mw��\x/�s���>���0��Ѧ]���`�un����=��4�m��ě㐔��#�
Si�9��>�`��/�x����ɟ�w�t����Cy��_<�<��EN�����0�M��MP$]�M�7��=m`�b��X�e�%?O5�ab�Ƙll7T16ݖ�ܥV��>�S1V�>��h�����&���Ki:�o�(� ����墖��	�	AZ~A`&�e63d� �I�X2� H��@~Ro74$���o����/��Ս���2�3��V�W��w^�O��^�#�� �pV.�(@��j�Z����0
9��C�ub�7
g�@�è���9덚FH�T��Z�0��#�5��(K,J��B��$��"+���#w�Pu���z�ǚ\mX���f�A��!Q٨
���f2�^%��a����f��!{��g���^�_ž�yL�S�⑓�eg�ʉG$2n��!�e0��/�X��cB��LMcrr��1�����Whnl�ܵT�� ��%���TRC���f�T��r�"-�#�4B8@��D��!$g
Ս��X���5�/m���o������y��糎���k^Z��)~��yu!#O�i&5ݲ�֚��(-���=uj�Wo�s���0���c˚�1�fF.��z�����u���LϦ�#��Elu�wx.����Ֆ��r
++ױv�:�:��_ı�M/��ܔ��>�B�Z���D�Z2gm���g�n���=sQ�(����;	�P^OC u\ҲG�,,�S�+:��g|��Ew���tl�#�]��DC�3y��)��Ӷ6f�@�(9w:��,p���Z�2�A3-ۓ{�/5�ؔ�������xߑ�j���j�B��FH_�9�g��
,�ʋ_Gܡuw�8����'y
����9����x��q���{��h��iLH���J�����99�S�oj�Hs2&A#�XR�.�|-�,D�[�L�����9}nI�՚j��ьժ�B����U_��y��}�q���k����3���le
��<r̭\I��~�����'k���L������dr��=ehF �Y0���PŴyв3X���;��m��v1�2��fmϬܩ�^����M|��N|3S��ym^ᖒ��[�7��f"llC^L���J�6� �2��g��h��<c6r�Lf�א,#m]��z�����'���^~����o�����/�F{�={d��P�̉�G>-K�G�q�2z���MN�شn�<����=[i�9X�J��u�����p�.���h	=��Ӳ�0kc�ob@+Ή*�>�N�e9C�й%�"pAu��pd�t
9�<c)�F���]�����l$���p��ꕙ^x������\]AY�OV@H��j�+�Q�UojC�z��5�lȷ���K6#���S���੓8�0'�}JA���%j���1��9�Zۉ'4��	4��]��\L;h��˷���k	#߬��S{B]mXL�Ls=��DJL�E����Fh�B�vYFա�U&�Ri\��K���!�Բ�DI5�1[�dax��:%�5�#ԅ�>��?��ΜU�����}O��x��i^ԳT� I8�-bv��+%\���4������*J�81 ��TPc����oa)�
I� Ẉ��^@(ǈv��U�+K��T�_GQj��
��h�ba���%�Ĉ��B�ᐙ�ƍeT�u�)(�M�F�l��6��d(��F����u�Bz�*ZB@N�9�C>����q�s9�7���_r,;=�^\<(����ƌh[�*������t��Ǆ�ɽ���B�O=x?�Ú��%�_[������*��m�m�.����A~����>�]�������biR�r����G�'�&̧e��J��~
�V��ܔ6a�y9�hf�ؕ���=A�L�(c5�5!�/}�U,ѓg���Ԍ��كG�w�G�/�M��#���&7�}C�L�8/��&8RS�D�D�B��ĤUo a7XR��&�ͯ��o�z���k��Z'oX��N�B��i�b��i��	)*8��X��+C�z�1�;{�Wnho���zB��j�,�nj�e�N]m�5�H`.�דg�R5��q���hƶfn���4o�K7ܷi!Ͼ'�>��ܭ��{�`�l�%UA�5��kz��F/g�n,ͼ���)P��۱����A�q����ď���ԩ��IT�5el���}�(��'J@(�ˊ��Kܭ_��fhߌ�[&���ة���2;[������n��>�k�6 [K��M���[3#�R�ѵl-��5���k"n�	�_��������Q�󻒭m�5c��{�`�6�%ϻ;15���ӧ�����<���=A��{d��P�jӝ��{J6��L�M��_v��`�֖��j��$����rC4�I�ci4�]�@�U������ ����k�U���~`)�A�)7���+�s�r(�M�+�K�7�)��k��ѨOR3L�,fh"}��H�}<��������~3�������g�Ԁ�_܀d9�1*8��5�83=�ӧ�HcK�Jql\�"�*T�5u,Y���Ʊ�%��(|��u��[a�Hz��W�%?0��b3�)6(�H�2�p��`�IOK�ᡱudó�Z�ؿ�6}&��Ֆ��	�V� �Db��J08�C���r=�\�`��v�f4��Vv� ��g��A�q��ig�\Y�������W�y�-͡�cvnV5)� �Pƈz�ɩ&��FQ2�$e��?��#��*8r�(�g���ߏ~.��]�>�����Er�E_@�>��:Ul�\�!@/ '��S��0��q����޼��y~ڰ��P:�%�+�
�|p^����'�
�\�l�R��AW��#`�Z�@�Y0�JP�k
G��ة��o��e�����$.D��HtG��㴖��������ץ^�������I���_�t]�0�#�q��K���9u����r/=L��d���tnU@fQƂ�m�2��r:&z.s�\������7D��9�[�<���zX��i���L�Ф���oF:/�Z��C[��xaK��77���i�2G�c#'�p�$�i�`�j�uic	�6(T����	�Y��a�ň`h]m'�{�Z�w,��l��S�}���/����	K�Q�/a��&ud}�"�֯iЄ��w�.���i�ī^Ga~�������7q�8#�yT�4'��_��5x�X���`)%�bY�cO�f:���Y����C;4Ai,���"�n�n"<7�D]nu�\%)Cj|�g�<�����hǐ�8
}+�z�	�R5�_�@�H;ͮ:t������j0i'9���Ջ=S���FMI��K��eH��*x���q�.A��47��;���K�N�w7���;fu��0�6�ȦX{�e�	�����
�no�hߔ���I�Β^S&���d��D��m%w;�{��of�L�}�=�<xp�7��wr~_���hYV�����;>���kd���iQ���������*���}ҡZ���$�?.8�V�U�Xt��
t��\�����l�Y]�XK��y��K��μ*#fd3�F������ص�9�7q
�	�m�c�M�䍍��[}Qg��'��M��1�p�]��*&����3��R����潌fEN�>���#X�^�� G�05ݣ�L&�j7k�m#@��h�4k��*�Z]��T�M" �2fd����1:Ϧ��9fc�Nʑɴ
���uu�aT�"�N��b�� ���D�?��A43;�vȱ��!����4_R�H��]�d�����ݮ�x�f�
	BH,rz��e�`7-TV�p��ZƦvªbr��c�Q�PK���S��Y�b&�ɃE��,ݙ�M`�V�NVA)Q����n(c�Bk(������+��p��T��cc�L���R�A�FrQ�0^����jy��|�queY7O�mv��س�8E�ח��0V@0ha���:�
�^�I��GԜ|������s�~0��3h,���QK�B��*�����ƪ�05;������:��\��Ǐ=�)ܷp�q�ǆڬ҈��Je,���]T�9s���=R٢j�ҥ4J�"�����4��O��޿Z6|��_0�Z+f!����M�>O���ڨ�)M/ ���a��
q��/cq~��,�E%��c��ҵ��ˀ+�*������]��d�4ٓ�r��Fj9~��I͜��ScK��)�%������cOᕷ_E�~錧Q�]�d�R�x.��.Xt�t�Ȫ�4������/p"����~j���_����SbHZv��Q|��x��w5(Ò�4�2g�x�-3���"����s*0� |��P����P�y����ؚj	�eD���Z�Y+9d�Za��L�B���h�G"J��e�$'��@]�"%�Vd��骗I�4����z㎲�ݖ)��2���uSh���җ"��
NG"�]ʱ�:�|߮#����������_�U����w����$��N�0v&T;�Ϯ�ym���t,�!Gb��˹��d��h�w�X�o�;y~�64��E���<��}'��[/�%�����6~����������w���# {Ǉ����������mh�f<O����EDpg�䂥OV�iX�;�Q.��Y*���7Q�������^z_~���\�qÈ=R���ߞ��`���M��^��q�\]M�C�m �<����:�uV6ՙ�I-�I�)�����@6kֿ��@�8z���Sc[}�}��h���{����������+8�� ��fU�1:��f;\ݜ;r�$R}�V�E���#P1�Ȉe`�H�ua�q�J�{�?
Ɨ)DW�����ۢ]��l� �Z��~��ՈP`�U����Ç��(Tf~F@��g�;@�C�QW0L�H��,H����U*f�b��k�1�$2<���~6V��������]�9%u!��8�<B��zt��X`t	��--/)�e���&��]�N�j��iփ�v�����C�����r.U��~�bj��Ө5�:��L��3D�ǒ{K�\v?g#9GI���c�T�q]^_S�v�%D�*�t�۪��d����|v��񌀽���ݵd��{�Qx_�oə�.F�yM��T���D%�O��pʽz��o���ޔy�o�ȧ���g��M"�FjĐ�K��U�2��q!!�R�2b@��*�q���t���E�7y�׮��w߄�\����~	?|�)��PK).\� �����1��Y�b��ex����9LO�`bjF�������'�n�-����OJ�	��3:Avұ�Qy��}���Mt�j��i�p��1<��c8|hSSڍ�����r�(�b	&��Y�OBJ�|�n�Se����dH��F��rQ�k�V0�b������WP�Te��a|zR�yU�z��iv����Ko��BJ�6	����O�'�W�^�m��n���E��6GdTZ����Nl�k-��s��	{�hO��8^%k�-���a���	�I�^N.}n-ӫA�!,����H ��Z4N�Pt��[��	S�|-�d��� �8���F*�dsT�nф��w��|��w�rl��E"%��2Z{TR�Wx����m?��u7��ݾ�wm˿����I8CK�
Me%�s���4(�Eډp�p�a��xn���E��ݑ��ﾟ*���{�ݷ^^�
��;{d��P�\���M0��ڑ�F���-�/��K}�:�Ď3f��f����)�/!L		��~�*��s�ܬ��t�*�t=K�W�;����@N$ "39��XF����?t�븺vIA>�j9���S�5�yRX�f�C�NZ����Ǭ�4h��Wؐ�H	Pc��з��Zv�F1?��zb�4@4�#���n^���wq���q��I���hDZw���C�O�P��g��l𶯶�$Vd�

�����"�i"fǉH�u$ifIK�F�о�L�ItW�H`D�G>{:Xis���,�})�'��{��*�NiiI_N�i4ꖜD�dx�Lkd�R�� څ"�Q2�2��d�s�r{iQ*��������#L�9���,�4B�<C�!�6y�]Ͷ1Z&`geyɀ��)�;w��i�G�#Y�����\c�� ���р�Cr���}�`H�SO�-�=&c�kR��T7*�
-1!�`)Kt��p_,i�G��7&�%nl�)绺���l]��>�{M��u�B��&<�-Ĩ*7)���:*>_���=�5��t��˧��X̛����tV�n���(�#�X�?�_����̔�����*@;`O���]�0�3^W�aΡl6�V��S�kf���j�}:R8�,^�u-����Q�|�"V�p�o�z��B�����r�P��gz�����,��o����'g�}��\Z�	!s��Ξ=ctO��B�4��QS�õ�W�6C��
r{�>���C��i!|=I6K�����p�ɇ�9��s�]|GH����~�G0s� JBI�H�,Z)G�epS�Slz���/��w��"+�wj_^���ȔWrL��t����|��8��,z%<�p)�W�'g5�7���ʥ����O�����*6�W�{��Ɏe�-��RMѾLVY���岺Qcš��E���N�9���^��c}� ��u��=W�5�-a��5㤂����|?��@K�)iU���2�<�	�ܛ|���=2���iߪg���mmZ�n?�-$bk6�^��w����wѬ��9۳'��vt�!v>ϻ�JFه����J�B-ku�|��SvR�|�ҫ��}�c���vgwX�9�?5m&�R���<Y٨d�w���# {Ǉ�(��6
ÀF�����."K��Q/b��^�G&JQ,�
�u�N]�5�ހ�*ￊ�8w�"ږl�l��5�~�31����w@�].
���]K+���.@�M7t�t:�kO��pMm�,t)��)
2@@N#^��ع��7���F�'oW���4��˚]`��AVM�T*I6!�v�����n�X��&h<���� \f����c5Z�.� pe��AAj0:�X�9݊����H�fa'�lG6��������t#!B"N��+�$����I�~t{
y��}I�E#O,ɠ�"�e3�h�%B.�u�`�^�����F�R���Vn�Q��2�aߔ�Da�D�d�&�e�$g>8+�RG��C��E��Qd���������0M�}��iI*��)c��������1{�(�u�x�ױֵ��$3���J�kZ6%��!bp���
����|�Ւx�n���v&i��f���@W��4w@sL����3�J����	�ԕ��  <"��
F�����$O#�J�H��1C	-KbX������ٷ�ŕ��o���>�d��	X_�r�}B�2y!@)LP�.�@�}Z�:J�X��5(Y���ϱv'gj!"�1lr�JhU[���P*�+�̍@Nqy(�j]Hf����?�@��ﾌGxL��/�k�1�q���듵���c��_�o0>>�_|_�������'~�'���o��o)�����[���Q���}Q~`�<��w�T�XQ�g�D;��N˽/z�67���(8����Ԩ��y����Ј�9����;{�F��P�]x�yDi[�,���U֏����lq��?|���SObzf�n��:��'T�i�]E�E��ֹr��U|�+_A����.��y�g�#�ج:B
"!,#���C�KD/a�F
��F�e)mtH��l��C
�1�vC<L�l�2����qc����jP�W�WQ�Pܯ��CyN��,�(�JF����ٶ�����Gݢ��v&;�~ �>���b���n��;��?�G�Ն�Y�r�Dj�ߣ�Ј��K^|kwtc�lʠv>�D�2����^3�o�NP��LJ�n2�n/��<sne:ڶ�! n�Z�w���# {Ǉ�x���S�ι_���;&;� _�YY=����D��W�
Y2`�)A���ZSL�֏{*�eU���:��_�MnHP���]6NK6����	�r'H>J��jd���+K��n�þI��'Y<�hi�yإ{KMž��T�NB��6��],�d�ml��
�)�}���5;5��F�N��"��������^~A�p]�������G~��(���ж��"?=�~��(D�Uu��&&��J�i�F��kLkS�b���4J�%`�������2��T��hI��H���@gv�d�R6�޹���	��.$Wb/��[@p7�`���{�$��j����|����}�~q��2��:��)|�[������j��{��ϱQ��'�E���XA�.r��܋�[�����p����\�}|p�<JS�x�ɧ17��Z���|����?�=��n`��eyS����M�5�	Rڣ�`���q���8:[F��̕���el��WBSr��kia�7�`О��S:1��!�F�75.t*bɛ팜���/~�L:��! ��I��%�$�Ck72���7���ߺ�����%�\OK�fЖ�~�^� �-!��}�<��s(�M���rC�[�2����s�U����Q��h�嫀��f�2O�����ĩCHM�������BnRz�,�!���u�����a����`a�;=9�����j����p~nNa����3<��S�r�
>�Ϩ�����?�9D�+�򏅠���ԩ��^�{U��� '��ꜵѨ�h�P,�/c��\b��F�*d�v����̧��4Y��v)��G��xIK�bY/b^�Ú��lNN�:yT�|}fi*Q�k��h�r����}\��&�.&�*WV�~�D�Y�V��Z��4;B�q"�`�xF�\_4"V���`�K�n���l�J���"�Y��2�Y���Z~	�:��0�x�&���*2\�����q�ߍՁ��/㕗{;��3=�N@�s�H�F�l'ڎ��n`�2���$d���ܪ!�ڝ��#w���w"�|ޖ��I����ݪyH~߱nq��ӱ}�F�n{�݈��=��1& �g��0��=�b�N�r�}�j�ŷ;c�B�F琔��B�F�(�% �>d���c������^p�����?`����# {Ǉ�x��,^��_��_������N@�]��
��� YHdw�~-ub#+F23A|�3v�a%�F�1ݐ۽� ~��ټ-�eC�
�����(�dc/�\Da|��됁~�|	$��)Ab9��\�tӔ�������:�9�	sC�c��2����Y|�_��Z9~D�\N������a�����F�sY��Q�Ύ�̰���#ጬ�c��&ޗ���1&�gq}u�b	O�#Z�
�Z�p�ہKC�L�t�&L����HU�������v�Y�EkH�j�t-f��F��ha�MQfl���6��E%���̲���ub�?�`��B!'�Ќ'�������I�R��� �~�X}�[p�����TJ˔���'�LbJtPk�����T�ÿ������0>=�#'�#��8w�,B��Lk+BNCS�x�0f榅pL"��⹧����y!"3rG�1�|׿��j��(�O�U��P����`0Lğ���p��WѰ.�|C�#�~�������fb������(�|mhىz�����T/2$�2��͚7¶��5��,/cbaR��	d�&��Kj��4о:�o�ΥRC�O�3k�u�=�v4LVC>�����K�����}3B�Z8��;x��P�Դ����s�1���2����$z�O|�SB������L��KאY��ǅt��!��X�{20�XY��vXE�0�Nu?��#(�R����K�f��,�S����s�?�C�ܔ�������?��C�U�E�7�_O?���~�w�	EҚ��,�)��$���[B@Vo`�^B��x*�'QH��؃@3Y��)-(M� Gd��G��㮂{���	��Ifi���t����ˇ~O���[Y��]��F+�ٕ�Z�Փ9�{G����$��f����)�u�I{��E���H6-��`��K��)jV�﫰6��:�s�`��-y���N��A�%AqҷDFf�e��Ʒ6!5]�I�!7j���nʱhn�U�r�f���&{�Vм��w:�5�� �H��Z�Y��;�]��.����n罓dd�4�TXI�Ǌw���gi˹Y.�N�[^�[����w��h��M�u��E�?�f��[]����G1�����t�;�h�땮X��y'�c~Nh�C?�l�<�2_m��{��Ͽ��'!�Gya{ǎ��;>�G��[��g�M��t�v���(ʩ6���68rl��d3�uǴ��Ҧ�&p�H=#�`7q"�,��E�=6(��ȗͮ#���-�� ��������s;�4r3d��|n^6��İ���FE;�H� <�-d��VEp��o�����۷'�3X��"���[٬e��V`/:�������L:��[iO˂���-j4�R��4=�\i�����z�p�|�a�eh�UE'wvټ1�k����3�YZo@��1�?�p�Q" �=d�� �B�6#Y��Q���u<HfR�T<,q������1c�����H[K����~=�7>�����1:��/abrR�I�_�,����9��-;��ɓG�pt�vK��*�:��:n[u-<:�Y�K���Ϡ�����꿃3Q��BN}�����*� ����Tf��DW�̔�F�dF�S��B1�RmFKH�!�t�a�(��A��X0R<��u�1��e��2�y!˦��5���k*H��Z�~R֤��V^�|��n�J�tLG��潈�6eĠ�S:� ���ĺ,ymV�Ű� y�M~��������f��}�?o��u�/W�����?���qߛ$�%y�z�D�9$��wr��k�h����\f���|��#�#%���[k`m�R�yw=웞�-�7?��G�cc�.�����2��m�y�~�Q������o�&fff���w_����3?� \�tY������xY��P=V̪��^��ɟ��K��d�$$���1�9�7n���W�0Cl�1C�gLu�k�A�����A�Myy�:����cd��4������D�FV]��@V�Z����t~DC-���8�#c�0��0��RF�q#��)65af��j�о��c�b���?'�
�c|��CS*�פݴ0F����` ��dF����nRJŬ��(b�v�N�tN椙�I����G�["ߌ�k	�.�{�6����e&v�ٝ~�^	��߻��ݴ[3$a‷ۡc�E��,m'{�v.��!�p�c���6��^�m�B�ns�rn�m[]϶�Od{��Kف�GQ0V;���h�{������(�-�I�þm��4�4u�����x�$��.;��M/쇦S��)�3|����N�z ��b2_ _R�%Kj6�6ή_EۍБ�jF-CY�܈�y�ŗ�ғ5-`���+-C>�im+d�@��!�N9y�zU�� 5��~�u�Z]�6����6�u���z7z��S�E�t���O���)�X�9/�X��{��&ӆ1:B��"�1��@��c�6"N���W��a�~D���w��w��+���H��&���ڮ�X���%ݡ� �5:fjh�F+���u���#�v��V�`�@�z����N9ZN�5]��v �㎜��䄾O�� ��P���QM,D#��%�BfLɞ��?x�j~G���İ���Gz���>��\���W/���/,]��5!!݃����R�>��/��[��P����^c{im0�h��,��\��@?ND�l����5]��Y�~�O_ô����mۨG���M;d^�Z2��J:�jܴ��g��6�f�2�$t���>6�s�1̲.�sF��zjfU��~�lA?;6.\<o:����g���@Xj��92᥍����f�.�w��W���zO>�>�c_�җ4c�R���~R�������&)3�4x� �V�ї�MGi,8S�?Iakd���H;2V�W�����������#��an6'$��Q�e-�~XƎ�Y�3�����]T���+��=.����$*$�,7b��RYWѾvgd�ڔu���'Ƌ�ȡF����q��!���55���73�|~�0��7f\��J0�~^җ�}m�<Q��=�:2ce��W;��ڰ7�7�����s\ی�`�ٛE��؏H�3[֕4�L!����2Oh;N���	U�É��`�
+8����=L�EZ s�Mi6T��*�2�/�̊f2��v�H�e��ɚ���4���^H�a2�A�y�2)�O�
-BY���g�i�y��&�U��n����\�@����[H	#�V|��7I,s?-�Zf��ة�i������)#��q��(�o��V�1"w��}����U;2ʔ�_�fѶi[��viVc�W���}�5w�hm;�qK�8�}�ޤ�i>s2Ϟ~�i��_�˅�~c�9����;>�G�R�l;F����a@�,�y�T�n}�^f7_mj+�����P�G�wP�\E3x���qb� �_ʇ�[�\�2�>| Q�Õ����eg�e(���)�P�r�(�}�U��țv�k! N �Q>'j��ASޣ�R��u�j5�X[YW!%S�t�aɓ��e�di�Q`D]�X��ߗ��+�'�x����ea������,�����q�ڍ�4Mm,
���Q&!$���m:��{��#�p �G�Q?j$��cҚ���:�w�����f�TOA@A�CzҬ�76�7a�R����4��%�3��L�9��>�z�r���5'䋂�|�����Y��o��.(1M�Y!&y�>�5ym��y�]D��t+�x�	�W�����W^�׾��:5,?�by��ѕ�*.��R�F�o��F�ƥ�AG��%��.�G��u�r--��m�n?Pƒ�A������k��z���N�,SŌ���і9]�N+��H�s�g��&����ڡ�35rN,�`i�+d�D.u"'��X��h����OmN*�Z���o��̛��M��Eb�m$�6��Hj�{�	|���[����>��OjT��n9�j�UyzF��r��f��ϰ;��Mk�?3���8¡���Ҟ��K}É�Ǒ��M����y.��T��q�VƔ��L"��x�Ǐߧ�_��_�k.P(Ά�ce|���RH����b�ưII'k�YV7;+��F�e!�r��ZNN��c���_{��ĲV�Ob�G�jt�
����Fd���.�R1�~��(��q��~���Yh\��c8m�/kB4����
�4���L��/K�r2������b�l.3Mbu6���L#��b�V�+�nR ut}C4e�d٥\^ǀ�rY-�	�V8���5Pb�e\�PyHT+ƒ=-ñ���| �X:��2h�U��)�#�-(�J�LO-�b�1O��8��gJ�ubSz�B��8nm���{��u�h<��K�V�q/��[��hMny�7�c�t�7i�N�b���N��g[�Ǵ|w��GV�YZ�y�[�'�	FY�݉���.�y�h��L!R�Y�4�٫#�y�c��~�R����?�#!�{d��P�_�(ԡBH�K������I1�s�ҝ<VPrw�Hqc(� �	N}�q��O�i�ʿ�*V/_G!e@�n>���do�\�򰋱�3�=����߇�����6�j[iy�3V4m.����4J>!%�m~,��GQ�|H��T�B]Ha��=T�%�!���F�I6��P�@PO� �\��d��?���P���ry�3*��n6����;z�	��m�5�Ad<�C�AxNZ#��m;�5[񱧞Q��l��V�ȹ	A�k`�7����( ؖS�؆|��0"Y,�'�8]����)��bi��z7���th��S<O�`~�c� ݗ���g�4��YҞ,q�Q��t���1S�(�����E��]\�TqaE�[.���aB���w^@�-J9\e#?�W2���t��]s_�sh�赻H�φf-1��r�u� o�� �X@Y ��#��)��ƅ������T�*`b%ZJ̒��l�H�si_	m�q��ȹP'3��RG�σh����e]c5��#Z�2�(�$��$%N:�ZoO��hf�<C�"�t5��M�\�PP='�.̀�K��Ԕ�F~�o����sZ����p��5!'���Ӿ�O,��'�y�W4�4�ʘ�e.��`v3EA�fm,�A]![���sR�*���Ɠ3�2O:C�<FB}f?�Iz��en��s��<N�?���oh��g��tK��L̬̕��w�6~�W�7�ͻs:����iu����!mtU��o	A�u����m.�_��%�`��`v��Z�i�s�H>Bө�"��y`:%dTHVĞ5l�~����B�ia&7�����%W��Y��V�sʎ�WPZ�%�x�I�zfYJ��W�ۇ�Hǌ.�̮9)C�X���BA����7�<�83:�r{�f W�6	��4[G]� ި\��mL���{����%�����,���2E�w��P�I�4Z��!c�j?�h3ä"u!�Zʳ۱� �V�m�'Ι�H����[v�^J��䂵U���F�n�7"����l�Nz℠����6�ڡ0]��s��&\�M���ַĊn�綟���s�l$i��m�`5وTgG3l��ؑ�ʊ�8A�3�����no���V������c����ccy�5۝z�#@1*D�@#vA��[�k�0�]w�~�S::
x����l�o� ���n��XS��Q�2z�Ŷ�>�C�y��,ceiO<��:�~��۸ּ7�VGA��n4d�o���J@Bj��2���fz����,k�� �Y��f2�Fv-� P�ڒh�J(�4Zu|��dv��'�d�sF�)�]�װ���%*³S!�-*��Ej�+���tq3��}u����0�{��	<��8��y\�|�{�u�8~�(P�zf�_��э�\����l"��<��wЦ�����eԘ���u-&�����$����/��;��nF�� Zf7(*�*D�x�ψ���-yρ|=�{\�"����e��,�s�����.�J�>k��m�X� O�e��t�b8�/ ]��Y����=T��FW����F���k0��W	�q "�غArs�5jW���u�ZMd�e*�\��k��\îfj����ZU�1�U��Şy.8�̬к����=Q�&�JN̫L��@���Z"AӅ���Jm]	NK �50�piy^��m��)�����_>����˚)�|d._�zEaF�Q�o���}�U�<���ǅeYպ����9���k�I�s�hfǨ�9w��?���^>�����J���g:	�v/�� Q��җ���:����ze����W/�_��vH�������
��߸!��:_�k��WC!��'䲣�2+d)jXZ:c�a�R��a�Mc,K����{��ګ�������JRCJ���bɖ��Bb����@ #��I�d�?��a r �aڤ�D�d�%��mf8{/3�Nw����{����Su��zfdYN0�3lvW�{�=�w��y��y�J
�0��k4;1-�^���`��^� �go�ы������Z|�W�S�9�ϡ����P��mK�������ݖ�֪�a���p*)U�6�+�q81�����6<]t���0ӀD:=���-��T��<�l4jC��d� aL�<�X*Q����D��SNN��T�tQ�ξ2<�G ��+���D���Z��2r2���)�$�˓���"���S�l�k��C9_����=������+�<|4��a�;Zj5N$>(2N�����>�d�E�;��xc�q�98{��?���$�/�EYJ�>bW��u̽~����GdE|3�Y1ۅ'���
pe�K����n��w:&�r��N�����:����u�\2�Cw89�� f)F��H�Ch��@	LӽvO�R���W�yoK
vB2
f���� #�Gu$����I�ߕT�'R�b2Y�R@R��_zU>󹟓��=-�7�Ҫ5�]�]ݓ@��+��\4�{T9�cP\�3��z��!8�t�Y�<#���r�Y9�zz�T�t���Og	F��v�8�N��C����eS�}H�in�a��3��R����DQ�%0��3r�p }�m�� �7~������ө�~�*x2���jS��%%]�ʦ�c>Wf�7�ۺ�3�T�Խg������\���v`c�ԩ�)��30���dR�RrBu��C�)��Q�������9�r�F�@�9��aP��$�� �;ժ�nm���Ӳ۪������wŵ}����e��~�Y�T6)�V�8�&�O�W�d��v/�
���z\h��BW��^�W��-�����S��OS��7b�'���|p_Q�2�!{D���2%�����׺Yݒ��畄���Ϊ����zu%V���[
���9(PO��2���D/�A�B�,
�csցhl�߷��!��V���y�$���MD�u�g/����QFU#��u���~��ߕT��2+ܧWt|=��S���ϰ�����ό�#��}��t�̲�0|A�i���N�e>5��k��᝔@�v
r�t_)%��	�O�eg}��n}wEJ�)�?5�5Y�ұ��z���bG�w�����R��e6�� �w��ߑ�{���H�7p}����,�ɟ���d��������,l?Hu�б�!A������dJ��������wu���2JL��%M(��=�0B UPâ����21 +�c���jcgMҍ��197sF�\�ѮWƒ��H�;��}Yϣ^k03R6���xe��/v�-�,�=�9Bυ�5z�1�B��$�'�-S�����n���"��xó�g��yv��	�$�F��8ϘgJ�҉,3��<�,Bgt(�ABjj�BAvv[aD>l����`6���60������/H$*e2c�y�>�z��1?Fؗm�e��~U�s�E���h��~����k�r8�p��y��7�;�q�2~(m���|h?4��������[��!����:������X �3[A�U�Et�:��d"���ێ�['0�@+��w��/4o�i����{_�����d��N�����򩴥�O��=;��B����0�bذ�.KcR T�o�uss���{ t�� ����}�w���iy�ܼ��k������2�/JF�����ʿ������<6}N^{��2�(H�h���%W�Ч=0����kyF�[�ۗ��5	�ӫ���^�S���H'��R�S��l!o��eY g �X������G�����5<r�F�6{����'���f@�Jq��PܽyM?{^&+����ܳ��������4U��nKL�?��zu�{�$�-�&s#���)����-�`Q�(���Z���U2�b������7��+�B����V�UNK�<I��С^ˡ^[0�D\�����f���we(�
o\�.B�z�P���y��Ƕ�@�X:�[��t��}"6�� �Gkָw�䷿�U�7�i	���_��[f�"m�,d�@1����X�?P2�s�J
=����T��~W���z�$'2�	�$
�翼&�f���XJ�%�(�J_-�\*�Df�Ƥ�<>\���υ)��e�ӐV=.?�z]n�mɛ+7�K�L_� P>�{'�f���r������-���A>���K�¨>��^��gh�����,�c�]�?��?�xͤ�aOB�.�-����u�����?�q���=@����J&�������.)4'�\�Ȱ�I�_��r,m���3�Yߐ�lIzz��&3+��E_� �ܱ����tzJ���9�l�Sr�*���^[���/�]���@ڃ���&	��֚�r��QS����\��K��b�!�i��{j��G��!Ȇ�5��A4v��+8�l�d�O˕SsRhR����뚝����i}&�R�^��ή�����@碞>���u[:6m9�X�gb�g	`%�Cd�|�-�{���b�B!�y	ٮ$ʝ��^8wN.]��l��p�2,Q3M�,�������F�hU����Q�D\�x�45<�̀���t��͙s�/�&�:w��,���g�B+!�'�c~l{�Wb���������#2�&��������O�~���dF�%�:�G�jW�%�  �V��T�up-�� <�����Zp�}�����Xs�~��a�\7�{H�]�vPq`��&׌O;"Ox����\�ܼT��zI�rB@ƶr�}�7ȓ��q{��k�w�R��1IC�6K]8�}W�P�҅6�@0�E+k�e�2����cy')�dN��	����������w5,p�iG��'�݆���۲�h����
N���Wdke�D�=�xy���c�20�4	�q5tY]H'&&�:W��y�ѣ�i�FͶ�2"����d��Huh�����'Bp ^(��d�E� xު�h�}�������3��~d��=��!ʄ� D�@2	9���0)��l�j27=+wn�f}?�%%���w�$��k7n�$(B)Ѕq$tcɸ4�-��Jy�^U��!"Y��wd8��1:�� 0協�$ h�7e�cFȌQ�����*��*�Hyz��nx�{�n1ڋ����0�C��A"FiP|~��Q��U"�ZDN����Į���2��H�0#���������yȴ�J�@�P��V�aY���g���=��+�������PA1��m�H�[��v���ʡ�&��Ґj�|�}rْ��g��+�A?P`M)�Rq��X����P ��ds}s��P����D�	�Tቱ��!�vO�t��X��RR��o�����ܜ������_������������^n߽'���d�E�����$/P9r��B�
�az-
r=�������R�1�����ک��²̔�dnfA
��,\Y��6o���^�ͭ-y�����'dee�٠��Y�J�67)������O��K��qW��{�ݒ�D\n�ܖ�kM9��'��y��U��٤��_��SϜ��w_P�a��Z��,"[)eH�6�M6��d���E@ �D���P2��ǉL.��U�HQ��D}(�AG������Oɹ��	�Gn��\�����T�j��3��ԕ������1�SVB��f���ml�H]���OH^�Y���y��3$���������)�T��L�T��1�b������(��ۦ�?����zC�}�a\����<#�9�!���~����$/����T�=�{������l��X��?r;�\*�/�l6���S��-
^<*�_r��N~O�(q#%�e+�Ge`|c>9.Y�c��΁�?zhXC��8����Й��ls�3�p��xj^��y�C�]��>�g5`��AC��LH1�E��8;�H�Ν?o߿�����vB@N���V.Wt.��芌;I�46 ��(Ϡ�#�C����+Hl$=T 6�� ��u9����N�i V��<� �ˏŕ��h��r��L���зo]ӅnZ��җ��ޞ|��Wd2���|Ev��e�ZS����rhH�g���L���4��~�nul��Z��.��v���0σ,%�̑AAf� OAK�X��B�� 䡬���둌3j�(!�#�
��� 0��߭�)��"Wj��У�{P���<�����
YY�]��p*diq����NG�=nyB��LONR�i{k[R
nY��C&�e�1B&�d�&RZ�q��)�W�ޗͤ���_�h�g�y>���;�ɞ�G���VPW�2�^��=���MLT��y��'�Lɲ�W�\e]:�n����yp�)HSv��K�$!�H��ނy��g�Y*�6/8R+�+�����v.�P,C0_�@Ѡ��^	<] ���$#���`b�ֻ�z]������0L�cӃ���jz��3Ҫ$Ö�T��;��2I��R��8N�!���WZ"B� �wIɃ����峒(��O�~���(��,3B�!K ]�pX�o8����-��g~�@���,gN/ɕ+W�~�����S��R �"��)�Y<��
�g�xa���}3�!At\,>�wI�#b)P���<�dcВ���ܽ���Ò\2��۔��ArS�/�A �pbo��N[	�/�XO�Ŭ$-�R��w����M,f�����?{-&��/KG�j_A3�(	}�>�����c2=�(���i��R2�/@�22Y���h�m*�89��'g�"�4~?hH��H�g�wl�I�ޚ��\����,yl�\�pEJ:G�T{���_e�sdѺ�볛ɕ8��KE����c�WwIO�^����,{0�S=�D@afV�PC�#}{�Y�cD`~LY?\�r����!�q^���9����F��u��]��K�	I筍�^�>�@y�8�ZmOf� ��{�L/�g�0��GDA�j6��-�"�%	���v���k0�(��(���mG371��)R��L��q*X�8Λ#�.�H/N���?�����x~o4&���爏�]ߜ����}d;� '��z+���±x�N+���l�����-N�RD���@�]�C���o��Xy�ي�
�'u�M�=< �	Y�x�b�fby;A7貂�[w���ߒꠧ 6'^�+dYt~�3B+��X6����-���j>[bT�XpA��,	]v��A�	և~�E��C˱7�tҡ�楋�ducS�#��[5�Ҧ>�M�
2 ݋�����3ߟ�Q���!��k		_��M=~O��@*3�`���Q9�)Y^:-�J2����G�����Z_e�@�a��ɢܬ�Hb������s=���,���N\o��?F�U^��-�˂�U|�1�2�2�QK�Kk�Ũ��fHG�|I�O��O?#+�^gYTN�c��i��T-���e�͐W�eJv\�k"�ȫ���}�(&�FB�!od�u���"1�gγA�G���ē)�#r_(N)�.�/K�A4y��Fu��I�(��iP�c�����O�ge���{?��|�?��JY�����5v���ץ������ɠ7X��O2@=ɍqP�3���=NLPYj@C�
F'Ϟ�&'K�/��T,"�̲(ݺ��Hl���1�ң?��?��߸J��ٹY�y�&A��<����+����|�~J�L/��G�	��a ���z�4��@vH��F�Fs<����y��	R�ި#~�c�^B�n���>���E��WDK���9��G)}k\>7������tF�����@�|Z��_����O�ͫ7叿�C��;W�85-s�is����g ��[�{S��hj��c4��h(�������y��񟏥dB�SA���Ԃ<�̧��-+)�q.c_U^�+>eD@�9��=ȴ�zUw79�^���l��qn=��,�z�D���H�h�M҆9c�>>,x����;Ơ�� ~ ˘�j�K���6I3�:'b��r���T�n���u�"��LS�(]ߩJ%m;{���%��sj��.:���# ׏�Hβɱ���<��9�0�~X&��\¿������q� �]t���FB؃�� �e@�y���7�O>l1����(�_|}�q��n����_n���K�?�_�W���L9s��_t�d;! '��{�CK:;H��#B82��(UAD �iwKAw���#��L:q(HV��uF2� ��Jd♤��,���:�u�I*�EI�t�u�P��T2'�W���������v���P9�3����xFQl��ЗN�eL��A�s��cD�;mdD`3'؏��O�k�'<3U	��fpgϞ��R����ʏ�x�5Д�U� PA�N�`��������+Ui���2U�Р� ��� ��ڸ��	������WH��V��:��9��������?�;��uP�6�

P�̥$�����Ĉ�kSn�d�h����Z�fCI]�eӰ��t����)$]AD��6E�Qb�n5HL�V�5ɖ*�q���,��ߥ�*�Ё�iY%/_�ٟ�o�������%���MF���(cIf�BD��b3M�N�#�	��g_��/>&�/�����J`��(!S���W��V?��x�`ܥ���H)�\�$�NO�,\��^�f���Ǟ�UBuK�dR����������5������8J�A�l����rT�a�XL�y�Nx2��ivj^f����Е3�����31it=���e�{4���<4zf��P�z�����~�7Z�^�.O<�G����������in$$Q�F�
h��3 Ԉ;����>�=}?���T^��<=i`h7[��x����]��M˩�3�5��1�0���ZT�JP��:����y
������:$��f�$��~��������|�%�x@~V�S}X�f�ʒ< �:�|���V0�����61�o��%J�hv���i�e�.��Č�Y>+��J�)Q���O��)'�a3SX����>{)��BE6V�����-�OO	2�w�P��A� �ZH��������*����yD@ג��!(��0>������is�@�$��P�����HerB��!	��!��$�� ���C_͎�:5�9K0QzȔ��r*L�6j?�x-g��C���_��>�����@}���$`?0����ƛ�?軏���灛��>����W;N-�c�d륉J���;p����ų���������oڒ�턀�l���nmW�yF 3)�a�R�AòeJ��:��tѝS�1(���u��D�_��1����]�l9��uo`+6��l(_�)����O乧���_�������:�� *��ݦ)��c���`,��m6Чd�	X���s�H��a�?�ǌ�!�$���Ɋ\y��i�. 's�2�(a[��t����j��|8�f�Ozp(�ս�5�9 �4�F�Fz�V�*�C�+�I˅����BXb�����tM�ަbj�P�p�es��~y���LC�o�����NQ���q���h�D��B��aKe��>���� ��|6��	B{�6{ �P*���;
hN�;+�RYzJTP�ȡ�
R�D; ����o���3qF�m��ӹ�H�'�Q�:d��N�q� �}!�����z279+����<&�)e��#��,�pe%*�o6�+!�;G���]�:�k���+�LI�nM�IN�vU��-%EJ2v�� �����t);!�g��-��k��D�$��.��VSIn�}%�t@�5��J> ��hrI�vfԗ��m�7 h������® =OJ�<��J���q���q�lH['���������򝗾Mxߏ�3��x�n�dvnN^x��ی��f�D6,0�ِ��$����G�� ��H Ӕ���T�{ڑt.��!>bcϞ¼�GDȩ$��L�%s~�xF�y>�ɋSpH����'�p��C���=��Aȴ���f��g��
�G� jd�4-��;V`I%SVb8���+i=&�6��Y!��-�hgM>H:�f2��e#���$�ȾE	m�HA��s�.�5��R�ը7$i���d�1I�[��<(�Ar[���uf6:J<���g%%}=����M风/<O�ʵu>�!`3N�x~}F#/>
I���xX�L0�B�4P�o+g�S^:���l���S�S2Y���;��\�eY�����uϰ��F2��U�=+$�`>�GB����̀�H���Əj��0b�2�P�)�5�=�zz�ބ���h2c�����������c�rQv!������S����c|�#G�{쐏fH"y_�'d>�ܙ]��H���p���'�V�?+,٢�{t<��[{�A�ɨt����v�g�<�c�X,e�T.65u"�n'�d�xo�1�w����� ���>� �υ���$�}E��dY.�f����ov�Yk�[�k��RV`�/�IKAۭ���䔥\����_�%`
`~�Z��"=�^g-� ��@�K�)d#na�?NHa�)"���,�~��>}Z6��$T��ZW�"�	��l���4�{��[���=S��T��a��₞�b>+i=N�:%�E��a�wmz���d��`"�IȂ���(P��:U��dqqI�z݆=���@g�d�g_	dT!� ����Cv��4I�1XÔ����sp[���v����	}Á�Zp�+Kd�� ��F9���A��+"�SS�}���>b��Ϯ��@���
�^�e���b֬Yݤ��@ikg��/�q�g�2��y���G��[	Fryu,�e\��c�t<�
�s�zBO;�%L��3Ȏ,+�=�pV�SY�m�c�ƐV���.z�|�
A�T�.��y�z9��� -�0�����e����E%�Y��9��[;7o��.�.�=pn<Yb	���0�w0b��	z��JBz��(��c�6��^��齞��g���Ɩ�{�A?�|)/��
��4���5���GR��eii^n޼F�_��_d�;<60�D�q�̆a|�Jt;#��E&%�z�k�0�s�>�q���KL�z<&�f?0~P���L:$�z��ގ���f�hr��������n���l�߈��(��&�����O0����}����>޶�F�b�Ǧ��4�Ԯ�o��v���vQ���,����w�Hx1,Av,%2�)f%�������>w������l�2ϟ6 �<�UB5��d���n��Yk���ի�eg�!}O�Ad�d�3m����įC�v�)�����{I���(q��	��c�2Y���c2�T���hؓR^ɵ�w`�9�cR�!���^6 ���~%Y-%u)%^���R*�p����������DM��� \���7���Dd9����G�^DeB���q$��#/�ȡ��(k��܎�>���x��)xy��T�y:z����8M�ooL���G��(�9�/��?	��>�	]�l�i�tpݾw��W���o��o��'|;! '��z+��:3��0|�I �I�F���QʟZ\�b
�K�(�����f��3h���ko������K[ؕ�٩�X&h���˩�gdO�����u�6Mڞy�I��P��6�0q�n�g��!�M�s9A������D�Y:��@D|'*�"�5�n�D`�?u%A(A�¹3g�gG�"5�V�u�VtL�Ig��BM鞉�IF��Z��)0�;4EH�PÏ�y�a�H�X�7�xK�x���^`�g!_a6��غ��F:K�YZ1'�<������m���ؕJ�.��ۛ<6\l�T�����j���%�3�� ��6	�qf�܃� ��h%mU��)H]�O�ۑ��4�-��nI{�&�QO�LLz0��}"���]*���B�2��V]FJ��l*ׅ(7)���;7o��.%}��wq�@��N�d��1���(���r�D0�+�Qm_v�{�{M2J 1��Jef'p\���<2E��1:��g
j�=�|*��L&��u���x�7�q��$��������q&�`G9�^����	ّ���<��J<;���U���
��Ͼ�'�z�&r��'��?�o�Oegg���o|�_��W�?��_�Z�&Ss�4@t�ht���ʲ����W�aS����'�<%�=�	�G1_<oI;�+�m$&���ݘ�bH��3�\㍃͘�Y%��BK�2��6<�s~�=�~8�gtl��)f@� �`��D��z�M��"�7�\Ɏ�h]*�D�R��4�:���HI����U�(%2#/,9��9�dl(����Z̔���R97 ���ݐ�w�ʍ7t^i)1�v�)m}�{��*y>�x�ڊ����w�n��7�1^k74�Ć��0�S"��F��ŵ� �=2�(J�P��+�}����1ɷ⍐F��aq(�K4`�3�{G�n�o���P��m����Gh�(�üol��x�����}����
B��T��~n|�\�����;�+��������P�*88���-l1�ኌ'V>�w�gk��n�\��$l\��M��������ױd��?Ο[��q��7����/����Ͽ���g;! '��zS@�з,;�2!x) ����Y?�n�Liw 2��eyz^�-���MK�?$�h�B�Q�JKW�P��k08ے%����j��ה�vC�wj2��(�m%:{2R��'��SYz�<K�`	{Xf��N��{H�`],�$��@? ,�YE�%HL6�&����`�C�z\ �> g
iS����irrB�g�轰��KþBy"�2����@D
���P9
����[>��-�l �tD���tY��������g�=I=ޜL(QCS��^��F��L@�@z�:����FX�^���J̢�� aG�=ʕ���� D��@Yk�G*^�������= l��`Җ>�S?�nu�}@rt�2�>�^�Mu�����;�啷ސ�nS�jOArL�{�%m�8��
����[��
��L������G?�=%
�\Z>���s_�Y���s�j�� ��Fu��	��DT
��&S��dܑ��g����W(�ǘ���mJ�+�ԅ~( } ���ʲ���,��XQ�������rJ�2�8]̓���mo���m�z_�8�Q��9}=Cp@z
lg�gi��45)��W���X�6M�z��e���@P��<�9����rYܻ'�J������c�����;���g���"��	��1nI��Ӳ֭+Y�e�ْk+w�O<�c�D/�=P�*f)�C�gc'i�^+F���zlY������)��q����1��־�������P%��>#6�#s4bT�A�����q������'��pج���ƚl�=Y�~CxF��4��dr�^�t�O}$~H�&�r��030���@�[ޗ;�ݐw�zM������ɶ�7b�stH#����Ũ2����=a������MȬ����B��:pi4�Ũ������=�(�1�l�+�S�߰�ܧ��Pvwwu�gEJ�	���!i$QL:�w1�N��(cP��H}�zs����k�U�"?���E�-�>����eL�e�=ܳ}��}�=fcF���GZ����<����������y�GztF$6�c��=
{?L��
	�X�̘��qٞC2����,�Pf$�Z�9zN�����VC�%��0�ld@��lfiy���V�O�d;! '��{��|.�
\׎'��p0�w�	(ځe|�F$�W`����jK��a���5�mD�u�=�� խ�:P`�k�T20������ܖ'�</+�y��7�_}�Yk}���P�i���}�jl����Ȭ���0�kz90��T�s�H%�8 �Va6��-��8z.(=P�o*h����ޮTQ�4��>=��i6i��k�/�� ������.6�j� �.�#���p%a�_D�
�.�� WZ��9�{fse���!�k"�h�G�
dt��Q�QY�8C�6_,�XplN�8Z�G��#��>����<��TKA�a1W����6?4�ؠ�{��Q�UO��6�)*�F_��R�g�OQft[	���ױz�ʈ���e���LN�|����r��y��}��g�}���v�T��׬%y�W7��e��!+cL�%���H��wh:�$���K����~������̜b��w�[��� ���/o�%S����&Ê#6��!	0��j�pH9�	%��L^�ۘo�z0���5��j:S��L����NeE�>���κ��3�X6��DbJ�@�8cA!���T��L3�O&�Nϴ�+2Q��~���?^�f�X2���}^e�R�ӤQ�B47?������"I=�AI	�������E���_��d�8��%��ٓ��3�e������{��z�L�ǩk� G�l`5���G�͙u��Y��P"! CC5��z����y)8Y
S� ���A7�����o]�V�UR�)��]*<�u��m�HZa;���b�B�w	ejfv@���^�}����djb^.�v�48�m���4�N�"	��l��ڊl>�#ׯ�%�oސk�J���sP��ǘ� ���ҕ�$��0�p�D0d��������	]�	�,SD�b�L�A��%�0��'E̔��@�W9�U�Y"ܧ����$K��ܣn~~��
=*���A���Y��G2�e?��~�ga6�+�%s��w��׶q���3fŎ�}TFu4�������g1�Hx�$؇���(+Q&a�o��<��1BWS{�'2v�������� +c2ǔ�&C9�32F��+�
�^�q�9��kcd�-
@L�ceY�D�$�c��9+s����+W>�^�c������Y�D:^(Y��=|c����`����	����fO�:1o:,c���-�]Ua��n�#+���3���y_ܼi%.������������%e7�N�ͣ�%�)��Z*�V��&�bj���!�h� �T�Q�QH�C�	�f��� ���� wV��%����P=*����y2
Z��Ӱω4	c2ԛc1�Nn�k�i�3�Pr(�y R& 2�h�����f�&迀諠Lh`j�{=��E�X��P�;P�c�4&�I+$>=��|�\�V>fiPZGIX��8�Z|?�Lऄ	� l<!9�1ƁN��xj<��H�M��@������q�
t��������'?�Y��f�K���Ұ�N�K.��ӧN)	���^[ x�A[�s���9y�U����~�f���-�#���h�����u8�����	:+�T��o^��2�{k��Y���)aI$G�Ե�ސֻz����@>����m�A00
J��N*����Y�+!A3���He$��J�ڔ7��)�dIN�-8�d��}�\��7��;�y;��[�D�cukCN�?+�ں�m�WJ,�:�p�*ZI6��ea�<����_�Hd��N�� 3�+0:~��������^πL��E�CQI�@���7ސ��	�Z��t!%����y�����[������ֆ���)�8� ٌ���p�� ��Gn(%l�o�@��rd,HZ���{clC�����N/�Jf��^	�c2���T�(/�鷍'F����
�Q�]؞�����L��SCx�Fb0�d�O�]Cfpn��$mi)���Kُ���m�Up����k�������(�s���@^{�eyp��ܽ�.�QWǑmC��#9�s'�pMFB���Ҽ��Xc�1��ærNIG8�3�m�h���Q�>5�C�B���#��b�2
h����dA0n��P򩜎�"3�v��zH���E�ǽ&��[}T_�C{�X��C�	����t��6���"UDB$�u8�;#y[�l��������rLf"" ����Ҵ�=�O̶���4���=LBL�Ɩ#�d����oz�CI��E�d0�$/���i�������򓽝����Y����cv����],|��p8��ݷQv��F��u,L�.��L\tZ��DjY��P"��B�NW_�!u�iH}�����tRn)�85����nC����Y���=J��,�{Ⓘ?�՝Mɔ��n+h`Jg���2k�D�������pD�Ϟ]��'�K�>�̸�i��X�cf ���ܹ���f�7@{QR%�Ʉ�>Ic��U����Y�m1j��ӿ!y:�V��b30�S	*ɸ6��!ew�l���PK&�"���qv	�AP�k2�q��A1���S4"��+/S	��k���c��D����B��H,���0*a�}	D��J�gr����YNSf� Qxn�[�)`3����u�V�����}P�����a�� ���-MI�ז��Y9{�,�Pd�¬��I��0��uIf`�6�����XC���j�;��O�S��,��,d��2;�$6w%_��T,-�d��myy��&q�2Y��x�lm���{
*+�zߺ��G=~�3�0�D�����uB�4����̜t��P=�\��Hh���Pyr�D�`��(U��%)��!!P�R��R��3SRR����75#�\� �
Y�t2FE8�ȹ:
���غJv��_go͑���{�R����9�d�U]�w^{MZۻ2tF��~��q[�۲���t���"��<i�������	�oU=��4���6J�\��ʡ��x(�7c���a���%�r�`�g:�赬����H/������96����'1��B]K�5QN�,�	�����8�TE:����)K�f.C�8��![�"���G?��a�)��=d�oܼ&��J�b$����no)��do��M�^A?V���${[�L-�� 3�o�CtI��,A����WY��0����%$J�2	����r6��\��`�A����h0vѳ�ϧ�ǹѥ:R��:���NO��jG�<�����f� ����'���'erb��x_�� �?h�0�GȀ�@���@6|�?�\�6 ܣ2aʣ�_
f�_�F�$��~X����y0�%H����HX�ՖC�{�0�p���cC Y��s���DL��{|<y�5?����|���p}�05�[��/	,�E���7��#J�J�w���f뺒Z\^>ɀ��v�}�7D�lŢ1W��w�
�����K�t"S��U�{��'�xVj�k�h���z��JmGz0�BI�gRi��25� kkk�e�b�)d%�dd��Z��F7��v���7)��.��1���	u����9��hsq�d�V�<�Ŵ�:n�"Ƭ�ׅ�թ�,�?B߆��G�c���s�����	�D��=|D�a��~���+��#ubԢ����Ԕ�v��@�
5��˦��CB￤ ���k�L��\,< C ~4�>D���v��S^X�c��- цc�%�-U,�<H����2*cPT��y��zt���k���#C4��u+�M/I{��<'\�r� �[;���V�E T�T(e{V�eQ`6駩x�,
?��p�k�ngeq�i�Oe	
�p�����/�x�	�:܁����E6� ��׫X,I�ἔ'&dnvQ
Jv���S���|_b����Yy��{
�-)��)PP}�lիR�b�����M�t�259��/'�l���hU�wKQ���@ġ��(�ͱ_E��\8���r�e�x��Y�����I�h�(�)+���g�w�V��Rp�R$d$P��R"3�����g�vl�v����Yj�(i�����Gy��kJz�-Y<u��zm��|;&���l�ǽ�b��̼����C�} }�3ق��J
�3r��]q���g23� ;U}n|�~0��R+2���c���Q��(f�9��3�%��w�>���ײ9蚞	S�t��!�(Ϸ���l6�>���D#�n\!z��{1PP��i�D>)��n�g0���4�}�2V��s��g�O\��{L~����[{{T��࿣�	���F/ʈ
X������(@���羯�6�����=9w��u*S���·��ܠ4~7��+7�yG���>g:�;]9��(��=٨�2�����^� vH@�R�bu��9�Yл���=:,e�#	a/�1�kT�b��4� �J�wfK\�\!�3ϊ�{dǺ �IW�	F�� Ed��c���%%���A�Y.�U�P�f���d<
��G�	�m�P����c���pz���� ��0}���[eC�3!����sC\LiSHb�i��q.�㯏��7%����9�Y�~����R��9�Q����렇d��d?cq�5zDj����3"�,��t�!�B�l��>���Ą��տ@�㹝�����������?~|���p�H&傊 ��A?�S ƈF���tBv��+��)�s� ��@5� � ψ$�AFJ�*�ܭVٜ�r������|��Y�hl+�{C�*Rm��`�&sP����d1Pv����~w(e,�ݶ��"T��v�L���iڡ�;��| �Ԡ���#O����X�h�S��2�:i�D��K 
�Ꝇq��/�?�*ʴ�*�| ��O�+p�$(ʦܘq��#���!A��=x�@>��,ij�y�o�% #�����a3jT��8��JPP���
�=p��2�Ȧ���4e[�Z����T�����^V��U��c�]6����M��(h)�\Z:ˊ�\9�늾d�:MMM�,�Q �E�.A��({^��SO>%]�jr��yokC!�7� �1a�1��M��dnaIArQ�=% ��$�����.���H2�E
��z�A ��� `�P椧��F�h'���	�1�5�;�Ƞ�w��E�v������iJQ#K���&�LA>��O�/f�{{5=nC
���3rvq��d m,Cǐ��]\%�.J��O
zm��"{V7�ew�.�޽+����ݎ,���������Ҳ,�/�'�{�u�� �}�L$ُ���c��n2r	:=�(�ܼ)�
���>;��	�#�Cٕ�ķ���=񀺒���@4*[���e=h���Lk�2���d����`�h��,:G�6�ɇ���`H�Kdv:u�dB8 b8�#c4�#ª϶G_�{�ߗ�������������=�Kh�Y�<��r��]��n3 Ӄ�2HP��{�����ޑ���33�J�\��~�u%�d�K�����o%�Y%���~ٴ�1r�^h��u��ǲᵘ�����iwp�L��3B����k�}w�;ay(�''TC����cY9^��r(�D�1X��(��P��I���~���T���_�S�EH��29^�dg����;�x�T,��C�E�Q �Y���}��G�=������$c�6��kk�<��a��� !>L����#"pPN����{5��"Ǝ�:;f=�y����l���iX7��"����8I��53F�F�f�q� h��z�A8�>��DL!�������}��ʯ��o|��?�� '�����_�T������.����ڡ������_����g̫Gt;�]�xב��3_����_�@a:j���W��_���tuw���r"60[>���{C��&fÔ-{
(��P���K^�?�ٕ��M6 ����R8���N_6��f�Èd���	��_�rE>��O��_EZV_23yi�;0e`��,�	�&���̈���z>k�}=N� ��g&:����6�g=.D�q�]CJ�ܻ'o����"?�fL�h���%�I2�b��P-���bP�s5D��Q@�{���} �U�9�F(�)!ҞI�L%NGX�ȓͤ���ɝ;�����|�9 v7t�f=�ޏa��&`��]��C�+��((Ή�����8ӳ�����Р��#��󘛛���HE��l�`�Ν;�n\?|'��ӥ����,�B�3@<"��mý
�$�*�����L�#q�FM��gzbV�z�
[e��'�^�-[o��ǧ���I��9�Y �@�3����R���;�W��'>��|Tp~ssl��LVh6�m���������E�Ic@	�uQL%�2]�P��m�:�@���>=}���g?#7o�'7��ֱ��k�ݤ�;zI0F;��ʩ�E�d��_��<p\<_:^@�3J��z��%)$2�5���S�tꌒ�!3�~ה$J%���L �|�U5zn �g��̹32;��R.��=���Ǥd%_(ɮ޳��w�{wߒ��?F"{JD��;Ro�%���D�6}?F,��3�������Z��Y�.�a	H��1�[�A"����03��a�@3�~t��.��x.��=�()ZY]!Y�óm�%F�oz+`F�Q2`�,����7���/����sHL	LHو�*��w�zK�J��k�m�n2&͑%�ڮ�6we8ۑ�Ύ얧%�� f��7J4cN[��	>��@1̣0\�ؤ� 2phڇdp���l^bŸO:�.KA�w�g�h8w��!�ƒ-%�	�������h*GVM����j�\J�Ⱦ7`!�����T�,)��tDGY��x��ŀ�$	��/J�0�"��60�����c%K�m�Q����u��Ʒ��n��q0y����#��H^6ڨ���C��"iG?�c��c��1"aT��cڲ�T�@@-��HN����{9�� ,�����Ͷ��>�Z����)G�=�^A�����<���κ�ڃ�M��@~B���g��򕯤���_�t����ٟ��������^].<�I�\,�r�
�Q����~jh��i���ؽd�؁)"��t
.p"X�[T�H�n�^_&&'���2`9	�|(A9�P҂ɥ���
n�\ 0��}�IFH+�����SҬ�|�,ՙ��z�ْ�.R�s6�7�������������綖Ig����G���U߶�R�5��r}%FXe�2f���/�JNO�Ӊ��s�a��M�d���bA��L?�M��$� ��׷H1W����#�kkR�̫��n� O_�z5�MI�4I�`"�xjI>��������,����F=*f��9�!*�R�nc �~FoP{n�D=�;#S�vFreE�g/�^�;&&*����c�ie1Z�0<�gH�/�J��c���`0��k�ԪV��w �x���4A4�:��T6|Cz�T�2nqe6h�U���O���B'rJ�b�����F�c�Ѩ�HA���a ��9�P~5��T���4��v��1���r�(�����>Jba�0�r��0��J�p��c��f�%|#�o47���C��2�o�
��_b?�����2TM��g����29!�׌�c�F�p9�ka�
�%	3:=�f�-}D�u|��%�IfjՆ$уӭS  ��4$�GA�d+�};��)��59}�,�R���a�^SPW�ɩ)�P:jjrNfgN1;��8[�2	�A���c�}(�*�����*P�?}N帬�������e;0�<���gB�DV.*Y�$q�ޒ[J�f���@� �����*�;{������$� ��GF&[Pbp>*�KrjjZ�{�)�~���ۑ%�ӳ�z=&����o*�KK�fZ�$k�R�{�ٟ�i���R1&�������r�Ί$u�[:sZ	\O6�9q��fT�B�c%�(ѩ�=�ʛPN3	���Z�&�^��&����K�\�<��n<�6Lu���	��j\�'k0���32�-�'����|�w���L�IK		��a���_�9���0`���&K�JJuCQ����Y�A���3�u~;S�o�&��X�<)].J�ѓo~�b�<��]8{N�3�td@�A��ό���01�Bt ��J����J����<J��:�t[�lً�1�	F�3h+���:�	(��9�!�B�����21U����D�Ì\�`�K�2� Q41f3���ק�*����%��
��A6�dX�!�u\s��Gy���.,�:�+r�>����̔	=
D�2�����<F9~;��(�e���(��%aѾM/�ä�!�#Q6�>d�G��?�[֡R&;�S@��+�>8��]�-���[&�s��$�^�oi���\��gm�5]S]+n9X{F�ь�쿑I�_�r��l֯��ًW.�Oӳ���L&*O?�7�女�P,9����u{��vWVV�R�L��ꢦ=��|�c�JHh>-�+l����`,f$*�2S��I#-؅�<�=�Q���r���(��Q�}/W.\��	�j �x݉�e���k5{yy��4-ʂ��F�G��=�C�b 7�T"=����D�L�9{��@4*�0���+FiI�E�0&�]`�EZǇ���k
ju���=,����>9Y�'MĒvq �R����X����@��t�:���=�8��@}�+���2iǕ��ޕ_x�Sv1؅<�ʣ\�sr�W�473��hOb�@r3I�A�ft�3�����mW2�ڮ���{ �N���0Ѕ`ły�W$ 1�����&b&>���Y��a�.���yDc����.;;��&�K o\cDs�Q�슂y�Ƞ'�&�dC�T,�C���c��S��%1��Pb��{�i�AJ$Bma�̉�7������S0j��L��NMLH�Zgԓ����N��q��)*��q�GJX)J�$������pejz^~�@�qIl"���R���g�}ɤ�iQ��C,��nܐ��/(I�쿣?�__S2�2~��B1G"577#��o��4ݦ��NU&de{� F�x�(�R�F�xԯ�|q@���m6W{t����q�����5N�$���)����;׮I�T1 <fJ�ғi�K��d�%1("��}�ņL�h s�!E	����jDur�z]un��/~���Mc8�Xа2n�/u\w��R��շ�W�W�����چ���A�Xf��G�LeZ���^M������á$�q�J���|2�ҥ��m�M<� ��W*Vr��I �JI�~�iYu�H��ʽ���%u.�8�����_����1��Ǖ�{���%��s>Q�1���>� ցe�B�����
�Q���t~��DUJ�b��upZ�L��PuQ�j��RX��M�����&��)m��|�����dD�2�^�8��0���������x}_�:����Y���E\�}��#-(��s����R�RSr��k(1I�c&��nt����ͼ�cjO�WH}�t�$M�%��t%+�RB�D��^��"��A߅^�^Qb<n "D& ��L3���@�S��%⦑��yfE�P(�ӄ�'#%C X�S�$���$є�x�#�c�c�tR,A���V��I&W�=r����9��oǕ���WE.���$4Q$?귰~� y�/�<m�x���xt�!���ԛ"�{B/�q�*���k�8��m���wt\�%{*l+�d���S����tQY�e���`�!"鉁p�����RƱk5�G�Qc|t�㛹&昣�ţ�-	?�	8Fq��9W�ɞ�e��zj4
�"��W����2��}�?�;��J�+��I%��z��֫�D�PH�˓
B�Ҩ7�f�����6��HBr�4"Ԭ3�R���C���@A�hX/ |;҅l���z)���5�U���xी�`�� e%�߹��] W�2�^g�O
09onn���h_�E� ��;����a$�F�R�8��m�d�@��, �tGF�3��j,L���� �������S��VP�d�e߱ C��}�O-x\[4>|�܋���o�GAAKH�m˽ں,e&%;��H�v���c;��)���T��JȰ���z }]om��V�*N%��IW�Âj��6� �тD��KI�D�=?Ң��J<,���#�~vvfN���L7���N7#�  ��IDAT�1=F�L�h6�+(�S�������� ��$h����A��9ZM.�h��C��Q�����iR����%�S%�B!�^����� �i�w�x�,�X�Dw�O��2�_��W}XQ��q���bB9
�	=�t�%g�z���v�jx����D�V(��0�9���5�?�S�'	������7���dNoՆ��۫w��:�y�[:J�f&*2}���*�� �������3����7�ުIUZ��D�m_�g��ҥ�	����UE��-��LKcgW�/O��
���9O+J���5u|��;zL�_ݒ�>��K�����Րy��>�\�����U����2����C����	6�߽s�}*x�1���3�ɋ�I��$�F�3f����^sG�P��������nT7(W}��+R]Y�ko�!7�x� �XD���+@0c*��LiZ����z�6�? ۘmH$zo�ߖk{�e�� ���9>��k\��� C�� �+�1��y}�����SC�a	�P&S�u�<b���aW��a�J��:�����&#�DC	S&m��j��L�fd:(*P��I����sr���H�Z)� �%��iv���o���B]��@�b�Ɓ�)�g/��AIQI�.�Q����Ʈ>�m��K:���+;m��P2��C�j�Օ�Z[��]�"�ɦo�`z��:fG}x���z��e&2Ҷ�H��D�N�(G��i/N��`���,���j��a�j��6�/���fI�דLYT��Ad��6�sdM��������\ca7�y��kJ�*����d�Fj�XIܨL�ᒢ��i�׎ۇH��������:n;�/�����=&���>����kQ�
��\�G�~�1�1~\Q6���N)|_�2^�)~�vs���v�q����Q�=X[�` �d��<J5��vXE`��,�a$&1��1����E�kZ�����a7���>����?w������턀�m��^1e{�`d�}�t;�D�l#ʥ�Tbrj���J6b$Ʌ��Qc���cCn���x2hB���n z�Fj�5�� 	j��IbFb��� ���T-l&&�G��QV������B�V��b�5@mL�c�c�x,O�"ݙ0��1�cM{����W�{�*:~���#���":6�91Ҡ�!r�e-S�Nz��㳗 �9����	'������4K�]� )^?LϢ�3`��3͊���A�����RrfbV�����=�;�+���[,��}J�
~��w�z&�Zw;�(�dC�G
;����Gm������b<6��Q�2�L�[�9c`v~�J37���#
{�1��IR��AR�M��������Ј�hlҀ� ��D�������t���~��.38q���7�c�]�ݕV/ES��7ߓg��ϧB�8�ʏP���6�8FlZ����sYJ���y:�א�@ ����X�Q{� �pP諫��{K�qJ1:J(����7�'�)���)�3�ll����ZXF�����)���>/�6d��#g�TTL��k��sX���ؐ/n��JMJ�,ϥ� go�;�	8�=������\����]���):U�~Gf�ͱ��eo�G�m�+!.���C���g΁]��Ҵx���ܶSY䒲^ݖ�Ɩi
��2l�tWCi�ayE<���iZWЊr"D�%�P�����_��,Ʋ��wz�{1�95�EV�E�E�8�l�-��l��0`�a���~Ї?,��ڰ �݃�6�n
m��ę,����2�*��Ȉ���Ý��:��x�U�ltU�b2##�w�瞳��k�Օ������%����y���ߌ��'�K�a�7��đ�yqF���*)썸Ơ
��4�"�Jx�D���*�8���ؐ��qi,��ʕK���(�Y�n��06������\�x� � :��g��J��vKgG@p������~
^�Ж��iYk3rbQ���,���F�J��A��ƺj�����5�onoȋo�(��-f@N���Z�O�w��o�Qr{������Ïcja��X�VX�Z5���?M��W.I[����M���%����?�Q�t����"]��?c�"�*��pWW�#t��agi��|w{�}j�ޮ̹5�EV��!E&<��>��#�s��Y�)�a�Aì��/�CY��RYfWķBV>R$FГQ��hkDa��{�Ҙ�4�#@�pHI��
AJ�Ӆ�T��R� ��P�xo�/�9��&������I��^@��
�#j�)� �H�L���|$��1I���$LF�J[W?&�[�)K� ��qW��4�ɿ�q�$ذ�@�����Dua�<�ՀoO~M��;~�vQaw��=��jU�y�w���#W��{Dp�΄������B��%��I�X��Z����̞ qؗ`0�s�H���}���?�񹧟����f� ����v��Do�{�U�+�O�����h��ibc��M0ot���d=��O���6b�EPg��|ʹ�4 �@�пaH�n3���e��Pi ����癆T�xp8��2N�e|V8�+�_w��4��n��&�@���@�����E#����H�"��53g�B.d	�Zs=�E+H�ȱ"����9z�I����PI��4�l�Ɔ��~`��<�5�_�i���c�g��:���׆���!hn]��¶�u+>Ru0���c\S��}	����ߖ��G��1PQ��
�BHij�s�bd��W��GJ
W
�R8"���-IQ#���ϊC���R-�����~? ??ϛC��~9�U(z�T�`�ڤNY�j���-��)���?Y-H]�A��������M*Uņ0A_���;�`
�쬓�$@��~���W`��A�g'����̔�>�*0U�����jO��
e'�񜪇��ɀA��M
�M�A\ �f�ijЎ�K��f�8P��M�M�4>��?�챣2=�����5�4�:~������>�}&��0M���/󋫬B�d�;��֨)��%��]$��;?�����Dz|�`�h4�~4��� �Z�g�]����V��/>//����+U�	��Sx��[o(Ю�m7�o�*�dI���^ψs�k���7�P�$ae �3�Q�}v����UP�
%@�^^��~��^-���A:�Ӂ���@�ʦ�G��JYƜ�U֐�����������S@��	��[��	�!F6P���ؾ�g�������\?ߖi�f��@R�&U#���QG��3����wQN�/���Ԓ�����WO�C+G��k����������qg�����0�{ҋ��ԩ����˵��\�%W>����O}T��s�h�e��b���r���pz;H��ӟ2TG�@�G[A���|���%�ܸ!�BYV�,˕` �>S

 �d�iL�(�2)Y�c�3����QR��VsS�3�P�t�J�1��16���^�Z�(Cu�-	u};~r����G0P�iP�
���g\z�X�`	$�t݂�7��>k�� �!!�]ˠ��v�Om� p����G����˵��洓Y%�}�A�g�X���d�����A�����#O���w�g��,��GEa�l0��WD�Y�y'�Ӳ�3��凉��cg����/3@�'��^��j69fV�H7~�I�WFwʝ���"��6JXy��΍�"Ҿ!���wTa2Q�t���$1ׅg�8�Ƙ7��N��s��f/���1H�[V?�B	���1���X�V.�A�Pz�������hO>`� �wt��^+��J�^^��;�K�����jP���>R�hJ�.g_b�1����3l�|�tC�F�3���>]6����$G�}`SAʬ�I<����LO~�4����0�f��p�=�̵r5!ln��J2:q�EYv &l��;L����ʁ��-D_�d�|�����4�YR$�_�ү��W5肁T��̢/e~��Q� D#�-�i�c�F�pZ7C{�H��5�Mz�7�	 6�q1���@gk�\���-U(0F�D��/==��^�ޠ�&]��׭`����k�9�6�6�l�iYr����_d�,#��ݭm�k��E��U�rX����8R}��gh+��L��ut�yf��V��lg!�{J�Vel��	 s��r��1�|^�ASH
�xV���w]�w5໮��Gu�T���� ��L�
�ν���8!�[��u��4���������a��?�%`�����o��+�%��tp�#��GPQ�Y����mqq�sY���\��.dE��R����:v�����������8��ò1ؓ��G�>)��RY�>%�^�4(C�j��=� ƽ���4��k�9�-]`���:���R��zTY Z��A|�A�����mJ��f�sG�{K��[�7eY��z�\��^�h00���Q��Sg���S�8N���H_�vI�-{�*�����^�ȑ�y��B*�!�F�R�lu���Y�Q�J56��:�u�W�IyeC�K`F��m]�vu��U0�T���g��ԏp=�AG~x�Mym��.3���y�t�AMC��.�SOʶ�#T�t}����Q�d� �Q�����x�\1��U�F��gyJ~�����4{s
��Ɨ��
`Job�v�8ř�6z���4Ԯ�=_=}J����_�嚂���Y<.���Hu���7B�$b�z�����=��)@v]j���|��S��e�ɿ���sP`�|L\�4k�3i�(�=u<��(�`!�.�뱐��������;�qq���^�A������FY����[�@�U���y5=?��Ti�=7��.��P��\�ԁֺԊ�
�M*,*U�C�`��T�o�J�K�}QQʽ�(;kz���M�B�I8ֳ�̎B��l��m0���^���ޯ掞ck�	���C�ss�S��PC�A*x��ի��4�u1����
琦�;�N�]�y7�rGv�>�o�^Sp2Y�������7tO�{�q5���r��4Ѡnz7L\�>��gv�bd����6Ak;Lsg�?�ʨo�����U��+rqL�5Q��U�:l\��fH�佗H���G�x���?��wtpE��γ7���ԉ^�k�?ntk�j��wގff4j�h��'C?M
^�~�dyeY7���FCf��ǀ�:�Q��:$d٨����L���mw����NqCA�"�KѶk���:�."0_C(%M6E�6:�*��E�[��� ���)�X {(�����t��ƿ un�2���$�@d���@9*�X۰1~ҏ,���|\f�8d��[�϶����W��XNb#dBf�H�
]H�g����$Бf<a#;S+4������ ŧز�SPBЎ�Vnh�'�� `�ga0���q���(#Ca� q�mxC�=!IZd3:��0���MݞYI/�S��3�l�k�7J�x��]@�-�Z:hC�
M�h�ǹǙ!�j�ҹ ��%}�\�`�@���<)�~�K�ϛ�81"�b�2�x`3��!�S�H��F���a��bC����X)in�:�/^j�p���Xӝ-1�H�E�@T�b��φ;;���Ч�l\}zʜ;*$��'��#T�`��t���ʣ>_���5��W_Z����FE`v~QΜ8��kQ�������[�.���7��ے�kJ�UG�3�^�R��?���$=4�#E;��k�Hk�7��? h�} ނQc���ɭ��,��`� �J]~��G>;��<����ͫ2�����kр�AʧӊTz���Q����)�-*0(ֹ.�K������7�dkԖ��g(gN��H�~��
ƽR���(0k��z�XG�lE��cA��t�a~O�����I�������`dFT,�vǼ^_�����N��3��iz�
�P)�BM*�Ym���{���b��	Y�����\@�R��=���v��R9�t\���O�csǤ���\X\S���I��^��6\c����ѣ��Y���0ؑ�=r�kz��.�*�Q����M"���
�gYe+Vx����>z��>�H���s�@�Sg���(�ӿ�_������z�s�8��P��,��F��9��� ���T���q�{%�r4���|�2� �����F��J�#*m(+��ػ��]�#*j8e$�I������(�H�`]=���"V�u��G��^2ʺ��FBU&��"�
㾄�Y4���a�w��
��h���
�&�{�{��UH�`���g���ha�%���w�w�@�����0���#S�}1��Z�p$�?�D����w4�~S�at0�,���;+�:҉jλ�i��Iխ��P���b � �#��@����7��`�TC�}3.�y�%W68�4HM"�а��q��c��}�zN�3�(���w|{��}� ��nʵǑ�UȤ[��xi�?�� ��9�g�z�n׽�J�^85���z�L��O=�,ܯݝ�f����T�^�z˅���Lsw�:'�o�S�����{RD`ڵ�e(���lL���(m��������e6�b����� AX�Za��P������4~��}��+����Ѹ����0��(
�l�\���!C�9ɨ,8��0�-��fy,�:�]���n����l�SbhS^�$����4m`m�M	h(�G�i�'$��\�^�8���k��d�Z�
N��j�&~p�!1�zZ�e���0�E ��L�g26�^�CYQC'�
ƃ@��~ԁ y&<����Ya굔���#�&=d9O?vD��fdk�%33�
nl�X	�L�z�o�� 
 �g��B.:�vs{W<㰎�*�7ɚ�a؈��b��-�8�!6~vz�������Ly\�T��ys[�1��-(���`D�5�bol"�b3n�E3z<'���g���v	�1+���B@�P�ZTT+�y*QxoTy򪛙m��`���[W�JeyI���������!�]�l��t�bPQ�����4n7�����5݄ѐ2l��~��sx��#H:W�����7"��)9Y����l�<-�e�}��G�e_�,|1����D�[�d��)�}��@�O�ټ$��W��l�����L�������_�myb�iPO>��$Y��ѐɲ��2O��Ӹ�6���l���#�v4T���7�b��*譁�SAv{-ޫ~�/u8������	�4<C��(H�.�{Wvk�Cc������Hلj4�'fG�!�9
:v:�	 @k�u�j�#��K�.G�b��t�����:i"����*��s�@Es���mK�j�;" i(U�����5
�z�QD��5���ΖM�W,Sp�mx�`�F�����=�i�g�e�2%���/�fڕW��e�J���1B�U�Pm-�뺊�G�~��+ �a�7�J�����lV�h��>)�T�G�P�;1��:WP�z>�6Pm�ф�� ��
�������{����9s��G�>�g5�3�م���^?�AcUږq!�2I&Ê5U(�Ax��������������v��)�ָOT�H��/L��'�I9{����������]��>&��R�1<4�x/ �߿�����VI9��;�'����nH�ӨqR�j��9������yF���m([�m� ��y��K�r�����+`ퟓ��qM�*2a�8H��9�|����0q��6a~.-./�?�1�G�G����h�}v<  �Wt���j��_H�J�v����,�:��[��~i�kH�j����/���<yZ�������I�s�۷(�ƹs� 7&�NO�?Ʀ��Or����GD.]�$O=�1�r������肦3�8ÌT��ꆂг��A�`R��z���F�R��0�x{�6ix4,./�uM�(�	�md� B�Z@�H�ׯ+`�9D �/�ؼ��5X����/�,�&[�1@&���B�tU����4�����e��v�]c7	"RD\�KV��e��\(��(�`,1��ɤ��5g���`���M7��"3��*eM�ӣp�PT����Q���RDL6	�6g4#@�>����T� �jj!�z���x:���=\�,-4�ɫ�gXY��9����K�^�*���ޢ�.�^�PO�Y����]�P+�����`�Zn����!@*k�W�Ue�s4���4�M�[��oC�4����y�̆fJ>�n[�o���8�e��ᢆ�H��@: M�X�w8G�`�b�	{Ob��c���������c�R��e��7F�� `��#�[r���ī�eckS�@���	i8b��C,��N�!�,"�a�g� ^�1=:<��b��s�V
� �� 1���;�</����~���* ��o�2�,s���s�����
���x�A�Ɣƅ�j :�1�=ؔ�/�!�aWFU#��}m���2�
h�Q��m���"��/��p�1H4��|+P�aKK����|���eK٠h���h!i��=S�����ߒ��V.o�K���WY ��������|E:'���}C�bejV�g��u���^H���`\�Z1u��ӏ���%�u�y��[[�&o�]nܸ��ﱕUy�������CO�鳏��hR6U��Y꣫ ����?w�����*Z����fj�Z���h��ʌ�X�R��Lqz��Q/��yy��O�g@j]��ſ����W�B����S�?��?S��:;@�J�#�G��"I��&��5�́�v�� �B����P�RP(PC�����n��I����jx��Jh�H$Z�뷌k;d�񬂶
6*A�Vǩ��eY�
T\��_���%y���{?�������y�� ���<X��RL�%V�Y��� �gUt/�^L�ϲN1�N�u�w���})���Y�&U���e_�!�i@7���WdЋ
Z��l�t��3��c���|�A�1Y)�����#h�� ��A�$����fw������̉���w,k��I$�ߝ�e{�~Q2�td�Ds��>I>ј��d%�Jsgsk\��{u%�4��e`�i8���`>�>���ի���.��j���[��|�� �o���
�����`)L��Tc=�o����;���A�W����
gϜ��}T*��+W/B!�~�G���M<V����0��޶$�h�LM �l�������/+�XO~���P�	t�[�/�n��~�~�)�e4���5�1b6�n�� �VtIAA�3'O���R�NǷ�ܼ*�]�#�G�������6ܱ��=��]�h��*�Y��F.0	*�t����<��G �n�J�q-�4�u��4
�!�.�ց%��k�R�]<��

�F���B�Z+��hqqL�~j�ը�/,=�R���Gh��l�25��|�@�
���"N��6^yXo(]�]Ȋ�ܻcz��3C����ۨilzl��DF��BAY�{�l'�d���^{�7A6X|�Ȳ��˱s��� �<Ә���g�b�kh	�Wc�(2�d�B��i=�2�ɠ?B�N¡/[�;��շ�T�$�&���N�m�[���u�,�c��vH-�������a[��-�-�c��s�P���v���Po�%?��^���� =�xm�
���21ѫS��i	�^')),�zA��Zm(��1�G�sq�Y��q�������q��̮�ʓ?�L\J�H��%��-�Qcc�[s.j0��KYT1exxhI���lƉ�A���C�n<�&�ҭ��w��S3+�R����4U��6����晃/B7����	y�P���pK�{�%�����m:�i
��sVQ ����Z��^��[��̸�8^V����+a0�\;����͟����UH'�f�%o�_�?��7�W��/X��A�k�D�`��Ԝ����.��S���|0%���dD6���ds�a��U�D�Y<������A� YnT)�c�]d����ϱ	(�=�������~�@�����շ���Ք%]G�f�b��-��U���U��2Y�AG�.�M�PfU Dl�*�g]oQ���!���� �����*�ei��u}��|K~���"�zC��˕�7蹱X�����S���� ��[+���-�-P�J�ڙ�`%AG�n`�q?�����x t�ӥ�O@�t=P���c�I���e�DD��[��Ҙ~�7st�$�aZ
�1T�P�`0�������JS^�ɫ�y�ga�Ϟ,��,���8j����~��"x(�t����}�&�c	���Z�y��YOff���U�LT�212"1��M��A^��{�QF&�弯q��d?(?\-�^�A a���R�L�&����
r��ϼ��
�|L~v����%o7�.������`[�B$��	Z��S΃}3�6��y�N︿y���˛�s����L���Ƈ��d}-��˅K���J�C�0�" ȃ���H_Z_��=��q;��d��ߋ#��Џ�4��Q Gm;9�&���޸P��GJ�J=q߹�V��۴_z�D7�(I-ͱ�y��v[�7��M~�3����^��o��E�b�^XZ���w���>��{۲���X;���3�f�@ɻۓ��׵�$	�����Sh�Z���cǢ[�֒V�Y��-�D�Ѯ�����l|?
���SY~	�߳]��8���w�;�.$~�|}H�ĲFx��[��\����;v!
�[IM&�E��4�s�Z��N��m���M��4xn9����L�#�q��z���uO_z����O~����Up�'|	x�G�.��8�cj�^\��\c�6
C9u*27��r��{3ƇM�Y�q�3�TRB����0N/��Fs+P<4�%�  �^\Y���C��� A_����Z/���Q����tݜkb��`I�=�QQH �3�0�����n�����ܹ��@ �TAB�;��lQ�2*h7������f�-/�uA�����8�AWQ���ecsC�w�oI��"��.�%}d�Ai�M���
$6����T��	�`����3䥒?���HTp �kTo̵c8Fz�f��5�ɪ��W�\7 �r��	���eT&K.�1��٤�G̈'ټ�Gq<��1ڟt@u U��g_���A�\ads1��_���Xt���~_��_�K)){��C�ۿ�R-Vz�;��>�T�L�H��(��&����[�7^���IT��[J)�HL*hE�S-8����o���^�SK�����>�����e��ˌ�γFb��?�HW��VwOn;T�����s��s��f�Ϳ�����9�|��S�˪:�!L6�;�ț<� 9_cb�)�����c��h��Q��T���twZRX�OC5���#�����RR`���'ý=�R�e��2{:�6ԪUt4؃�X�ǚ�^����S� ���79g��ڲLp������L��(:S� /�U�����) ~��3����dT���Y�P!$���
�3���I��%l�w�b�o�&{R�`L5���M�:t�����d��q��kѧ�P!$g ��^�=�'!��3����l�ޔ�<�}V\�K������*7&��W�Aطm��n�̈7"Ֆ�с^{9!0�gt=Ce��L�;_��@�ґT˞i�w�����c�ww�m���3��N|/�=�q�����~���ú(���xs���gd�����^���ƿ��`<����,fr�(;�H�9��y���;�9@3�u�n�5�sM�n�\�hL�SМ1(I��� ��*���I�f2�܍ӌr�l�~�Ȩ��=���s�s�y�!�|��FSթ�'θW߹lg�'�~� �o�`mxmmik���ƍ����K���T���;x<+��Z��<��jm�q"��3�N��xa��y�Qځ����ku�B��d� :`��eix3h P�m����[҇����>pJ�,����v-�/J���$�H7,����E!M�`�4�/������VO�����P���nC=�в�@�rD�L�w����oZVP�,E]�� x�ȹ�crf��Pak�d�+����u΋L1�թ;���]o�6l�E����E��(q`�i�CBd��RlS5����l�	[k\V^t-r3�ԉ�7��9e��$7k$]�l-)"�����O��ǀ=)hT��Aҟ���(���u�!Ш6Q�K��.^��ᦸ�
�ޠ�c�4"�C�H��6�?���D���G
vd��qVbB���q�ȸZ�bZ.y~P!s2�c���@��Aڵ۷����|�K_� =��~���uٺ�&m����{j~N��H�8�8�li6��֡�}eyE���h@Gr,F�f0P��^��^!a&���s#)"HGp�@�W+++�j�؇�����Kџ7��]�1��E�	���PQ�F�j�dks���Ua�3�;�}���>�H}jP��C՘_�*EJ�,Kg���Nx�R$�S�]���b�~��+��5�y�/I�q�FQ��W��d|�K�|��|���8D�|%�}���-�"��R/�HA��~���Uy��%I_2fb�?����.U���a��q�9W��

2�q��:#�ѿť�� bU��p=�<#R�\ҩ�����%��O�eh1C1U�\ֱ���+8`�uv����$�n����dZ�gײ�|b�VB��q��y��y�(�uܔү�33zm�|�T�3UTclY��6�N�e��%ɂ��d��M`�=�|�(�29Pӯ�.z!��[s�s��P>��_$}���f����C�2��84sх�T@�D��r��)7?g�!6f������*ڪ�ge?�e�?�.EJ��1&E�I�:zt�U�n�-�7�]�9��Ah��Xt#3m��lH��b� 	�7''���c*�{���{�Шɥ��VJ�hds+�X�_��8��F�Bl[��OɻU����;+y�}������������~�~}'��fy���� ���0>v፫O|�h0�m~Ƶ	�X9�)���q�^k�L*�R�ʫc�w�5�����a���s�s��{�yÌ�Ί�Ϧ8�{�䉭ǟx䅍�o��� ���H���^�桿��|���޶�Κ358�R�+l�h����j��rj�9bo�����5�bZ��d`=ˮ�e>=�WӽL��$q��Ѝ�r9x��{[jA����D��j��1jAb��r5FU#���#�6f����}(��N���?��a�AR!�(\h�j���.�H��',@ȸZ��I�(7sS�eB$6�ɲq��!�Q�/�
.�	��l�k2E�D����=(���X&��m�05"L)�ʃ#p�.?M��}�����l�����S��[�F����Xⲉ4.l�����]7n�ԭL��+� ��\�B�^sΨ�@3?�B�0p�U�mܒ�o�*O>��ܺqS��'%G��5��R��%�^�T���l�dogO�3�z�G�x\���r�F��H�a�X{K4FCf�)j@G��1�F�Z�N�-o�o3�@%
� �Q�u�����(0�en�~��25)�:M�J,���Tk0�qF5�TxC�Z	SЬ�=�؛�dK��
Jj�y�uL���)A+A�QVQ��HGN��Fi�sfh@�Sdvwo�)m�M4BC�8�R�AZZ`[6s�iT���[-��=�s�G��~c"c�AO����J]hzG,�q�ՠ4:���'6���pnb��gDwp���,x�d�JsS^����IQ�-O��q�wb��X��}�����IQF��2E%<��aO�AA��c��#/]9/{
&^����6��ѢZX�Rc���em=&��O��� �.(����*!����G�=Wx�b�J�8�Vj�JYr�P2��g�=*�YyCR4%���
�yy����K?�7�|SN?!�~6o�qM �?�#�@����@2I���ςI�
Q�Oa�s3�iZ�J���u+���	���.��R�O���>��
��g>!Eo�?Ǐ�m�o����e�҃�
�B�����;s�&��y�����nP��H�9���z  /A�b��f
@���wGc)z>�iFrxo'�JS��oB�7Ń�R�9��4!g���>H�َ�֧�^�\�k^�A�8�LT�0@��j�[㊆����=�Pt��51d&AG�}e�(�$o0�2�!z�$w������W^IʀH�/�SǼI<����V��H�p~�=�'���1�0)L2O�|,�s=x(x�F����K��������� ���x|��_͟�h��oɭ�����{x����{�O��ZC��J%�cR���֪�:#���4[d�L/�m�|Kk�qܓ��`eu��dm+�<g�Gn�bzX��H�yF5'M�M����>_kA#=T�2��LrA��W�[��UH���L�4�F�W�԰��O:��}R���.��9��&��E��f�R-��o��1�&i�4j�Ũt�T)�6Q�,Bd٘�_7A�@��c S�+�nHW�}��#C��4�@u'�K��c�Q���㲹�#�NWuG=��<��,�,���7�Y���a��AX�^�1����*�|�.���~9�)�����U| �0����!Y�jH���_^�V��M���o] ��܄�;��Xp��E)*�CoJ��Х���ب�;��a	 @Ԣ�{��E�T�H�O��j}?�G�d�@�+})��@�h��zZ[�k���K������x�&R)�葧�hQ/�43��?�@S4��>�ú��~%v,�pD��<��a��bS��<E��d�	��� �ޥ4�U�,)b�`�Y���$iu�����*�:.�����P�4&8�B,V�B�����K�g�^�����"�߈N������ӑQ?ೀ�Aٖ*Rz=�b�����������\���oT� �+eG:��P�1J�F��O�ధ��A!0pr�k��u�E`\@�"�ao����(��t��}X�n�)������1ϨwLJxOI�`����p-�^�|Lt.\��eX� ��*i�-��P���JV��I�g����OMV����:����ڕ3Ǐə�U9�r��?��&Wn��zh�a6J `�Д�(�ˍ1�ع��������P����!��x��u�.?��?��w��g�d�����;9�7������N�����&�Ɇ��0��=��N�� �0P�nJYw����5�*;�8�~��9��t��/�� ��Aa��Ŷ��!cw�1um����9�Fe����sC�ɟ��7/�)T	{脲���O^��U��l��=Q���<}���χ
����@U?p<  ���Q��T ��[7��4�#�(���3�qndT0L�A������l��'=#�)�55��4[��*��^��Ho�0�e)��э��!i02L�b6eW����J�Q��E���v�� r����@}8�����
8C��dK��d0�ܖ��U ;A� �����|�Ӂ����@i��Ab���Q+�,<�]�ۻrms�M�Q2����q���mmK�P���i�IdjfZ޹v]Z{mYY�diiEff����K�~�,,-(A>�4�0`E�јf`gU'8q//a0h�X2��R2բ'��IE�\j�cO����n�˱Cf�V�v�%K++�������٣�����`��`�R*�yz�ʠ�h0w���`���ͤtj4�j��U�jГRQ	s+ʲ� W'���8SR[��^�>�B@)
��,�4�4���.�-Tc2���a�l�����:yJ4@�
��ӳ�<�w._��۩t5���'�@��e�U��JI�ef��!`�4EdE=/��A�!@e�2.�AF�GGy�8���a����P�
�i�K-�׈P�E Yf�0�A#*I8/P{"=G8�SE�1U@p
�F
����@�{�'���^A*�%9�z�j|.�oF
�>�U��<�I��2���/��/ч�ȂS�5�r�#�n�K�1/��r' Y�U�ސix��^U@2/��9V ))�Kɫ��̀2(��~Wb�c�cX����� �J�髀�[{-=g]+������ćǬ{������,�aS�~*����<t�|��' ������:�)!e��x��<��,�C�5��B��X��T�Gt�+��@�[�uw��OE�������6���mV f)Ρ� M>n*���k<�;��1��^2���<Ε��w�����q���I9�������#�`�Ϳ�;�D8�g�S�>�zdy���_��%y�	�qb���j�؛��R��5�}0�N��p�(aL�S�<�s`|\CN����;~7�'(�{����{o�i��|�x @��#�C�F�\���;f��:�܎��R���m�P�@�̢0�A����	0k�X&\�䎱q��+�V~:nf?�~ȯ"�^*�۔��^������	']�~[R��em�Cw�fw�>Sl)�r}�A����#PS�t/�΃L{�?�|Z��q��~W�\�?��?֠�(�~�MC�7#P��~ǔ��$Wu�*�&��Ϙ�[���9����VoI��������zH���3�OI�ݓ���2�dg���T@��oG�;PTӀ����.�7��Mf���:Ơ����@��͂F��T��Τt��Ϥ��"ۉ��|���`S�}�h�cF 	 f齽q�� G�%����ه��uRC=����T<Q`B�<����H��XF��aeu���^8���+�K7�{[�G(���
"su�����uv���i �_P(��M��i)0�3������4�N3?�g++���#���^���-����}\�8��\�yCnooj ^�@z�P�B������TD�W�Z�����c��J�Ȑǜ��E�p8�@�!�IMP�����W���Є � 4z\ؤx!��
|S"/"M� �j�&�U���hE��A] <?
@@0��>�� ���^?�1����O;):��(�ͦ�;vWƁ{�}��b� V��Ǡ���k�Ȅ�r�}�wGϭ�cPe�:��K�g2k������ͫ�V,�\�� ����/�2{�,�͊�ɩ��s0&|.q���~A�T��E(�k��j�{�(��ֲ)ԯ0����e���@�рv*U�$�����;�ȧ���,,.ʣ�������iC%�@n��J�	�!�g����!�cN-a�K�A�����o�y z���� �����>�]�Y0��uH;s�@�K$kDώ���Y�24��?��#�������w����F��Ͻ�k�x]6�}��{��ĉ�r����a $��R��3����n�I���H���R
�l����ٷ����=:�L�s��`��;��i[ Ƚ���Ѷ����u��e���%(��u�N��Wy�7�}t<  ���1??cWK�`{Ћ�ĩ��5���J�� 	�Ďc��,�Ea�*��z�Lz4�d�V��Χ4e�e�6@_e.�	y�	)7��s�j���+ϢQ��2���`XL�{b���Ӯ�+NE.��؛p��;ȸ
N�������\dEt"6sI��2�/;1��&@-0���_��\_�IZ�@��ӧO���te��"m�ϔ�hH�o�O<��VW$���g~A��Z��v]���u�H䵋danN���غ�.L�G��-�2�T�YR�CC���}[{�Q�G�<sE$4&#S���T��Ӏ��j1H,����8!�������̞֧ټ�i�bJ�x��
�n�S�䋿�y왧��8/��+�&;�-o\nq�*���5p�� 	��5�c�X��e��*�u�Ӓ_��/��Ξ����Wn�Mߊ�o�*�|eOj���|Ef c)�9����oI�j���C#aKʠ�o�)c'4;����5@!��͛k���?'SՁ�_�*����岷�C?��cL�P��0� �
z5�EbL�-�Li>�eP������@=,�%��#̞�SF �,�~fv��/ �\J�*d����u�����٫�c�>dO� a�>��1���P���Cc�Y�ʓ^����ԭK�S��̩S2S��W��3XNe,sͦi���^[Ǽ�c�����@y) ���	�Y)��D:�â8��!)R�J��#�Z$��~^�L��2�ҧN��kk���;!��J��
k���Z+�1�񁀙Uk��AnUBb��͚d��S��%�u���M�x�F�te�-
Ź�W��s�8_ɥ�Aa�]�W8·:���܏�1]W��()��t��D��}��Ql"y���� �f�2����,{M�z�64�O�U�d�/S^M����L�����iG�;���4
I�t����}�3��<4��!a^	�Ӭ��>�c^��ߖ�"k� �����$�W�C����~�]�\�d�M8�O��$�8��I�Pu�U܀���U� a�%����s9-�zy��7jZ��A `�]�d�ʵ_����nN�r������Y��nLh�8��� [�T"�l~� ���>���6����N2],���m�`|�;L"�b���hJ�I�0+F	?d@�(�18����$䃃΀f��q��Ar.���q���.�6DxM�k��+��&(gu8J���`�8${�i���3v�B\� ��dK)�H�d-x�1�w;k��L&���hu��~��dS7�o|���K?�/��"v�*?���t圌4��] ��>�7ʎ�X��������}DV����K?�s��*=�]d�����}��+J���F]�����`�TS4f�S�~Ve(U��rThN1e�`��2͓�P���u>��`�h�q��}�n�l�g5� 6V?�\-��������§��ŷ�����I�)�/�h���P�?ST��e�׶��;w~��xxT۾���6�k:� ,TI��F]f���Vҹ!l�E��hK����W���W݈C�2U3�W��d.�|�{p��v[
@PQ:s�4`B�W���1��?�xDZ;-�R��#�d@���+8���ffd��n��l���x��^t0�R�M��;Հ�����^�Ko�%M�Q��N��y
�
$�G��h�dw���2V��
G��k���o3�=\(p'*6Ҳ�,қ`N	P�d�K2h6�r��uy��qY�V`��2�X����1��lJ�VJ��K�l�\ѱQ ����D� M��<�1�B�
T�=gL�_�$�O���א����33���g� �O�V rS�����ƭ5�}6c#����Aʞ��[�Λ��;�4�,8(�P��9�Z��X]Z�+o^0��A��'�z�Jz?b#!� T���P�9�_9�����yA�5�v��+V�{�����9y���_�5(����?��ou�L��
-=F���"$(2�p�9�/�� P���G�y�-]���t�Ap�9���v&FZݨ޼yKZC��%
U`�b-Ii����3�	���=��j�fCb$ys����9r�{U;&��IJfN��<����������Vc�t)������L�=I��?���
�6�溓�������x�
�� �	Qَ-w���.�$9���ڕ�?��9�^�^?��[���8�	��xA�\@�AװBd�(X����}{W���]��b����I�P� 9��n/�|Ć�e�L��ehT��BCiI"c��1n,���.����V$YJ,��(e�`��qƥ8'��ʌR��>�GŔ/�����Գuc�JT������C}�<0H�Q@d�� UlJ�љ�,�%��w��e�Z���f�5t*]����ciе�M���{?,H�B�#W����[q��� ��i��5��e�R�z�"�-�������L���C#��@�NEa�@���A�0h-��� b��"_	f�����{|�Q� �����ړ^#�tDJ%d��hY����N٥�6���=�H���;��u�G��4���Ԫ�6veΩ�����5���hl�	�+�L]^�3�N�*�ҏ_�����Y�Ԩi�{�U*�J��SG%-e��� p�k*{��|�m�`],<�+�����x��bЈ�������� .LBkuq����My�ɼ����%�e_�9�K�ł���SG�
z
z�tK������#6��5@O�yA������aJݹr�A#�+7� ����A�B;:��߉������N2���F"��&�	�%4���QiHI�k�j��!�(I��~� �T!�.���=3;���Oi:�*��o�3���Ա�e�ښ�Ӕ<rV_�`�>� C���;�r���
��x���C'f�+еb0�e89�+
~��Z�\T��$�6nJ�}����mn0�]�G��){
�|�mJ�"������5�i���̌���{<\�����{��g(>U��9#'O�%�/��n��F�^d�nFi8q3�G�}$`��Ѓ*�~*��{c�F��D�2xVvwvduq^�zEfumy����ƥ+�Z`&OLo(�Jeg�������S�?�RP���"��UR��PY̓n�yE&�C"���}�ӓF�"!�(܂��wl�o�yvH^7+��� l�{ ��oh��M��,h���)W���;Ҽ�w�U��÷"S²�����IFC�t����7!r �vV%#��{~��)O�R�f��UI�,$�QKc�.{-E2&�@��5 �5����8"�xy?K�3����S2 ��	��~=W���|� ���>~�!��}�y���,��=&�.ia���2�VHM#$) c��C.x1+"1�ZB*�P�(ېB#�"��䋙'	�fk���$̏�&i�g�!�u�� ����R�u6;ep����� \�zQt�6MyO}�)ټ�.a(���S253+��Ǥ��łI�/���{����.�ک�\�tI���yX�}��T�A�:RIA� <p��`��y-�3k�`��ۋ���F.ݝA�����,NY�F?5�A��]#]	F�4��H~�#��^��ݮ|�>/?��O�љ��Uc*�׆�����)�f�AG�h6<T��Uni�
�/|\P�T�@�c圾.u<ggg���GdauQ�*x��qyx���9vF>��������� =*}�I�M�<��#�L=�pT�]�$;���F����ݎ,������v(�#���H�Q�MM�7�d��+bv����4��N{�7�q�:���@�%�����Nk ���@��W��>��̗g�2T��5�#aQ*Q�
8�RE#�r�AIQ�7��ގ�������-�ҹiբ)7���̪��)��NI�%�������T��J�D@�|@�H�AKǏν,ooޔ~1�%�<Y}A�zZU0��,�z#�y�2T���2�>�2�gl�xM��
RL�\��T����+�}�z�4Gy{����?%˫XC�2��
H6���s��
2Z�s�v�`A�y8B%�� |$�꜂�HVN�5�B�A�����@�x����C��x��ST\���sfN�rUJ?�����T_���.��|Tc!����߱�yaE��>�4в�^�"'�3����(m����.U��߁�,ȥ��3'�ڻ�l�*�!���ɠQ @M��0��r�|�ߑ/��*�A ��ϱ���W��*@\cL8�t��Eۘ�f�f�ϱ���P���^����	͠rB>�7��ޮ�O]�������K�� ��> ��xw��T��s��n�_{�}&�-���}���~5QQy�#�x�b(}�\�}����{�I9�e��2�>�𚞬�UA  �4���+-`#�Y���  �"��<���bg������[s�5SJ]��3g��x<  ���ǩeS.ֲ�(��%tSy�����(�m�$�D��Q�¦��{�qa>���~M����P�A�A���TM��gV)1N�C�(�˾�x� ���m}�R�5�\� ��9vJ*
$b;K��hP����&����S��/|Z�����dP��O��4������LJ�BNTߣ�ے�����x�V��o�6�
u�7�^4��LE���IT�/R�{�@� #	���`Ӂ�wI���2,\�QI
�$h4�bS�@:� ������F?T|P�B�8����ߪ�>{F��o��8.kpo�TF_�@�����Z�{�' {�\G�)+����~?� ��P�j5[Ҙ�J��0�t}�Aw�s��g>/{����~�����v������� .�}�B��؄0����*�U\˓�{�i9�v孴)��s��2��4��G#�E�Y���ػ�!�Kb<0�  rKb:l'���Pg�M�!x��~��K�����tJB�+�,�����\eZ�#�����@�e�U�_{�M.�g,�o��-ϝI~r�%�5�rb���/����>"
GX�1=N)���|�6�e�i4�wX`up��rnU��_}M�o_�y��8�&�>_PM;r��Tku�;ZQ��i"FG;&��-��2�ts��;2{Ғ�#�]�Ԫ��F�S�~�����*T�7���X�,ך����6�w5���>7e�ew��̩��!�o�;8 �輨����k2��tz�!7���
57mzAG�=qF�N$k�]ix�l����}�M�(S������ܤ�B�RV��� tQ���� �@P��L<� ���i�n�!Ejt��QiF��3шTN�@avi���``�� ,m���L`�&pJ���tH���o]�_��/L�}�!���!��:����c ���n�Me��ʨ��B�J��1�l!sG�!(�@4���({�(#i���Q�.�Y𹿇`M��� r�������q�����y��aǤ���>5�a����ۻ����c�����
�����M���N��e�G��,ӓ���I_1@i,�Fu~e$��Un�hg��w�����ț��<׬"�$�Ϧ�E|Z�ەۗn��x @��#��862�n������}I
�ze�ӌ2�d�WQV�Ep��xt�n�"�?��=A�=���~�~b��l(A�Pc2Y�8��g��琥Di�}zA9���wu��*�K$(K2��.]$h���5=���ۯk�DM��$�Ǝ�$�zq;qT�z�#4�h õ'>��lip��iQ
�������x�%�G��1����,/�E�����DL@ahT�[ "4�[�̍2Qʅ?�Q`�&������YAP�կ�_/��R��p��@�gJ��r��P��ڶ��>.����ѣՒN�a`Cz�m�y[���{���˗��ʱ��r~k߸�?t������ 7�<�$s�����	����,��i���#ȨC���էei����=�4ؓ=CFT2
�<�!���ޅ��(0���l�g%1�4iF�)1����m2�P�B� ��j�m��CK����yD��((��W�N�퐙�Y�{	�s�b
� �\}B��ݮT��f���R�\G�
~)�3/�%���(=�5�ynܠ	�[Q�Z>+s���O��g���5�C�d���-�o�V�J�����e1�i ��!<�<X\�k��@e�P�K�
d�(�'"�~��%�i}ڐ��BV�l�(�u��d���(X��ҨѫLi|K�q�����bQ���������ʦ>ϐ�ѧ%<=�s�W��pϨ8���i��jC�4�������j�DJooG�"�y� �U��T!�Lo#<��"��^y�E�uTП隖 �u�z�T��������Y�
R��b�ީ��Pb�(��T�B�lg}H� hV��R��ī�e��$Iő�����J�̦p��[���9��z�d�kjl���Ϣ���V��+}J��Ò�i�gY* ��)\�
��T�����Z����c�yw ��t�� %���`.N��N*&M�˚��k�}�> d�Y����4k�&Mx�e���$����{�|��8J�+�wz|��|��`�`��r@�.
���n��ν7��u���lii"cu��繄��]c�
��J��x @�룳�a�? �����6y�̒���/6�4Tf*�\��,a�'aw U8+5�9�zT��=�рN�������6�D�z�G,���ه�Lu�fɟ����"h��-�R�����S$E�Z/ˑ�IU�_P�A]j,,j���|����	{C���V��g  ���c��H6w����c��⟗�}�c�ors.�:����/p���?^�o�k�4@4^
�#��!��I���Ǥ^f�PJ�5Ҵ�JC����@���m�e!8а�Z���=*$i�83S�g>������f�L%>{8��IA�J@)3�K��A�����`�ֈd����N�+;;M���+��+�;z�8)b 8%g�:L��0�HP��,z��l
\�)"��Ѡ,����'4Wл��3�DR�s�_�S�
`%�����;��sEF��PU�ŊO������� ����Nr�<���z����3��E9;�"3��7��~>)���7�?��x��zA��՚ߏ(!�N�P��ӓ�λ��ՋV5�N�Z
���k���d�ZX�V���777g�͢!���Z��KN]��s���{�MXM�Zvw�t|]qJEr������NZ���c�U��v��M`Z.UdjzA�N_�zϋ�s�u?t��<�ćdnjZ�a$�V�I����έ]���t����U�SwLC���+p{�VH�"�'V䚮ͷߖ�^g�����+���PtB�=��@�:Ǧ�5�:V�<]CT�t��	y�u�a�O���z̰�'����>6����1{�*3U��ݡ�7S�Q�h���PϮ,L ���BEO�M�)�v���ǂ���q�,ܷ�� O0 ��+L T���T���yJ^�~Q�֮ɹ�/�������T0Y�����Z�b�³��L>�Yaf��Ǡ`!�Eoo{�
�?��\.[|1'���x:��Bm�'`[f�%y/�ݴ�\�Ng�%vY䵲���5R�&��^��6�����QM�ỽ���������m�7�du�������&iO��r*��P�Ȭ4P����*t�{�b�q���v9e�|���˳\J~N	{*��컺�ث�DBb��81戨���[�Zf�� ȃ�}}A�*����l��R6k��k�������ɜ�8�������7���u#�RQ0S)�tX���R�uQ ��RE�@��V)�`�5�?��-���1��=d�=��נA!��VyЊ�,�H�*3X:z��;uF��>���fWv[Y-G���2���/3���f_���x��4��i0Ӈ�l��n[��=.��zUJܽG�~@�3H�96�􈤱�8�J��3՝���af�� 	���ba_�.�P���@�~�����i�����ˤY������r�ş���|u��r��I�v�A �C/�����Y���Ɲ{u���aTc,� 5��E��Ӄ��^gW�Ͷ�i�;�0;��bo�z�Z[��	(K#�l>�<k%�}'��d]�4\��܆S�M�o������P��ј��<��O���Ny&�N�_zN؆�b6W�{s��)*s]|�"G��o�ܳu�s�.�A�gن����P}8��:\ͽ6�.�}�
J�\{���ӐƇ/��z�3�GGOe��e�=�$��+��3�mey���L�`�A�	�E� �+���#�o�����E��n($Qd,�KIK���`���i3m��۴/�s��s_VeUW�v��4�o�讪������s~�;o�z6}#m�`�1䔤 BBuk}KVWפ����ޏ�%����H��3�e��|��ɔ�rggS?��S�0mSJ��D�#�G r�M�>�c�t���$�W�",%�9������t+�ǉ��
X�`+�:�%U4�/n�)��$SPb���1��{F.�עd��{��!8����Ҕ�ŗ_���(a-*�7�)�u$j�Y*��z.W�r[�p��,zZ8�ԧ
9)T�RR���;�����<��9FE(@I���dM��8�JJ�a�J\bP�2�vZ���tu��s�F��A��7ҽ��u�?0.������@1͕l� QV��<JN@�T�꺡|�G�@鶎g)S������Ք�҆�i��<�ẘ2�����(�dy����c��p�lc^��m��8�׉�ޫZ5�����#�`����<!+w��Ǐ{�{d���n"���r�GdW�cJ��q9TV5���������v�u>X�4�z�w�"���G�F��g:{>��,T��|7�W�́k�)�z������}?���{�|���Ҫ�Ϣ�y?�	���=}�A�D7x;���U�)�U�0�2��e�����z��?��HouW��]�Z})[ݼL�t��ߖ|�*�AN ���7-�u�u�b�R��M� D��s0x1 ���:�ڶ��B��M�hu��dPKn�+��2��������@._yF�U����.ǒ��l^o�l`^(�@�MJ�@�S���0 ��}�VD��A��:}E>!�M�Ҁr�FZp���dX���Q]�5�,��dL���&j	 �ƚ�5.�5����@D����,��Җ͵M��F;���X�ʅ���M)e8�+�G� H�b�xC8�o�r�'�ϔ=���A#-���P�49�	�"ߋˋ�Atwym��~��#��`�5��TP�L�(�c�U����(Պ��t!#���Eo�ēE����k)��xK�c���%3�P��P�Nf%�Sb��3frp�yZ^\w|�Y��N���'����2�q��k��K��<�����Kt���
h�q�������I���I9v��}O�����L.�2�WE����4�V[�3�u���A�jnnA�@ַ֥�%Z�zO&&jcxD 80Pk+�M�-�.�Kuδ!Kk�$��<�轳�kd�XBY4F��:^�>��y���xyB��<�>��L�34�9��� $� ��]%CJ���>C�
���\<wE����h�5�Ю7�d��I�;�Ή@�
�s�~�&����k�l*u�}�7h�GD@�[lrW��s86=#5=�1,�.��J�_|�UF{K�\۾K#@���٦�}*��珧כ�s�?N�bFb��elrLl}�6�W�7�)������gB�k�t-��g�tN@lB��P 	��S&8���"(�U)��g�T+�|�%�(��3�>�tFɺ��"(�hGJ���Ĩ\e�72J`Q��~������A�t/(�Q	k�޼@�J
�y�?���y6P�HŻ-�*���2�������P��${�$�܎CU(��DQp��v�x�`��e�d�%j��BJ<��}&Cլ����h�?�L��0|��������0>H���r����a"���D�lX�5�}aƆe�6K##����' �'))3f�I�|�k�&1G����1�;�$1Q�(�~�0"���b��3�<#����+��1y|���f�+�\Qv�}�J3��Fe[����Z_I@[l\��+f��f��(�X�T�H���X*/[!��;JI67F�@7S��3ܭӺ�uL#-iNxq��� �N��F�>���>J��%�8���4�B:�p�s��8rm�e�$Ջd�<F	ʹ~�R�0Ҋ?���ﳤhyeM	T�&�R�1�wza�*U�."b��L=5�g�6����25u����$"���|㱀5�wDo-	'O��3���so�,>\�Q����@ |�.��e��C
�(%A�X��z.(�������]�p!k1̒���\{�M���*�H8�>T��D�3���9���Ң�D`R��r�������׮����)Y^^��;q\�ggdu}SV��%Έԕh�;;��k/д�@izbZ�?%�J@f�'���>P`���ɒ&c�ؕ���ɶ�g�&�y���� � ��L�5*<��9�%L��h�|]ڀ{z�&�aT��^���5����2�VЕ��1%#y'G���+���7^�M�'��-��� �t�z�:��^��􂬬�HFIEVA0����+�괔� ��i�G T���~,tW�D#���R�T�~�� �#+�դ_�b�e��1ɤq��>?�ܧ�ϘӭS�����eT�7$�M&[�gR�Yޘʱ�%0��UP|�JNO�W���?��
�u��s�C��(K�MhhH6�h:WR�\�6[)�0�ݖ�x�u��_�-�0��{���~E�=���,�Q�eGM6u!���|��l w��A�� (��z�9�ڭkb+��z���z�S3=9)�Ҷ�&��\]��UJ�B>� ����������Q�֕'�^�_��/ȿ~�_Jw�-Qk A]�ʮ'���7��=���Fpd.Y>&�C:_������섌O�$��������y(�D�
MQq�)m�����q��q�X��@d�n�k.X��3yĈ�&����� _2I����K��mˮ�����w��R��p���%B{-��2%�݃����Ɂ߉6�?�{��h� :t-%w�D�يw�؆x%Jsqx4��pO���c��#�g�X�M9|]l��½�2F�������a��䄉3��r٧��spGu<��bc�(��� B���Z�q[އ�c��xo �aDg^Ԫ�ձ@�8R�cc����NՏ��Ӗ�궔t�L��i��x�"�8-�TA>�������������oISA�diBA�%�X7��l��ŇʌO���J.���^�5Ǧ��,ĉ��1 C��O0?�ͺߣ!����cM�z�k�J�S�%��l7�S'N�����	QA6i�f�Q@5�����jMN�<-�b�(��&B�e߂!ge�=�(47����q� b"�V�I�2�:�Q��%� �:b�8UN"}CV}����o!2�@BΜ9'�N��/���_���$e5n*w��e�e)����8�B������7��VH.8�(����V ����;YZZbumsCR���s�W`�ݗ��m�.�cr��M���,�LMǤR*���7���])*P����ʸLVǥ� ���rz��K�����o�\�I_|������È�L��c��^ĔjO6�g�{��%�3�q>q�՛�uG��(X�+IE�������@V����m�nn��,���,�땔!C�r��Q�/(�F��粯
��V�u����Bt0����3=�1���ݼ+e��enІ�dW��y�S�d@D� 
9峟��\��?����߁L���bc����W�V� �xg�����(9��sߒsǎ�|z��������<T���h[9(E��zo��g�9��h�R�������C���?�I��S�Y���%�n��@%n��^���)�b��Z��=�fR��d�?����@�J�t���@�}#~+����}�i���slG�e����Ά �Y����7^�/~���_��[������"�]�tt�[��Q$.@���Us9�lS��JoH_"4��VSF�`�N��><E��ҷ�#t>�Yd��L/`(�˻J��̶bm��۟#���JX$��y� C��c���=�_D�(Ǧ�R�ɺ��a�1�̤��г�����mh�C#NT�L��'F�}��{}:x�
[�DD�:���$�M�5y�#T��H�n�ј>h�c(*bH��ug���G4����Ɏ<x�>1s����D�/>Z�8:�Z��>f�,�Qf����(�"�T�D�;������=p<& ���������0��0�V���pe�*6�Mq`:%.d(�]�v�U�Q̺r�X���T2U��<9F�rS�Uu�<�ed�¥2rN���oE���7e�[�N���YCZ6#������S��9N�9��y0��}�z�e8⤟ W,�l��v���e�*�X���8���;r��q�k @�u��2=�S�=A��F��
Z��hT�M9����8*ʈ�.2M�R�0V�Y��@ �d	R� ���0��7L�?�a�P>�7��}�H���"H�)�X�d��j*P5�����c��M���^}UΞ9#�ژlllP��)+$9hO96�*)���+W�,I���O�x��nq�AE���[�duu���Ч��x�,��V�-/_�kK�dr~V�5PF�gI�!�_33	�!qQv3>��T�m�&O�9�km)�����<%�Y~S�JAz�Qo��s"L��{2����˘�7U�8)f��2i4FO^p��-:�w[��}oP2�r�a(���s��09��Z���E�;)9ql��h�FV�bU���<OzQ�dK̆��*XC��~,l���~~���כ��\��Ɇ:�J)�T�B�!�lC�O`)i'cKMI���%5d`t��\��E ���;TԐ��P�%�}�Z���养��_���ɯ}���䂔m���)�����Hb��\)|J�|b|Z������XY2�-iy�|������e����z��A��c�H�W��F�����ȿŬ��箽"/ݸ&cs3��gǏ����f�N�Jd-r��s�f�����4�X�#�����S?�)Y[YQ������;�K��Րp�#Q} E__���qH�l��Bu��@�����XI�.��TH�PY�9V˙~-�?86�}0�z���)!D���7����V?����Jn�](g��{54����1��+�(P�j� �87W��b^"����P�{���u��L,�5�8�8Ra*N�Ψ��h0>�9���%@��������G�b�I���~��j�Q�Q��3��C��Q�hf䑥l{},&�a[V��a2:CWr۲��GH ���=TC��}(�1���޽��l��H|`��<\�y3*����D�?������c��xO��m��t���7�=X'�y��K$Y�#�v�'eߑ����IU��rMfK���s�Q���e�zR.�8+�_`4�ѴJN*�JR>�yf.����H�JW7�0��*P2 u% ��8�!G� %^��;E�,7] t(��B�h? I������`��uAy
/ss҃&��*b�S_��Xnd�*� ������8��R
8�E9���L7���Y#MlIF�P֠i�Q�P�=dɋGU#�YI�A0��a0�6�%qh�c�^��kCO 6�����6�� J��^Wv)(1k)I�Dd�Q�D	�L�ؿ�T���ni�(���Xc��(!�G��N۲��K�q��Y��2���i�D]�w[��8�I�T(�5�����R�di^�3�{/޺&��7���u�(�k6vi�HSi�O%��o��b��	X�t���3�o�򏽲��D$�(9j4v����dD�Ũ��%���.α�Ť�ޓ���M�\�HQ�4dcY.����Д�Q�2��m'�2��u,�x��`lܔ�:�w�m3�I��t20e��D�z%S^�r�H

R�\~B�ުλ�;��	uΡ\RD3��ͨ�Ō�6�,u��^��T,/�{K����W~�?�'�����A�������H N i%��D�(�doP���{�kr��)}��V �����������t�&��'�c|���	h�m}n'�\�:�����P;����r�����|W��[d�9<s�)9s�<qbM����{��ܡh�d�̌��7�����������JY޾u��>0(ХtLz�m�v�g�\����B�I	SV�d�inh�M��C��q�+d�a�z
�ut�I#�Q�p���<���}8P��d�a�U�#��� �Pr�ɵ�#�fb�9O=դ��(�u�g��(�if4��&�@�� 4OQ:�g���ղ�2�������|5<�k����F�YJ���D�k���v�$:r�U��zc�����Xֻ���ǈ�3�M��Q
W���?;����x��P�`����^")��k�;Ǒ�Q��Q�oX�w�� ��B�N��=���������v�z�b�8pl��v�f���A%-�����`ԗ �nȵtQfu�-eb����J2U�K�-���M���"c���^ZAʻ��۵l���c'��;���k��\�|ZI@6/;��hF����Y�� ���F�Yw��I0�XiF�Q2 4�	�O�^�t^AG햼��+�����ٔ��������s/|OIL�!�N�b�J;P"��Z�r��&ՌTH@���94����Gp<�	`P��w�r{]�w��ifDPz�P�/ 8�v]��6���H�n#�M�eQ�Z ��?0�34ʰЌ�ht�\$�����)ol�w��4)egiOQm+I�#"�-(���g�){A%��d D�riB�J�*�^�䢥��V�_W�鋧�3O?�w^���uk]jSc�(iR3��O�������-[%ZȦt{r�ؼ�ڞ�7�d��˲|+��ֲ���Ih$�I>�J.f.#rN�e'fYI4(1&C#��������8H6���c��,UKR�L�w&��_�-���SC�}_aO�Ѫ6��vh���:bJ�#�/�7F��W��R7�a-?23^lJ��Y�H��)PGvr��`/	�R�LMH��J6jJ�U���Kҭ7L�>$I_YW6$�����;�7ձ�N�I�c~��*����_ea|Z��6C�)$m��+}^��=>7#-�\�}��ɀ����Z,�	ٝDO���~�������?��������\��V���@HH0��a�X�g=H3s���l7�r����;��Զ�B������,�2{R�O>!�c��g>#��ɯ��|�$��X���Z.%c�16���䣢��|A��NC*��������@����Ѓ$��;�UA��o%�;��-�(*m�s�C�'�^n��Bz4%��qٮo��s$�43k
2����1qP��r*�N�x���*Q�3�t ��R@7��ːr�\7QR��!�)���S��4Z����4���s�f6���F����ݖG���`d?�F�GS����5�wt�e���FK�?�]���+�w:�M��Q�{����5�L�&���=o+:𾣟Ǒ1x�,�S��K���a��1�o]�[�%��\]އ�c��xOh�H;ۅ�C�e��ǐ��ý��aDc o��nA�R���d�X�r*'Y���S�p2�󌮢��� �[���jK�H��ə�34<[�^����m���#
�vwM�"Nq�d�h�(�E���Qϰ��%�ɤ�lS��f�kdC��jsSAx��dd���2Y�He`� �V�ug�>���AKN�:+ӓӲ�ّ���J�R2�_��DOD��ꭻ�a+�2j:~�s���{
�{��p6��ig�l�@��kE��k�xYg� �k�r�Q��E*6�A^7Ԯ �| |j6K��@���6�u � �y��S^��� � �x_dj�W��҆JO�)m����iH��J�ߖ{k��֢�X}Y�]���,^�g3� �h�g��e@,�z��H���տ*X���i��5zӰ����3FA�u��|O�߉�|8|mh�"�0������-C:@S豑�ʘ��d�c���Bƨ�1eW�10S��
��UB�a��c/"���z,C0h〬$bqv�)Y"X�b�xIN�i�e�K��8��ą�g��Ғ8gIy�*���%�d���i�F�v��8O<8y�3ab����͠-vK}�c�@0�$8P��AR��7���s�l�y��!�h=��OĚR ��T��8���Cp��o�ټ#� �}A�-\��[���hȿs�|d0`���]:�_��{�b����GƑ��ɏIE�� t|���Yy�祯d��Yl�H�WB��x]�ĺ����^����2�k���9y��i�|�&�Y?����m*����(u�O�ݕ^yUz�F��5�k@�
��,fVr�2e}Q���-���k�?��Q�å���v��ӧ�0����혾�'9����,����A�s�$ml��NW�S�[W׭L�e��P},��ڏ�mI�>��x�Ң��y�d���AB1z>��ߋ��%n��l=*����~7�QM�GI�u~{�\�ޤ�*!4��Q�õ�f�F�+�����%ʌ<�4��at��u.{�X����8|Mrn��%�bH>F�?~/���^�G�L]����?ۖ���<>��GZWW�� �����:7J��,d���ܐ� R-_jvIfs�0� W��R����F���N�Q���k�]*�I���r�,��)�h/��Ƚ�2ː���esi���L(C���R���?K�>�rI�A�T��]uج
`�����kJo�.�j����u ��)P X$���b5v��iɆ�)�o�eڛ��o����L˒���Մ鈗�N]l�QQ�5ݸ!���}'L��7�H7}��1CO4㣷�:4�f��)���j��R���:�.#J�k��y�ѹ��	d' �Z�67����o��4�g!3c>��� W�
�+���:���`�>���m7y^��ސ�DA`uvZ�3�llސW�n�������d�Z��4A���>HZN�����N������TE�`��b�_��Z�D�����͒q�%i5`L�3z�\�Dn!�
�\:�Q+� q�d������5%_>!=�8FE
�b �Bl��? %%����B�����h�͆��Dd@a j5v�>�/�
EJf�lQN��?)��JX��#sO�-�z�#��$��9��Tfk������6Pq-�4{J�
�a\�A��´Ũ}�G�%H=[ɳ�q���A����Au7����$�.]d_OW�^�2���q�µFIoUF��s��疯��n��Yߒ�����	 X��0D���\.K��5�gY�悡��k�NL,�����������ǀ��KO�G/?���SBx��,��?�k�J��k��^hrYm���]9w��T�����t˓��v�%S*R< ��>;�;�����������"*Ta�
��f�^C	nZ��١T�v���D1Jz8P�J�������dʍ@�(�pGI)�Ƶ�N���o�yg�X�H/��(����T��(�x����Q�xX9֣"�X�`���,���G5�<H6�*�~�PF�a��C)��s�����������l���G�e|�K��g�S
��4$k!AR¤��!��G��Ǭ=#��5R�5��ho�q��~��X|?G��hem-�����cx<& ����l>z>, � ֯<':X!K�

���9W]��j�g��\9u�ݲx�m�|w{Y�\��߼��ZII'��8/Ǐ��˺ُ�L@vmS5>9.���.v1%�V$�q�~�f�
Gn�dM��=�a����8�k�+�@��ɾr��|���f,�V@����$;����|�c�Y]d�!"�"ܺ�Ӳ�ң�~c�+��%K��u����S�F��E:�6K�Q�
J!B�Ql�6P�D�%7��%D (y�He��.�A����0��G	2&p�����f���.f�HAp���1L$��x�|^�����K����fR�u8ƍ`�3�$�7̹p��آ�N�{���zGb�g�QO�)���M(2+xR���S����7�^{]��2��bT�ܴi�f�E��2Vb?��bӋb�F���^"G�/�$,Q�
a���1�����-3?\4�C��_r��@���+j�^m�e��HTӸ~�W�e��暾ƒr:G_�m*��w�Z�)i
������y�f����,��/�(�*&A%)�6J30*�m��뵤��9]V��'2)�q@&2ٙ �����	Y�Tڔ,Y:f%xH(���R�ӹJ��=z��0��8H2v��ݔ��|�6r� �H���M����F7 iS���YE��ݓ�,��,���u��:L�T����>g}=d.�.����k�m7xm�ȧ���ޓ\���!�R����y�\4N�x�����k�gy��3�\����mq.�H:gN'����4s��ŷ�"�6�S)���.:A��ӱjnn���E�c����ڸ�B]
��NK@!��Wr����]S�"�I/P�Bv6��#9�{9�ߐ�����sE���!{���Wq� �TFs���)��t��j�s
" ��|#Ё?��4*XF�*�2�E��I��{}��?I�P�|!@����f�Y�H||P)��d�ҧ�ch���R���ۨS����A�X<4��Oz��}��\�!���F�V���y7�W����:L6�MF%J2���q'��X+�vbl;z_ 7�y����K���0cć��h��5����9HΆY#��Pt����
�L�}��1<���{�(f3Ѡ� ;�]:�N�G���b4XғB$�4�NI��|I�;%S~J�<#��&�RU:��,�l˽�u]D ��*��|��ܔ��x^:��7��inr��Ӳ���E��g�aC~�71��L�(0�+N�A�א���]��S��������e���E��k����:��2��6��7�\��s��C��| ` 14wZ-���I!]���Y�$��mw�7���=R�P�E@�bh֑�J+����*�B���1I��-}�9I����PB���G�J#n$N�1#�u���!כ6@�&c ozM]�������,q�2P��*��Z�N_BF���'����d���T�Hxv�z
,a4���~Cf���[k�ey{I8ܣT�f�������rL�@�� �2*g
�X>*0J��P~�4�"B��� S��T��Q���1 ���1���	:����M��m#WjJyR0���U�U�u�
)m�=%�y%���%^��ǹ���4����O/�/V c~I����<j`��z~���(�s�����8�T�2��k���q鶻�Y�2H��x�gi	�6��XU�����l�%P��hJ/��h~���+�_R$ݑ��~"4�Qc��K�"���B���*��D�$��|����M���Hyz\2 �AT���b����#:o��T6-]%�'祧s��Y[�#��Ie\�cg:T��܇�pX�(����d�s����?q�}W$Y(����I�'>+�s�T�)�e:[U2�KY׷I}�W�����>�)�0=';˫��ڦa�U���t�2�r�@q���u���b�����'��յ5��ّ��~/;JR::oak��0��l6)�ʜw0
�m�,�9�V�J���.3g�1 ��SWbO�X�_`^�@����_#{>�j&@1��x� ��ͥYN�����Zm���>
&m���b�f�o� �����Z9�Yޏ����J�FEo�A�'Rۖ�����$�n�2(CB�����i�f���9�5E/�Ob��M��5��F��(3;����D�(ߒ��&��6�_��0�Sh�ra�`���F�ᱲ)�{T��2���M�NX���H��"��(J�2^�}M?���{����Dχ��{��v��V2�n6������ʦ2�.��L�46z�En���M]ۻ�y�.�&<���t�T&F��d�P,3Crg�.ݖ�g�T.*�3@�B����+��ࢅ�zFX؂�'ib��oo�������L�+��sb��lq\����b_Ar�M�o-�5Q�R���R�xg��I�I a4����"b�R(d�Є����.}TA��z�
墨�+�B��},��İ>Jq0�BXS�%�֡�eQ^7)n8�' 
x�vC�ٝn]���cĺwu�ʱ�N؄�� Q�WP�cC*8尡<�����}yq�����S)5��o������r�p]&a	!uP*�HF	��M�O:~�^K�w�|����g�_�7oHk��X`f��F�k_��xC �;���f#3n��n�	���d# �UB�U�۬���$�׏����/"� ��	(\�����#�,7t�Є6��`M�0T������ill�ܮX,���)wW��g�3�RT�F�J�\<3m��������jd�4�����x��4Z�h�I�<#��ݓ|��������������T���|L�����*o,�I��8�,}(���u��LIY�ZKA��d�Z�x0�P�ql0��lp���@24�Sz��*a�Т�'ʂ�aZz
ޛޒ�t���5i*��X�7i�n����&e�H
b%#Y�^t�T��҈l]�|~r �P��υ
�q��|fP�e�����mfj\Ν9ì��[��l��kZ:w7u߸����~�c�JJע�����������{tW�2V�(K�픤��aIʡʥq�� P��ޕ�`E�z�J|�zG�63�s�r��m���?*��ҿy�M�=x �
R�-���%�+6�8�^3�*[6�-t~z:�PP�}`�,�6�2<@������l�k�����H�DV���u����e�A䌼7T�,%Q�Σ1@��~r�}��6l����8zH��(�������hߙR_c�h���!լ��� {�1
���H~76�Y��}I��%�k�T�|Vt@�a�g��~�{}K,k�hp�ݶ��0�=�(��@Vc}cp
��;4�E,�p6r�ƕ}����(GX�]�:�]lwZ���o��_����<>��Gu����"`�B���{=��~в��(���	DBnp���lE-)�uK܊(ﺤ ���E��ݟ2�Me�V�X����b�ӭ�x�Z�t����Z���y����夠`��O?-���� �4�FΈ~ �52,�DlQC�e������7^��g�ʌ]`�ŧ/~H����[�����}��#�~��=ȩ:�6z_�o�Tb�~
pJ��Q���%���XmB>�ُ��'/8�l���]}N�4ץa{�C�2��l҈�Y��F��c:QK��&w�,��\�Aɦ�4��P�]���A�?��ɊXݐd B_FcӘ�$Ɂ7 P�'��rrjVN�/0�A�\2?z��7�G� #�_��ؘ�:y�D����KrlvFA�M�r�s[��0�K�f�.w�l~��o���99��eJ�~��o˫K�ŭ��A��82�!&��qbl�	��-�y��/؟�Ȉ@�uMi v0D�9'�+6�;{�Aʦ)_kS,(4�l�At����)sC�	$OQ`���1�n�
47۲�Ӑ�������������A9�㆞��Pp���2	ᛷ��<�t���|il6p4���|	����'�T�ʼ���3
J]J�vR����
����
�o*�4eugC�d�ƀ�3e@~ܐ��m�ؓ��H�-ˌ�F*S���5�J4w;��k[�{G�j��Q��[�%�h$/�J4	���*"��I4�57NH��P�t�t�YmoI	��4�aW	�@�����voCN�8)�����>�=� ۨ�Y�����e��Fb��̬�/�-��2�g*���u����D���)}�!��yWAw�ݒ�q�K�	���c��t[��o�J~����|�y�����s����M*�Ҵ���g�K��g���3���d=w_V��@ш����ױ}��������s����]Z��N�jj�<�O����s����\�1�!����K��DV"� �V���@#XV6�8�dʘ�b�u��P��.��P:ʬYh�r�u!�d�kz�:�B��`�T��=$��
�8܈��!'GW�ˡ�aU�G�u$��sφ�Q�	SVxX�鰙���?�t 8�;�u�t�0[��u$�^��ūws&��z+Y{P^k�G$FM����h�w~��;�����G�j+�U��<� di`h�z�������|��c��x|�W�b������Q;l��t�E��G-�.v�D$#qV�|<DJB�� ,�/AwC�u�%�����ֶ��%HJ@JE����S �Оn�-%]]���/U�4ݚ��J���/�
N:��腉ܣmL݈(��8q�&�&ۖ�s�^��y��9Q��^�"O_xJ����ޟ��lyM%$�v�����SYSnB9K{�15��Q���W��KO�T�����������+ߓ�(��}6��;2�)!����P豘�v����N=� �$�n_AG�D��� e�htQǖ%%��JJ#b��\�9Yd_�-}���9fW����7n^�������:u\&/���x��X���;l��v�L*)���d�ȓz��T������m9w��pF�Z���x��ʋ�_�ݰ#v>�רc`�͆�Dc�9�Y�pHb�M)�İ�K�܈�'Iܠ���-^��I_GBN٬.�wA(-��1��D���a�G�~���K^�BssJzubRB�[��x(��v��s���Ɏ���������ݒ��q������-ٴ�U@����(��&�g�9j��J�:��ͦl��XO������xe��7(�j��輰zM}����7��X��gu�߀�$�d���d��I�o r��f\S
���aʇt�/=!����ĦiԿ,������Z�/� I))z�d�����v����̞d���00Qx�J��]	�V�.�����o cM�{}̫�PN�����H6�@��'��\jV�Ͷ���N� ,�)p�����"�$��M9�<�{��Y]�@
�ΠH����'ul#��w�*���Uq���Kv�ץ�󣷣���E% ����~V.M��3]5 M枞WI	TV׼T����re�my�@T �W_{En�}CI�QD�A��h�w�/~/�/H*�	�����~iڜ��,�"�)������"�R��yd�o~�bf�a	k)T��ǥ��萲�/L�^������$���Qcc�2�Ԓ���%ِ���h��Qҷ ��j<f>8��/�:��x�GC��Q� �������s��(I:`F�g�|c�&�$jd�G3Rqt�t�Ii�����\��{<H����\��׿Cyِ�X)�.vҨ��d]�ܺ�u����������y��	���=}4�J:r�t..�v���p��N�N[,�b�|F����'���~�Ί���TR��hh�K��`�(���i�x�*Uݔ��ɥdwcMnL���OKU
���)�Kw����Ț�#��n�y� 6�nl�QY�E��d�%�u�R���?{��$_����W>"g��%��0�����?f�ǰ����a�����)"�>Oz7x`kO�X	��_���k���g��(��Ñ�7�h�vR�I {�ӓ�h�}���v$��1zi��fn}�����̧LS����
�X-�e�'��o"G�L�\�@��+_��ĝ���
3 � ��g�E�u�G9#�zM(e	{Jnt|+�M�pͷ�-R�v��G-xi� ���G%�D���������*8��׮O8��İ�4H$cʥⰓ�df�6�c0T�i���mp��Y�a$��|�ĸ�+�A J����(˳)���ɜ��g�@����O9Y�S� �b�螼�xO�o��sI��%P�bgK9�aXV�����lȲ�!��]}�%�Ō�	�@#bO�������F�!��{67^�byZ�tNz������ko�$S�3'��f�6�d#m���܌^����2����]���i������ wn�%��o����x⊜:sA�>:!���_��	%�~nIϽ�dcR���I��GZ�k3�ect`��O�7�a���F��z�<:���g����+���}]\F��^(O���/���%�d�x���Juu�QVTRr~��}��R�"�;�Tz����ʲ<���T�B6h�ՠ�t�ۖ��M)*a@YX�:Ʀ�P�m��H�6��r���5���Z	Ǯ46��蜁�ǽ���g?�)	[{a�u�m;�ǐ%T^�M/�b%O��y�ItemyCf����̌ܽsG�Y�;%^0	���d��8���q���l��hj�vC}߂���-�R�$Ғ���$�x��@��AR�
�lF�ˈ=4�Q�����3b#��fe#���pxOM�aCǤ�ߑ�y�����3y�4�������h��'EIF3�C K���åWq�C'�w{�-�_4�A�����z�2���a��^��SFn�p���� |�����*������9���u�u?N��(ճQC�������|�ʙ#�`u���ݻ��+�/������1y|����7��޲";�m�YL�Y7���h�Y�C#7��
8��\�k�-Y��[�R�^��X�-��G����q�e�lF�m�k���ϰ��"ǟxVv���֝�����+��|AZ퍤~��{G�]ol�Y|�܀jQ��:�����ͷ��������I�2�x��4m�_R��^e	�4�����%j������(��(d���$��տ�F
ҡ��}�J��Y���!mJyX��L���Y���81r}rjA>����9������[�oK��� h��~t�%n���'�����)�BC֏���v�*V)�!���r����,]�mF`]6�H���9��B` �/ Q��9ͺ��={�ԭ�������$hP��N��Fg�"��L�G"0&��H�N��,�v�p�3�k�[�sc�8ʅ8�N�d�d7ظ��(���;0�0��#uj��M�8�LOϵ�l�g������U��ɽ�U�䝽�$Ƕ���%07Q��oI�QR�VB�s=���XI�G���Z�g�g���J_��}�(�k���)��NLH�R#��j�H{u[	������,/JY�kN�z�T!Q2��!�7%Y��e��Tr�����s�d����R�ψJ�w�u̧dLA:�Z�U&�U���k�%��/~�����'$ӷ��)���Ɔ�s��}�������|�̖u��R;yQ�\����w���L �����ą'�S!�Ff�M�o��8��8�^���X���%q���r�N�Ѿ��������o�%=�+�ͯK�g~^�U�E�K3�`i~v�Bu=�����ޓ�W���.�lqvRN-,HN	`�7N����l^��ed��	����s�N͜P�	pjɥK�����������/��h�$W�s�[^O��������#�6�=��cm��d�d��4�kK������
Q���9���J�AZŦ�z�TI(�t�f�()�{��!�bLӖ��	dunf�,�����3,J��=���P�}�x�hxR"�N*T\:�L�Q�2=;�bIB:F�K���0(�~�C�˰M�yk��s8cd�Ȭ�@�2�ލ#�ҭ�4�SY'�%�Gc�aV�p��(Y-�#CѾs���k���)+�r[s�Z��L��m�.��7�|�}M>p<& �/��ۿm��n��m�Y�jt�O�>YT���){�����]��t:�'OFq>����n�7����n����ri��n&�V��~v\���zϯ��|�g�n�M�y�z��5��Z�Ъ׳
�Ү�:��ϳ[��0�� �r{�J�WH��^�(c�w[�P7�@Qߏ����{i�	�� �>��{7��AH��z�vv������hB�'B��lu��Vah�,eq9�u����#[^_�)�i)���� AD�065	N�&�ԍͻ\�ɔm˫KoK�v�PBr�L.-�����<y��Ҋz҃��r��HQ��8�-L8O7I�q˗nl2"��'/�\��_��|�'Z��;/�T�`��܃PA�e��Ԥ�0r�f[��`E��h8m�m���G���$.����R���f��k0��Q��G$d�r!LS(�%d�N��Ze���Z�����S]F��= (���Kd�2��D���H��;�@�XO�_�Hj� ���(����\xOo��9A�诂F�~�g���NLΈ�ϋ�S{F���o� �K���X.d��,� 6�r��=!t5�G{#@V���?4���"�4��G�͜Ʒ��ˑqu��²/��1�O�fq�����(�SC�嶲�f���Gi��l[��|���!_���ɩS��:�Ȁ�Wd���^Zb(P��R���k��(��$h59���
7���>�aEIʑ� ׮|��?$�\�^Oh����ރ5}�ӳ�t��8��-����Z,��et;���+��hu),017/�޾%U%΢D	���ZU\h+wf>���W_��r�<#�H���s�eH�"g��ߊ�S�C�!Fف;�V[�'JEN��S��[[��ڔ|h~N�)�(t[b���m�M�抱�/�狛d�b]C�I�����TA��g����o^���ߒ�gt�·2�.��蘝��	��b+��?���������9O>������<Af�\�~�gƆ�:
c5�*����PF\ �Mg�29s��H���-�V���믰�ll|\�����t�����{(�y}�ٴ��>$�3�	����!�!����<��q ��`���`���(��{����� �Vt~�]Y�q�M
:���$]x��z/B���6w�T��G����@��R�$���z<B���������WvuT�cT������Ќzx��`�8�!��m{�1�<�z��kH�d?������u�^?���팖n���%u�{\~���^�����2�d~���vwwv�B���»�����1���	h��o���˙\�ٸ|��ӗO;}zmy���Ul/v���D'3'l�(,�Hyc��pN7�b1t{6�s,h��+�Ỏ�KZ
���#����Ͷn� =�fO'��^�#�r��)��B_�h��4�0lnm���<z�9l��Б�(��#F8��������]�ܰLH7�v��A��'�߷��~��z�b�ۉ
�B�j5�t&��@�@i@���B]PG��`����G=��~t;�ɬA���kC��V�ί����l���e��;zY�\���y�2[�=�����ܫ:6��.d.�YE����0k�f��l�H��L����U��GV��zز��I�/(j�u��-O�ֶ�tS����J���NA��I ek��k/K�����$��r�.VK�l�J<BICY�n�²��v9�:W3kHD��k@ �����m�_+0Jx~��T�r�D���Њ��I��������!@֍<���@�u����.���dj�C�4`4f]8���ᢋ��S�0E��1r�7k���s^��2�# 1	����V(	�6th�Ŗ�b�8En#���$ݓM<�2�nD�u�M��i:��$�������5$ s��NƒR�hz.�J-� ����X[5�I)#s�(ۨ��I���H,��'4[�jH�D*�$����ܣD:}�,�@�
����+?0���eWQ~C�����`=���A��?���X:�S�G�R-��˿�%��rWז$s,��\��e└�yi�}����K�fD��~ ,�:�n���t!��1dh૓
]��g�q���z��8�}�d�^�ZUV����%������3e�)xf?�N]�B���X\��.Ô�P��j��ꪴM���ˍ��cxq���65.�7�K��II��7��kr,W�B�Ҍ4��%Uݮ�`�Gh�i�7G���|�q?�1�49����|`zB�ժ����T�\�Pֵr���q��}���fm�>���e����gΑ���L���+���oIS��׾�u��������/YH�C0 0%���xߓ���>Č&K�<]�����+o��x�D��%-B>���
i%�:�2%ji�Y�t�e�W��)-%&�sJ�k5^�������:_��odjУp�����2���t(b�xoQ^z���x��f�1I��l�ܭ�:K:���1k�~5;����^�[�ǲ�����}�����C����n]�]ٜ�"���e?�p�D	�=l��'��4o��4�<�=�������wo	��� �V���+O2��� �h�T���0�AY⑦s�˶�̅��cU���1tF����G����9,��/�2�q���=��$�aǁ�8!��~��!G+3Gއ�����J�ӊϼv�s��g@��Y���J�����/��s���h�>�ۓ�qI������d[6�w������!�Y�6& J.�Y���e�$@�Ӎ���dӔe�\�����:u,�,S+	��m��9t8F$ɉJU�Qэ)�A��0�v=�|������Z�A6�9��@\�1��L6e" I�ixU jC�ޔ�D�I�.BP�т�j�T ��t����b��JD�
������nWAP>�	詁k�+[�\!����r-�_(Mf'ܻ� ��T�U��c(���3���� 1��]��� ��{rn��L�LJam[�B$��i5ven�&%=�)���ezW��+���ސn�(��@���g�����K]aُ�˲t�E}mČ�gЅi%��c�{�F���&a�$D��\U�y�eYZ]����_���))(8H��H��g ~S7�Y9-}��������r��.�T����942���S�����Z���Bd=	 �k�-Q
*;���sG	���E�v6��CWc`r�
@��P
TLc(@�2#�k~�x��&�E�L��s�Z��"��d�7��&������2�0��������Pu��@%�����ЀS'��۬��3�*�){��4���s1��c���� CSB������3�x4��񅇅�PA8��"<��Q���`1��C�iJzz��/ސ'���1O��,O��HO�QuYzEO��.��s�Nl�7Ź��+�w��kC^�uM��}M��'�J�����'����>�z�97������T��YT4��#3����(��>�B�`�
����P�eGC�����IC�¿����s]I��O�\�S�\���~$ޛk���|���RD��N�^�-;Jp6�W�,3��:����^cI�dhƫcR���:��UIX&���TAfƞ2*q����-��6�������F+���])��`,�
ڳJ���ץ�ϓ| ��h��55����uiV������������ԑ[���/��W2W����es6=Lt̌��_x�XΟ�Do�?��?���'c���ۯʸ��X�U�Ί	h����I������sdư�o�ڃrǹ�y}}C�^����_���NK�Zұks��(��L��ӧ�\�33�zr��{��M򙝂�7	�%�1��_�U�[J�����on�Ɇ��]%���t|pS���8z^OZ��d�t��G�cJ%Y���z>�eV;��cT�� �m֕!zx<����ɡ���a��;��a��;�Ś�:H8ը�޼Qb$#q|����M,��9�~����@_��<�c��f)ec�z����[��H�ʁ�4�p�����0ϒ�s��� 1|4��٩T*.���X_]]���l��X�}�����=���S���������oW2������dCs!_�J�d$u��W(���ȡ�<� Fh���%f �
E `�?�<��pH�"&u��Jd<��������l��`��6=zds9�Օ5:H�""�8)O���tM�"�v�H^�� ���/p��Yߠ�,%݌�v�
� `
���
�Ⴌ�vL�k��3�2ܸB����S����� 2Q��������H�g�n�$P�����	n��1 ��/�2���D%���|������|�K� �/�%o|�99=3'c���v�I}�9�e[�ǫׯ)��@I��ZC��Xҹ��k�Kܪ���E�q�LOȠ�!X��(~�������8J>`<Gb����<�lZڮ��������?'�<1>gd,9O�L�P�����wyϑ� nv�:�=��^߸'�VS�Y��c�(r��HB��6�~*d���~
(���(!���o����o]��|��yQ(�D$݄Xa�`�\��DL�R�.�>�?�ۏ���8�Gy
M��O�F�9=�1j\ �4{Lz}@�Y�R�<}3B��ЬMAՌ2Jrs)����4���!76��r{S���06i4�y#CI�o�cd���e\���p^�i�5ۓ1p�KL���t;2d,0M��EM)Q�G=�����dМ���{"��n���C� r���0�s�{_�����'J&��P�	����<�e;]d��@��t�Ja �W�R����Q�HwraBN.��������$������s�ُZ�����B��X�.�!��}��i����m������JK6����xU�����\����b���q
�we���2w�4E.>q^�˧ٰ�E<0����[PRP�O}�Y���<�������^��_����2�����іޣӧ�A�����B��c�sz19h�5c]�P���xR!!�Il3Z��nwcɇ)9}��J�RQ2�����ٖ���$�3z���xB��O�Xz�^���|fr�Y�+g/������7޺*WCd�rtDG�%\O)x��'��+��܎��GV��e��9�u$�iyu��.�R�M�p{t}t{��M�s��hI�ٓ��{�l����K���˖�E�N�Ji�W���s�8_����ymE^x�u儖L�����O�:�/�Z�l�Av%[ ��;Jf��<3&�zs��d�	���t4x�Ȍ��9�Ay�<�~��/�;��j�%����$.��O�ٚ�b@o­�7��IbJ��!���k�~��Ao��@�hSե�K�{]FM�Q�ü)F��&��09Iư�m�����P�"��*�^m���my�8Iȑ�2b8x��f�z��?F@�(i�{"G}T�*:��{�s���� E��<�������At���z��_��w��xL@�����E�`'��UK��Ǣ��vfrJAQ�Fg�x�f��|�ȟS~��
^��d5�[[���	i��n�^ �B�=�KK+IɄ!
��d�X�+�����=9�p����ؔ���P��*�7.�����l�d0�J�߃��s~��4����Y�l�u%��sd�<ܱ�V�,�8W��(R�(Q2��!t��d�����~i?B�h�a�[��[��-���"Yd���<��p��k}'�F�ͼE5��R7+3�ĉ�|����{�2c�\8QOAh[�n��=��*��f�������{�����x=���L�g8`�k6�����'y�ʼ6�hd�nC��sЊ{��]kT}�IҲ�h5[`�g�E`�l+�4hK5��Ӝ��z�	���-���ًߑ?���ˇ>�f9[���X�ʙe���`��2/��X��n&�̡���]�@V��7Zw��7�d;�I���ݹ�t3n��^�����͞�O3cL�͸(���4*c3�4��`K��eԾ-o�ߖ�����loni\��v�w�z 74"�D/Ӏl��d�e�^� #l�pR��Fx,�[F�����
U�5��=�Ʒ�L��5�i0V��(ֹs7�}(h��,p�7fQ¹E:b�r��aC�|�*�8����������%�)��;��	�7�r�����a��3�znC�NH�`��rc�\�}��yD9�X|F&+j�|H�0ó�*��7��MG)��$Hcc�H�H|y����� ���%�N�0g,��4�끔/��2+�'R�7�� �n��\�o���)����O�����ϸ�jL�%�їÊ��2�B�{�Bf�ށ4;&K���9��y+�Ь�0V%0�w�y0< v��t�*�@g���~E��ߓ{�t
zm:�"�	���͸����e��ug��i,4X����4��	זQk��iM���G���9�Q��9NFrg���۽)���2�~�*M.W�ָ�"���K��:�jC,�x$؃��]Vز�>]Ě�6�`r��%�KR����Ҋl���0	2�FC*���fpp(��e�sdA?ç������Ody}Qv��x���5��bͯ|�u���%��_6�=��-��0�o��;�w��D<s�Y�B�k�}�=!�������V[P�/���{O�v�o���X�����#�^�B����Î�͖�}�6�P	��<�u=�\�"+u�U��އ=�܅�4m��97� kk���3š��H�Zcet�(��+�=$,���󷶶��*�V�� V�k�T��� �P�ӱw�;����!�%��u&�1�����q������1��	�%Ƴ�>'U6f��N�b���'�n�t��ǯ�led��P����x�l���>�h{�{�$e����,���\'�)�G��ג��׬��d��>��I���+�0��KT���G ��ﰞ}��r���F��ʅ��to�^��>6��+聎=H�B/���4e6Y[p�Q�Љʾd�O S��
>0y0Y(6ȐG �
1z�eV@OA��s�R���4 3��Y))8`�����ں�b�/��[�x�p����0J�!l�i1��k��f���?H�f�Ȅ�A�>D�pML�����>p�!� 0�5X(dlr�Ƅ���$�-m(�\XI鞣�Z��E��m�)6�̍�Ý�>X��jN�L��<��c2`��hcS'�vБj�$�{�����W>��|��Srn�#R� �`�l�(�hޑ��e�i�$�y�nAZ�#�����V�5<���1Ԁ���礮���7%�F#�
-��^���۔��i�5����<�f	�񂾟qv� h$��P���fI�:��(����8�����
�*	��q:2�(�G�o�n�Y�!
ܦ�Yc mOztF��������S��8�QdJ2*_١C�����B�p��O��"bfbM����B� �YR{��m	��R���Z�Ю�bn�g�"J����P4��U���x�8A�aAi)T9��-���2�����݃M��ih�kL�)���z14Ls%�'{��40#<��9 ��P�М;YYr<H�&��j��;2s�-�gp��k2�/��>�:�b�Wp��������&g+���OJ���/˼[#����xf<1?�z�oMBZ��q�-���-�-	�}�'���w$,!S>���M9��&�R���ʣ!Ʊҁ�������x�OIQ�z�?��_��C�>ڗ��Y������^#Pi4�G�ູ�-��-�zt=Y?{VA�<?�A1�h�P8�b��p�B�5�<}�q�*%m�$v<����9��_�q�'�-�[�����R5�%��2T1�U�UȂ�a_|a���S�Z�݃}�G
��Z�a���z�@�st"����3�?!��
�2���9(J[�����x<�=T�zB�͐�X/���� ��߾�	�rxБ���rq�	�H�.�ASΞ=O��H>P��|��[oK�}ȪCW׾^�#�oߖ뉮o��D��@�x3$���/@D_����Hn�H����(�%/��U�r���
SY�
,Pp�>Q�5�o�
|�o�\�E]SG����d��HD���!&
*��B���V0_A�
T5�� X�<��s"��i�z
��6Q���&r�d���<�Q|6.=A��8�x��2��C	 �xv�7'����	�O�ٞ���P���6�YW�:�N����AjXr��M �QJ���M+]�L�PnV�]�YQ8�g�|����4���f�/�� �����Od�=����a���|UmYgد:>7|YV����K56���lV�".�h��s��JB��nl���@/�G\,�����M ��v��к`��yxh2��8o<6�ޠ��Z���Ac9�qC7�6+�-TH|�ٰ��Q����UO�Ftf<B�hF�i;`�A�ǂ �;�I!�������&�פֿ�1��낮�ڈ~ȠY��N�  *�N�e��8Ե�����4ّ3JKu{a��\����4��!6�	������b�W�����ơ��[ߗ�^}U��9Y���<��X����Cү9���.{Bb]x�����mY�tA��y:g����BϹJIj���vP�J	Bs]���M/IYu`j�6��	%E E	
���EJjB8�Y4�;c.��U�@��[P�I��3U�wL�^gLT�6r�\M�IO`�AJ c�+#-���չ� ;�I��m����6����vp"0`ӎ�zP.��)-b���T�<�g�1d G�Cl�z����T��0�6,����82��RQP©(8Ӏs���Y��Q{�����N����}����3רV�����=7�Do�����N����r�T��������%���6��tr]~{F߀�=Q�N�_��6=V&m��s��(�8)E$�p_v���\nߕs�+R/զ�M��[�����7��̄����+�;h�/�ZgS�� /��e���[ߕ7�ޗ�J�:z �`cEA��T�Ą�A���I��wK�ڻ2 ���I#����1�R,�3e���	i�6=Nl�#�T��G�W����s����9#i�]6</�F(Fm	�$yp�������,�-�:Y�-Ь2K�V�s�w���F�	�C<����i�������M�蹨(���	��ʅ2��@�RG�Z�� �6V��.�w��X��7��{��@O��������(�ڜ~��	QY��I�Q� dA�O=�P�s������K�����!�ef��y��D�
:��Hn]�#ۛ[���#�[�ҁ����/F��0��gv�sp?��F�J�b�y�G0cI������x���{\�����x�'��[�@�E�녅P�C%��bh��g�^��r&���m�6ee��R�&S���!����>��Չ7u����<Ǐ�Ն�c���0~\=��V���M*S5��s�F���.�� HOÇYzJ�
�xX?��cm?@�:�=N�K9�}2#��$T3=����{������o~�<:x< ��a_�ب�ϦI����.xO8Y���^X����6T:��	�D1���N�n����(b�Ԩ���j��X��;�,���������j����(��c�D�36�Ã�4�M>KKK�X9��@m} ��o�l�@��VSJ
$j���t��'��B=��ꁍ�\1*9+++znc4�MܵM�U�^�*�@����e�Y.���`�F^�q�F����X�@�7�x�B�Md�\cn�Dd~?v!&��2޻�c�Y��L������n޻g/|���i�%,�Q��+W�A�� ��e�q��CoG7�ۇ[R�%
�^U�B�n��n
�q�c�,��k`�Ȟ��J���n̠�8�ҋ�O_�C-k�� ��|��sK�����
Bǹ	��,����2��!$$��`/NcSQ��f���E�P���}���NCc|�	50��3�4#�.y�S�C��!@*�cظ5���ɒ�Pۊ�����M4AL�4�R
�S�(ة*
�<�#(��5�PpB��9[M|�o�e��p^�r�l�Ο�U"�@���w|F��F�y���+�P�%H%c=��.��+*�h��k����I�)�〕	=*Q��Vt�m#��{ƾ�E�%�m*<z�1�CO�b( 80� jqO)9���j�:� fJv� ��^PY��Ƥ�vX�K�'zT6��P�����[�_f�ͽ5~4�=uIj��
���Yd�b
f��0�âΟ3qSc��?�2����%C��574=;>zM����h�G	�m�����&WAv��Ѧ����� �gǣ�B�kO�T(Y�qNr9׽w4�-S�kQ�$������@&�^g�����yp��y���_"�c���w���Z&&����}��9f:�3jD�j���h".vΩ��O}�3|���ݔy]�����K�����<��/D5t.��wemcM��+g��������=$�l���tG-�,�ɽ�%�/͑��UG�u]7:��eOF:�{������+������H���x~��@�����xHJ'�r��@%1т5��' �|�r
.�UT��fYA��j����M�1��c�< ���Ta�=c�C�\�
�k/�wo�Hx� pD#b�H2�g��x��| ��y��ؒRcE��q���4��l��S��\S��u�bd����L{+���h>'��I��T��l����D=��y���߯�M��O�>��փ����մ��>�`��^s�nk�`���<I��F�"�����c9��yp�S
�����>�+�c�il6|>�� �/q�={���ϹV�Y�..0f*xe��zU������E�Lnk8
���Ho�r�n`���e�~_�f�@	��5�A���>*����/�Y[]�E�L�
 �z�T&��Z�p�Yi���<�0���d����&��/p��f{�yh�y}�M��z��������X�	�� ������`4�� 9I�p�q,��Ud��c�E5�@�d(`��ܢ��9��/� ]�Y�\K�hA��.�Kv0�5�[\�
c)���Vf�ya��a�u��K��L���j�ӑ��M;j�[����`7���4�� ��Q�����ź����R��P�ˋ�"@e��#�n�h&o�VЪ��h�e�db'�Ah'����L+$W�ُ�C�'d�	�A6�>1��jQ��3�&���WЀ��Y�\bf8�6���)�@@�hI��M���cT/���\aG��h{rX�m�B�5 ��V�s���KV ��5�H#�e�w�B�g���3�N�-9y�t&�G��@^x�U��k?��+$xo��	.<��u�un�A��qD��5[��Gլ$�޾X!��dWYq*4���%�+T̛36j���ަ)]� ��Q'q.����ж@�ɫ!�U>�]��.���W=';�|��e�ę��e�C����G���t��l�
t\
L"��ڿ"s��8� U4=gu9�'�S�Xz n�z|T����fU��0��40�v���7�îX�^$�EDe�jo	���� �q��b�U>����f>#؈�J�"{&x��ƬqɌ�"���]�=�!���~fL(S#�@�b(��5�0p� �cO?K�b�чz�Q=�X��'� ��Q�-�r!�pa4���,�w1)����*~y
M?�3�x����A�������*��Ue?8du�X��:���KqeN*h0Ϡl8���F J#�qG�җw/�\^޹"{����p�9P��t���[Wu�Y�ΰ)��;2h�e�iK��`�:	$!�
j[
�b�$j�Z �C�!1P0����X]�^0�d/�U�k��g��g�]�7��/�K1��9�UŊ�
6@���r��ZI�ӄ��O�/��C�F	�"���g��5��s�}k�����8.;9~���\�O�J<����R��=�5f):�Zp�\�'}��}��>����Ǳ~���z?>@"w�Zf�1��=���5�$�iU��?;yl�&��4	�R�h��j�?| �� �/qh�QL������T[� ��j�{y������a�"��P:�߾sW7��J;�����r!�B�*T�ʵ�!q	�	u�" ����w�e @� ��;}n�П��.ύ
N&�Q�҇�}nl��h�U����+{�He�� �NK�u��ߓ��%�Г��~-���uf��<�Rz7����<xh
�j@�.O
�� ��o�T�/�4�X���M� ����J�@�@5�̄Պ%<�}���x��j��wF�#�\O��$�_.�����[�,�#���y,�^a�5e���a V�*D��Z�ߗ<f�c,���W�LQ-I3�m1 �y"��3���ZAo@��]m�J��a�m�I��c�P�{f�C8M��k����^GL�#�:f�@т�(g̈��,��T�B� TO�+�=��R�'��ĖQAq�> �oԤLP����A�DJ�k���0<�h�ISR ��������<^]�9)��<�}2�;��5V��qR�Dr�a'�����5��*x��߼���օP��ب7�=.g����Y���(}��-+
��
 =�"%�(ˋ����eqSPˤ�e赱bi��8�2������7lw���w
����@�9@��(`�������gb���N���L�3�~��� �.��� W�p(1��{"��L6f�*�����=c wҰV�RX�=�up�Y$�F�<��=#X����l_���Yy䣑�G�[�I!���aW��@a$�R�T���"xw
T��3xsD�^ )WPnt�M'��|n裩^A��i�����Ԇ�O<E��s�y�~�솬./���+���q�	�y���?�}��b9Ɨ���	tr�!���qȏ{���$$x�9idT�~���^o�P}�=�d8���}�y����O='�
$����zB�Oǹ9�H/�{�w���k:��H�7>���������\O�����%N�ͭ�9=�ڢ�z	w��HC�q������Ŭ&�L�'�uͫ*p����ʮ��W��
��!�NJ��cxX%�H���XM2�H^����~ ���ѥ>FЈ��.�z��@jI�U_�����T[ݯX�b�/��y�F��^��3 �(W�;��3��G�W3� G3�'�}��R :[٘���O�/ք�{���K�ڣ�0+W�Tm���%=��L�	 -W
�iNS����mMհ�\���8�?��Ь&�c��~�|bΗ�f_���x�'��_q^�ʍ�H{���^y%�z��?x����# �Ks�:*7�['o������������dC	���/&/�G����s����aˮTkL��4�U�<����޽��07]8wc��i:8�J�ZH��U�}���0���6Ҥ$��'ۇ�T���<l�a�B���@=����OC�g�}V�]�&��!�!��)��Կ�������_D�{:�l�H�t���a���T.D#tci0��8,*�n��(�5q����&�wcs��������h̻�Z��  �j�2r</�F�8��ѭ���W�(nc�����������(�W�K���c=���^G�P.j�$��!U�f�=.u��P�i_2R3@�w%��5(կ�����F�_���n��̢o��`4� &_)]��ʣ�8�Ѡ#�R�z2�3�Z_V0�gR��-H'�勥�4�4ˑ_n�D�$��8q�M%���|4�I0/@�	�#l��Hb�8"f��_L@@�*��]lȹ4�m�����Je�f9��ʕ���4�\���w���\U��/>��T]�E�u���$VX@E�L7$[��_JƆ�\�6W����~S�sl�19���.��_��sՎ���NO��k�򧟓3
(Z
�K�5��Ag_
��>����l�6���=5/�n�����u��P��_ydĉa��osl��G�  �[���F��P?J����6�"��33�\ 2�����Ӎ٦*����6^P���P,UMk7�NęF�+MI��U<�_a� U��AT �-2�h͝6�/n��LH.C��\*�Ԁ���M#&`'�ƍF~T}PI���jWp���-2p��SA2е��?i�F����YED����48�%���"8(���:~?�����4�ͫDν�ܹyO��b�&���Z�IKPDC��P�
$l��u})7�8ր7E��� �?Az��
���2�d�r"���@��O�s���0��,A`�y�� <�Zm��� �����T(Y�����c���������4�]�q}�^S��}��^֑��'��
�k?�]�y���NqP��{0j�7��:��bC�z�1�p�q���VK{�|���+�=��k5Ľ�X�VW�e����BP��/��ЛX�ɦmL;Y��hy 0��4��r�&b�yr�3=e4����&�U�RE�����%r2c���fݫ�=�a�����3�=Ǌ0*�M����G՗���>�a��^J��B@�h�9�s�'�'�������z>N���?����9Z���lr�*_���?�mJ?~����ד�͞ h���I����s`3{�N�z��H��ԶuBT?ƺ�����7o߻���(b<:f�G �8�ܹ����?�Ǻa?�<8�zj�_�i\�, `��Me�h,�`L��X7��誻������
N�~G/E@5�mdК��To�]�����̏�w�2��q�t����{�l�8,d�]S���ễt�mf<�1��{�����|�ph;�8������-�iD����]]����q��@�����H�J�1l�;�W�#��F��Jlk��+wG���I��:�IÜ5�������d��tC�%�[r@�e��>0�!_~~c噏~�B��˙Ɩ_�$��H#��]`����HJ���O��h�g��U����,�
D&���l����yw5@�( H�݈#�2�ٹrV���ȂV���%��Cl7`0
�%�����.�y3�ڞ�F�s
>��&3��a *3GY�y�f�>6z�\j д���7�5�E��ff�����6�:�6�g�W��0r�&��[�Y{��>9��LL��c�E���c��g��)J�&��$�d���f��Hn��a�Cg��r�Ɣ����������|� �3 Ͳ>;�z���[��0[=y���o�	5�s��g��d�0'�qVm6ʺuO�X.�����|��������Ȏ���bɗQd��U�,f�Q%���
���4Y���<!0c��677N�l"�����"��G���^��=>��Uz�P�
��T&&�%NJ2C=-����b���p��4�#!���7��Ybh7�V0��W��(#�B�/W�7�,?@:䦗�$�*���$���Hm���V>����`���tl�J.D$tLB�e(�A��-S���o UEC�	%��@��a�r�j3*��N@àݖk7�0�0W����x��`��a��;�I���Þޣ1��'�Y��$�4ɸZ�;lN�9'hDYp(hYU��X�Y����3�j+X�ڔ�~�,��i�  �}�`_����*�Pћ��TpB���Q[��^{IgA9B�������,����s�+d�ݓA�/���t���u�v�>"A���T�@�'�y(U���z-E}6�+��^O���s�n�9C�{(U�b��"�lHCg���#.� �#ܣO���<V�,��<��R�m��� Ɂ�G T�&=U��� �K�L0jۀNP���?7U
k�S��>���S~��<Z�٦��M�M�}������	���	(����������Fo~o��Zo�����Ȝ��ٲ.5^J��q���54���,7>ړ����鵛�Y����?K��}N~�ֻU�]����q�x@~�#}��W;��?��u�����]�Z�\e5p�������j�b/�-��mǍ�3�������ۺu���8�ٲ������	�I@����7��G������ѩ��I�� ����C����|�Q��e}}��i�4t<�jv����h鶬�i���/ꇭ-{���M�-�����0z�o1䭙���A����88���V��F�d�$�B)�����O�ZuInnݓ�6�K�`�j��ؑ�ؒ��ߑs�E�;�q�6W����1�[
"�폾+w{��/6*0��_�=��c�r~]�|@���]�o�H5�j�b>�@Ð��	�R�a�c�6���/r�)�b�%�gvCؘ,�T�2�T��z�΀�EL�\�@	B	�A���|Τ�0�����7Gvߚ�&�nZ GLZ�e=M�H�h4�Y	 H�9w�FT�J�;&�y��LLF^�,e3�3jRi�e��P����I�T3=G�/Cf:��l}A_X�����@^�ַe�ގ��V{FNO.�=&�k�Uu,R���Y��2i�UD��R�F��P���>(X�_$���C�7��轈�~�� ��80��NbQR��4�`8C�Pd�i��3r�i�Z��=�MS;�Q�`��I+i��&#=�E~��߸͙���t�N��!�I)���	�RQʾ�H�'�T�XT�>zq�6�9q<M���=	9�:˩���,������
2b�\�Ҩ�Hm�(۷ﲑ�H��Ј��#���	U�@{���)n��ߣ�K`<�F��`0W�
��ժ	>��ȤB�oayI޿��[�R�"[w�ʾ΋3�����Y�\\��!;8�+�"��A��Sf���$عTjV �8 ˲�չ��N���'=��u?�jjЎ���]9�Ֆv�/���ߥ,o�X`Nb{gGn���E��Ų7ܔP��P��@zÎ>cYb]A ��B�/�i�����|��!�}�lwdtdG���>�}#����Ā$K �Qe����x��_��������< Q�����ʟ��g8�i��k*��zz�PLC��ջiw�ՠ��u�iH�@�^r{K�S������id�x��aY9���M��g��*�/��M���4_2�|�I� �1=''�՞N֨}�oNz�DM�#���>�M��Úi��Mz9�_,�8��S��}�cc)dR�i���mg)S7e�6B�R�]]�={v����#
ֱ� ��9�W_������y�#/�\oE��F�����1��Pn$g�G!J��喆s�����[*Y UA>twg'z֍+���IoDnl'�j5im�2T���$n���J�<��f��â�Ff�i�k��Y�A�n�n�/��I�^!�_]�<Od�|���cceݳu��=[Z�k`�c�"q�-�K��?��o˒T%��ʟ��W���U*S������%)��5����\�6eV��.��^(���o��߼�i�C��jʆ��~�c��ʇ��38��m�W��'���%߿��Y����u:w�[�1��͕�|^��4�� �r�J��r
��25�c��ҏ#6 ��g�v�2z��M�\�;lfN �5\�YEIrߋl
@��H	�+m�g�0��e1�c�t���Ж�A��? ���݊qgt�tdA�j�c�4�δ�P�߾�@�ʨ������T��ѿ�{5i�%��~�?�w�|G^y�52Kkz�֤�Ӓ�٢��U�ԋ�vp(2���׿��[�s�*J63� ��m��e��5c�c_�"ǘ>>:��.{"`�$��X�(�&��^/Ї@{C�����e��4~�����n�5�1 ���@�Jl0+,*����a*��:.�K�0t��M�>+0Y���tA���=�l�GI\G�#*hYFֶ��:pi I�(p��=�dm�,e�������^K�rF�~jUn_�.Y[�O
��Fr�H�4�j�s>�H� �Q�3*͠/�$�D�P� ����f3s��eɍ[7e��@��Y�lsw_nlޕ���"���t�~�ʻr��5�B�ۺ�9�gt�/+���бJ��Ӏ�&zϸFp �LR&�����%�'�A(?}�)6�\'�
2������eia�jQ�K
J�\}���s�=���|ͨ��ONPF�EH�}8��H�&xv-P�t^��:oJ���I&�B���C
��� 4-�x�[��P�P�N�G<�ɠ'���7�����дS��M��(�����>{�<���g �=,�F����J��L�4�כ��bC}
�Ġ�����f�2gBF+��o�;��;���h�x���ײ�_7�I�r��p�i26'�9�w����R�Nz���M����C����d<f�(�5��?��j�0�1�5��EM?�R���39�2�,�`*� Ǝ7�?��_K�:+��g'u3ҵ�8��7o�z�Z��EńG��# ��x|��ޅ��n���޻���u����k�ݻ'��3/%~�[�%���657mT�v]7�y)Ȳ�X��'�M)����n�+I�Wc��n�U��~j^cꘙͬ ��d����d�s�����\<�Q�ʯ��<�|Q
�F��X�bN%0U׮�s� f(�����C�4Pi�5�7	}��àg�v}�؜�M5��ƺ_)qL���
S�}�E�I�$c~Fj��gd2�ibԄh�D``ҽ��\�d��� �}D��$�Q`�ـ^��"&���qW��?�[�{ҳb�C����òI�a���e��AN���")Tp+�����i��s4���dN?����;=�����',��V�K�*�P���~J�Ȃ�
�F��K �(�/5�F�,��ˏo_��6�"��	�tH(� 44x+��r�{B8�L�`�IA���G�P'K\�Z�mU�K�F!�8� �a�7�Gybxl�@��W�Ѓ7�����ҸSh�	}�Ȓ�RC�X[�������"�-sS�׈q�F�H�f�1)/P_��e�����+6%�G|��U����-�M8
v�l��+cu,�ےQߗ�?�����>/�̌�4�;_�H13��f�0�l�����ԡ����I�j!�lçE�ۗ�K��ߑ�aSP�+V�����3�����_\6���4f��n�PǶ9�ŋe"�;��l
@Z��eo�+ V���T�+ ���5�MC��]fd�� �ܴ�s������*� Զ��*h�t!�ۗ��m��G>*?�����i�:�Ԑ��?N���b��A�3���\  Il�(H��,��S�9�_�W6�'}&�4�B"�b�"EP z�����s�@��Bn#H�@U��7�C"`͌��cP2���lC��z���q�&^@�H�*,l>dp_�lc���ɌdR���q+���(��H�,f3����5f�i���*�ױ�ۓռ�~����1�D���Mސ<��:���]*�A����ֱߥ�@��ސ�j�������>k���i�:���#KF@�޿ٞ��T>>�j2{�o͂�)�n��Mb�Қs�c��F`"\�~m����{��Ͽ��o>�~�p< ��_����8!ϕ�K��cǺ��8c�}s�/�*u�����ǿ 7n�V$�]+�>s%��8�����%����P���̲������ln|HJE_>�|I�@�"f�{`�1�	�-�1pE��g��V8���7���F��B0`�1Ȧ���i�H`/\��s��E���Q��Г�	U�(+ �Qt��D�A1״y�5�Y�{Bz^9W�@n΅��pY�HH��@{��B�Rf�LUV�tꆎ`��-!W�ʡ3���]R��y�:��|~T>xo3����#:?+�?�� �-q�fЇ}�{�h�ZDe��zG�X�/oH�3�/}�P9�al/>~^ꍺ��~�P���~�K_�N�,���H[oMA��R�8P�(�!�Źĳ���	�Sf|3�H���+�nI�����Ӌ�X�J��@���P.Q��$I�tz�5؂*d�QW�F����O������H ��w����ڛT�b��+T]RO>|�q���ɒ�*!d�=��%ulf���Qg��M��N�܍��ޕ����*����	T^���,k�aG�5�l��� ��G�x���?fr^,SS���:}"@[����]�����=�!�������z!t��U)Z
�iN�1�!�Ch�/A�O���޾<��GĪ͉�:�S�JUjK�ro�)���9�=�����)��|��A��P$�IɈU@��.R���K��&g.,���� ʤ���6�ܖV�%oݸ"g�Xѹ�yO��H�Z���+���̨k��Ӷ���$�8Do$�+��OU�tm�c�?^��E�LĐv�� ���e/��y�&C�<��T��4��;FqbdfB��5IP̴F-L�W!.�����X邨jf�B�%�F24S�+���B���o&�<���P�����\���_PUc�C�b�ȾH�3�B	`۬�'�Xpn�|
}h&�=�z�mT��4u���{����;��0K�J�ӯ�>�T��'��<_v�*'�GHL����]��]j�)��m��u��g@�q���&3cq�2��e�bfϚ�*���$�N)�b2�f����;���֦��P'� ȣ�W����s���.�C���B�Q��Б�Z�n��q_����^���|��gLV9rd.�?�i���_a�'���/^������hh ���ȯ?�Y���to>�Qlh@l� �)}��[�_��W6���59�~��gE�����⽷��P�9!�X#�-T�P�Q8�^c�����64�3n�VNU`��ԝ�(_q�Av�	���Yl�+��A��s������C�`0�Ftd�Qm![��{:0|qM�=��	|n.4�-V�Y�FdR`ކ~�%��@Zn$}�D�ɍQ���b�i�uݱR= v$�Ih�Rv��4��B.�F)Gz`�e�z�B���JMz
�Ӥ��ѭT+|4�G����c��	�{E�O���m(y��Z��ew�y  ��IDAT����X�U7��b1ϰ��hl`�h���E.-��?��oɆΆ��0��E���Y�7���DLk�g�������$���X}U��q���)Q>�tQO�̙s
>

 l)%�$�)}�1ѣ������M���HP� ɁOޜ�yI?g1�Zi� >��w<I��W|���9�FO
l:Oy��3��8R��{.9$e�m^����z�m#ul�ڣ��Le���m�hȶ�����*:G�������uaiyM*�K�����mY�_�ų��I|��K'P�������1�k`���V`���	+U�P�L�"�5��e)���oTmY^=+���\��#vŗ�'��ޠ!�Kt�?��<���=1 �6A)*�S��z�����Ą�VF�^Yb�Rؓa{H#\$�h(��lC
w*`I���~�$j2�jC��7�z�$�Oü��؄5΃[z��#dރ�S[�8�9æu(~��1̥���8�tH�����:Fpc�� )fTuQ���T���b-/�F��y��D�����)
C��}���U4�8�8ԟB��d�S�a���~pO�)�t��LU���zeF�cZ��DyZ��k8�O���yx�<_��N;~�#jYvn�h���㴊�yL�ꁿ�f?B�������1����;�Q�w�޹�X���<�L ��S�G ���+}\�~%�qy�j����4,��:��]l;�=�~:��ΡLZϋ��Ǻ�!�E��1ˡO��r���XJ���xW>��'��\!�z�����h85k w��-��J��)2n76ok2'�Z���n��}>6
h�T��f�	�Z�R�"��]�"���4�
�BHie!�	A6�DC|7���+汧�*�A���i�H�W<(oɅ٨[����fw�����&c4�C�1A/Ő�'�1(wX�p�>X���{�.M.���T!��:��R`��B��ò��6 � ,�#�oZ1)P�
G:f>�2��x�sO>K���<��G^�D�{;
5f�4��aK���ގ��;K�}�<�ɠJ	ׇr��t@�lV�Q@D}3�&et��XPs8�Gf<!���(U����ٲH/���-i�z9��d��>�0���\`�x�5= �`�, �N�Z�*�'�*Հj�)�ɽv�A^N#�����Uuvn�9%�:@T���ST9K�?�C
��E�� �J�@Y� ����J�Y��Y���f�
�\ ��(E�%� � ;�-A�
��|?}�*~���$ϨCHa��!V¨`���%��̆��f�]T���"����5��x��9X<���M���^�T���-I7���/�W��٧����Y^�9�s��:����%��LeE������+��C�c�<F
�A�D�AIʋ
Nʲq�	��v{r�j��h�׊ ��RP}�2M�ñ���h	�c�a@���kJR��T�c|��grV7���ј�
�́QG�Xb &�7���  ��jc��@TQ�$Of�[��mc�dh��0� u*V-�ESd�����>61�` G&�m��`�k� �훞�Y�H
[�����\+�Ջ����&i�,��Ri�HbmB���jS41��|�������`O�����IǬ������8���w�,���H mM=�fAM`��'41��O'T,|9��@��1�`���L*"�[�W'�����L���-��Ǆ|�B5��3�G@�Lc�D�*������?dwqUq^�G��a��^�y�O��ƿ~�ҥ�<:N=�Gǯ�q��Z��H�xI�1���}6�=�$v�p�F9�`����oI��1ꯂ��P3��ʾ5�RiGCf�/�����2Ԉj�c3�o��`Pu�eK��z��<s�C��2.�>6��PZ;)]�7�-(#��$�p����?����Q�n�.@��4� �!���ܠ&�$A�~�&��������Ź�e��tt6�2�3%�a��p�I5�wo���i;�DF]��|�$\�m���U#C�|Ӭ�
�;�
���!���*M��#&p�EJFu�ͯ Ty��h<$��-�7C��J���[M����E/�P��)L=�;wnI}���h;n���\�a��ǲ��������^�����Ѹ ��%�Q4E ��� �VD��t��|���Wd��0��6)d����@�8�*�~��L.���^�˅��ʯ��T�u��
 T,��e
��z_jzN(0��J.��^��[�d��3>'\��������js�����(x>7k�|~�+�'�u�Ɵ�\�1�*��t{-}�P���xAB_�Z��C7T`�˂*\߽�m67��cSA"��/ץ
��В��Ͻ����+.�iB����ވ��r���0����u��+���~o,/��:��,�,�|Ke�١_P�*x+.Jq�*�nG�Gŵ��p��Y$E���
:�u����?��x�5Vh$���[g�Ґû[:�#�f`��)+u�rQ.�mpfh��k��M�,/�PF4�D�@�=�@FM����*�1T�@?������"�1cU�Z��$�&+�J��w��V=C�-��c��ɴY�-s�75#i �E!�p	^�=�^��5 �AZ&d���
_�{�0����#�Q��2*y�yoTW뵺d��,����d�1��+~�ºm� `�4Ũ�gr20�s
�}�������@/���X��4}����1�ˑN?�����;9H;�2�Ks�9f���p~;�N� p*7oM�lz�)�2�7�M��g�ƶg�v�����t�f���������&f�
���_#><h�������͸���G ���+�QzF�ı2�,)���c%���`�J���"($�P!)�j�@$R� :��aG��PbG��n��Q�cF�nbv̰1�9>��I������}�M�X<ԌaV8���Jo3��zݨ�:�#�Y�X���%������f���V���n��L�\��� :������N6��[f1��a1�bLR�Q�ױU��Z�������М]��M�'�k��=6M���Lu��Y[1M�P��GPY�hy� 2����FA�4�X� ���ؤ�#�n��S�t��qDP��k4�AT�o΅�>��~�����`Qe@pm2�FJ���g�*��H�cz���'���K���<�=���F͸��I]���;�7l�u&r��5V��	�>+hF_����loo�C���\ڶ�e�DI`�[i2Ɂ�A6b��P3bV�6����W�.ڤ��$HCV�u��sT��P��4��b%��iK��f ��|F�
0�����d"c+��x<�\�	DQ[���Ng_�;���E�u�����������	��|늼��w	@
բ,�.)0+����ܻrG�]�-��y6�ȭ«M�>�ul�2j*��aW޽}Ug��2�Pt�.���O>CWoT<}��~��>i�J_A�|u�����Ey��S|7=��z]y��;r�>��"�,��@������u�+�1�.	+{�$񚳄�qiu��W
\��;kK�RR�Xѵ�g0����/˷��J��P�����AM���?hG�B�8�@�2�'��8Hأ�=�Sđ�q�2�<HNC���r؞k$�C��X4��3(M6�/��f�2땘�	�A�0,l��S��%���q?�1�u�F>�
����>�|�l�g$�|�3��Ȩ_�ku������@�N�n�����D�����w�=��"9I���pR@|�a�����$��M	&�r�\�e�s�p���s���$�b���=��Ӫ@��ML�7�Ϻ���&����h�53 �x�)ڛ�	�7s����1��(�0qz�k��ך�=���`j��0�[�W�1��tEx< ��_��x����qdcc���k)@�m�+I5*�UY����y7��o~U�AG���4u�9+����F����cc�a�qƀ��r��bw�l��䓲��Fj ��ˍy��(T�����wI?��o�@�F����Z��a�E)8�T5���@;�(����eS��l���,��L�=�k���^�YЁ�'Y��Q�	��kbv������m^3�V冂��8�NA����r(oݼ"��,ʒ_���=+��~K��XEW�Qj2��r�F�`o��;��p���7�aSBo�S��lVR R�M��Fu/�����9���noJ��'�;���}9�ߖ(=��%YY[ˇ�2fz�/����ln��$e�4�c(�1 �8�f�q�P*b��mJ�T��K�o��[\� KOAP{БO}��?,��l޺#[��l�����1���ʪ�y�ft ����KG�,����0���͹�ҟ��P���Kl0&�P>G�~��A\n,��w/K�1k��؜�j5C���}��y9{���"���oI��-[�[r��S�MY_]��u��&���kbB�~�2'A�.�O�^[A�u��cok��;��T��t��7*��_�M�t�1�y��t|vw%��=��Oʒ^[w�����Gsc�T������
����w����i���z�c_�M"�	:q�8c0�6�HO���|35����/�7�����o��D|����W>�EY/4�Ur�<�	�<j�M\S���#���G�����t$,��H�P����s��T�~N$<Xa�g��(<���L0�,���C*:5�|��=@��R�=CX$l��ab�)QE��|=��P��=�
XH����4,[F��*~bhW�P��ZL��\�6#5�șAsrj:ا�)H�����P���:�X�.e.��X}񨈇Jh�q�5�
2dOn?^�8)���>�������S��IO��?�w�;�I}���O f�ي�,�j��ڠ����� �,��ח7v^=���������Î�Q��_�I�p��n�ۉ���ks�K�ۇ����� yt�jx˥���"*d�4
��Q�竛����ї�s��,R��Ɋn�_��/�g���'/�(�{��"�.cJ�rQ��P�4��g��,��B�{Qz���앟2��[��%`�ٞ_^�♉�R�����ٻ-�y�G�2��!���+-��4`p��xe_J�2�`��t�c:he�EL�E:!�:�{A&��_&k�F��B;�}��$��`�{���ԣ�L���7/HX��(a�����u�����?��?�qa���k/l�K�ߔ@��**�zE�BI?[wj@����l�M�Ya`��q�dM�D�`�T�@���W6��#q�`U���AkW[�r��5D�l�ݑ�8�J�,��fl�Č������Z��!0��{i&�'���f�!I��������s�+�I>1��rw��4�R.IQ����H����z� Y�3����ll�J]�	ԣṳ����נw�ln�0V�	�p/h��q,���l0���X��U0����x
��^�xIj�V��Ʒ?����\}���5f��Z���a`a��P�e�$+���9z�m�lI�tL �m���y�g��
�쒼������9Y��V��.[v�K�×�����ʕwޕ�~�A���^^����������|0*������P~r�u�>�șr�}1^�N{������z�>��C�>����ӌ*VI>���ȫ�ߣ?Ǚ�u�����~�
�W�%�m#^`�n�yr��� ��d��EO|=�q_�ٺ!?z�M(��#)蚄g����������G�3�ux�zG��$��0A<�;��H�Zi���g��|jR�񐢙�l�W*���� `TOQu�r�P���c;1ܔ�YI-��fR��#&�$E4M���e��P�d��G1�^GdLv@�b��r�h��+(�B�G�*�C�٠��'���o�|�{��s<x� �M�գ�5����e�\i~벣�cb���l��q�q�*ͯ̈���Y�,����s�����(� $,�-�2�f�I���C��U�`���<�F�����Fr��>����8�G�� ȣ�W�x���Ї����Y��G����.)i���6�2Uv�0�@��lfd%R��n_�0��DQ6��i��ԟ[2?� uj�}[n߽+������Ha�!W�I��U9�X��ڢ
�$��H�]y�������Z�	�~-��� �KW�B����O�A� ��W
��/Ȱ�5��\��[�2�##��,C.�6�2��g�5j:�ZLK��]2C�����nR��Msf��!��C�γ�����S�@��J�E�4�l+���~�'��a!�Wt,^�uE= 6����/GR�+;iJ��Ci
YQ8C9�����\�Y��ѐ�j �u�]���ź���ټה��~] g{������� 㩏=%�v��������c��F��[�\n8�����ld�)����iWd��������L��>����s��Miv�����RV����<�pVVk�2��Tq�w����S*���k
lWe���f�'���)~@ʋ�p_�k`]����̞R�`�&̚�e�&G���(�.�dkwS^~�g��O>/+�eV?z������P	��$��瞓�BC�ܹ-��&3���ZX9CZ�.��S�Y{Tr������i(X
R,��p��c"���H�ʂ>c���/������e����ɧ��g��_�ybկ�x�����_K�������
�{3�x��ė� ������{׮���.�W(�k��GaF �d�ϨV�o�2�x�\�8��Ϫ�U��ߘ`��� 1���5���]�1/\��1p ���$�P�VW�v`\۹)?x��ɻ
>�:�6|���>g>�sր� ���z�z�^���ox��LY:������2���1��q_S+6}=vB5,4�{�y'm&\ð����_�FM7Wd@��\
�gT��D�	����D*Yd���1 �	�^&#�y���
�P��nw �s�d��2c'����h<� \L�[�{��s��f�S���ې�U���>x��P~~��}��U��2���g�s��c��eN�= T�\�v�<'�����=�&S<���?�,������'*U"��;�8J)�VҜU0*)F���EN���(x[���9�Gǯ����W��ݺ5���%?I� d��d�&TXP]�ve�X��B4hc�I�X�x�U�|�m�����u|�/0+��9K7��C���}[�ݺcK���E*ͽ�=�r��|�k��$�x��`Ȓ����������~1fs;��0d���ۗ͢@�����),I�<2�q=����ب-�c�n�N$y���L(V�=�\ߧlMWM,��Qךh�m���j��P���a��&ɴQ������B�A�XlNQ�*5�G��Y]����\����h�6���A	,��)�%$�+	&�vU,�$�������N�����(7�S X���\�yM�
>�<�o�ߑ���O���A[��~��~�+�_��%�HI��U*~%0�+�i|$#��Ѩ��/�u}/�\&=��5�1613���k�逢��7������l�Y�O<�پrS��@�+��u�j�7ޑ��m�_���"+�K�0?'���,.�Wg̱R�j[*-CK�sK.A>��F��m��)�Ĥ��mm���\X�H0��o�?�����9�`�A�r��O���|�7~Mέ��흻���#3�f�E�אq��z ���Z���*Dz-́�t���t��r�΁���ݭ-Y]Y�?���B~���ʝ�[r�+��S�3��\�~Uڇ=i��+��]2��p0���e�����,��%* :���%�g���{�o��|��gu-�W���Tx��!��P��M嘛l�N�W��
�A�%��ُ� �*�����u����}��ɂ�[<ڸ��Ja��X:��S���F�Z�Ym���ԓ�w��m�?V��v���FID��(�ڄ`:ds�����t$-<�HP�@F�tM�4H��u���2<�afz ��И��BcJ\;hh
��N�)`ad�	�λ�t6(��Q�@s��ӯ�~U�3����ޛY�_��.�޷/�r���ڷ��V�Z���D��Ad@�[�f�b�`��CG����F�3C�B��jm��j-��Vwu�յ�R��}�����;�{3_feU�����ۑ]��w�]~��;�9��>Q��X�]�[=�R�C�=k��&��;����(a$P�����|>^� w�' E�}q|��Q�f�(h��ёό��UH�K&�P�]���RUG�p� YQ���9x����{+��T��,/��P �A�4���½�����`#��U�v���1���x��l�)�hCx:�ϓ��ȑ�h��d�:ޯ��j�������#�����v�}��T6��;��֗���O �׸ ���u�9��Z��sf�T*�
S�a�$��rp�r�s�_�����[f�����ЄU��9���p�%
RJ��S�F�k��2ȴ��=��IZ�p�q�>��	z�[�FY8��_��i�ߥ?��'���
�YK�xo8]Zs���ɵ#r-%?	E'�fN�!�$l���AOe�xe��08�vQi�;�H���hЖi�P|� �C�V�'��#M��N&K�3L .a0(U�PQ�4EC���D&*��>ЬM⌭+J	LI�O3���B?�+S���4��x&C�v�jA����!@��:������`���+W"���mj����zG���`0�C�H�RH1��*� h2�=�\�����!����2�?�� ���A^��ҕ�+���hjl�
FU2�+�MZԨ���/�T��x�K�O�#�w��R�R�S�Pk`6X��h��߮ߡ���sM��9�^���r���e����r��%Ps4?5/<vP� �xk���!��LӉ�g8�]��R�=�3:�����
�1�9��}��?#�#�����#m��Y���8� ��X٤�}�2Ξ{����P�����,�\�㧎����)O���l
��glɐKR��Y�ߛ5�
�3cҩ�iZ��2M�9�������xsC��s��Q�R������Ng�?������MOU���k_y^L�<ǣlF�14��A�Ё������	Db[���ק��&]X�)�!��'�v)M�����S�_��#g��Ѣ�L��nܤ[��0��6��3df=�& �[#���/�ֿ��} P�?Fc�O���:M�%:}�}�gD��b64�f��ߟ��!LR�����'*t ���/x�A�X.��k��j�+�RZ|���1Β��,*y~ �Si=/bx��Ɣ2 ��.�M�К �M�z����~VJE���������I��&�|�Ri�҅�<7�B�c0�/�
�b{�iƔO0�G����� Y.�A$_�zӆV�ǾJN�O��CRq�����B�LM��Nxgv�wm��o��j%X�p�{����ma���V����O�G�ڡ^��Q
���~����$Ҿ�����_e�~[rI5g�u��m:����=��~��k�߮�Pij=��:���ƍ����>��λ��n��׼ ���u�ٶ�3� ����[y^��_:*./L�{kԼX�G~���"�\Z�Ɓf�Bp�[�nlq�<NO��BQx��u��N���*Mq��S��ѻ��.��p`�9���2���o���]�5y��<���R!�<�1��M��h�!:���R�⨭��I��	2yE�m�fRP*����ŉY�ê�l�_=��e�ӌ�E��f�L�2֤�[��*������l��E�WF_�t��R���!��8���-Lл{-d*�fЦ����P����ǀg<�b/ρ�+���n���f(�z *�$�9�-ezl���}�ϋAKƔ��	��X&��C�|F���'���r�F��'h��u�Au8�P�q%�A��|2�+2���"��'��@�y=Z���F��%	 Ã42�(��J�G �%�R�J�� �ʁv�3i���\qPil~�����8���i*?��2E�f�R1S ;��KC���#8>{�P���R�"j`�q�w�!&{^ԑ^���X� n�}�G x�0��y̿�7�٣����[�0{�RpC���  ��`��>�\)�	�>�G}�>�я�u4D~cPd���O��62C��|���
�Eۢx�w��_�GN��'Ϟ�`٠G�=BF�*S���P1��'N��ğe|�A�;��W�R���(�n+�F��_���u�
��zE\������u0��@��
�	�����)k<#4��2��W�����T��R;�㦏k�6���sחgD���/2������I���j-��G<��<N�M=AK~��\]z�|{!�?H2�TSK�4�����5`2}ɗ�yT�b���U+�fx�@��������9g4z��@�ܠ	��x��*&� �uT��<����۴͙�Ctwy��1�%EEzYl��*ay�w��$�O�ճԽ!؊*zo`~�*��+�Q��O�z)���8|�'�^�w�F��S�~��wB�/@�$E����47'f}D��P�i4���Qy����U��gB��A�;|��D������v���@�m)�_�]u�n���{������^�L�����"�v8���GD}���K�x���� #!�9/-�ը�c�u�}>{{B@�[`���ޥ�H�u/
�F?*�������f����w���:l��v @���f��I�'?���`DY!Ra�7�D��@��iҿ���IG'	_�lQ�� �=�����yJs�lѹG�᱇�����o���}��_��������)���9|��7��_�/�^����R��r�Q\���G�@���D�&��[k���� ��Ga��ţ�y��g��K��=դI O�I
ږo�d���(���E����xj��v�%O�F^��ƫ�'�~�uh^�����4���yzCy��|:E�L^�ɷ��LV�􆅳�y��*M�+w)�����$�9�I�p��@p�9�(={�y�}�b΁�Q�A���b��Az�!�v/����K담��ʆ���OT��l��̕�G/.�Lx�ى�;=���]���b�@��������=sG�_�������*���gT>�t���c����W�YE�j�@|�i��o{'=q�^Z���49GLB�R��*��Ġ.���QM���)Z�Z�N=���oS����7��}ȁ_mm�����u:;w����;%�玝� J]T@f�f$[�{tdf�n/�R�ӥ�O�FC��[$R���ړfg@���V�N3V�l�&�Uz���h�8NT���ﵡl�*s˥��m ~@��r�3��ѵ$H !�
���sD��Ҡח���YU;�4@�Y� E�ѐ}@U�_�B.�cϓ�����ɇ�Hv�L���|����qa�훟'�j�A���eP��pF7x��iX6i���j*Z|�;���w}�q�uE?B�R�8>H|�q�m(%:=�3m
��@�H����!>"G� Ů#S�R�
œ�� ��ͱ�˓��я�4BO���2�I� $��ē
j�����z$�*�m��T�\�tƒ����:��9ُ)=U�R)#��*aD�'#�� �F��M��D�gc������@�	rlVJ
���TRH ��mA�D���\elC�;���XUK�;H5qڽ�co�]���4�'�����j�ޮ.�@Dۯ����ⲇ���1v� ��u9ϑ=�p��� 	]�k�Q��w�?��7QǒP�b ���܏v�l�xp��~>*����w���뙨�	]-N�|��yˌ��Pd����V����z�����o�گ�@۷� ���u��z��XY�
��k�@�7�}	�H&/����uڼ�AU��Z�R�N�����;h.;A�.ߦ�z��}� l
���4���lu��Z��|�	�ugI}1i����焯}���R����˟Wh� &�b��Z�A���x��\g
�p�-��y��h���y��Oٴd'C Hz�~rҤ.�P����G�^%�M��	'L��cꐼWe�%�A��R^�<� d,#�^Ie)r@��rj.C>�/�B��u8�G�ns�t��1D ���m���qj�$ӄ��Z�Pnv���,�N���)�Ҝ���m��m���ؙ1��S�4p@����� c0��r�03dp���ݧ��-1  E�kq`���ӌ8�����rO��Q�6H�"��ɮۣՍUu�p�)��y>m���C�ʄ@J�*��w�h����E�H�����m  @s��|.pFo4����fp]��I_|SP�@�G�����A.�@���V�P���>B)H�������T8*�����C�͟53{H�Q*�̴k��G�@YHh�M6��8 �T �Z�}���F��|Nyf��I)r �̯�_Gd��l������J��]������vib�@���� E����z�v����e52PRѺ!���G9<�@�"�7x��Dh:d�h��ީ7�җ� ���&��!d^9o��0u��̡�T������rB�
��C�=��?�@�HY�2Ie"/l�UE�y�S~ ����@5
�ڨ^D
�R�,3XF�/�Y���C�/�wL�TC��|͡(711A/��2�ݾ�8�~�%���� �Phyq �A\�E�sD$@D3����L��,?;���lb*�`�������\k8��3��_q=��&}l��3�B �[T�M�
\J�,i��נ�����҇� �I�а_?Ƀ�gG_��N����}SiX艴����>�dS
�`�+�ڶ��Wy+T4`�
��k��7U�����c���v۟%>9�ޥ@��b��1��-���I�ǳs��������)���`�+m �`{]oao~�M���a�p+�C1~�r>����#��zhR�kRj��{�#t�X$o�F����k7)J������F�:x]�t��.-��W9_ð�VK&˱r��X8C�a�>u�˴<�Sh@1ɡAAKWj����_�QI�xɤ�E6h����{arJ;���B�l��j�Y>�p���MXdщ�IՈ?� �(cJ�?Jt�c>�d�R�1W3#D��T�sP[p���dy���h�(�����@.���[5�7h��Ż����^ R����ߵ�_�
�p���-:<1+N�!�]�Ǣ���#�b��u�t����m�����G���VT94�=��-A|Z�K&��l�&�U�2�iZc��`���
�ߓ
BG@+��џ�^�<P��[kT�d����]i���Uv��3{�̺P��$��Sϐ��a���~�+��@�M��I/w�f�\�0e��d����r�h4T�aFi�+py���-��B�N�lF$_sfZ�5�Pus�4Ԥ/!͠�p�F��c�9���:Mg)�)PA d���it��3����A��\1�$jy��3���HH�V]��|N�_�ZR=�<�H�{.�G��R�+d@���tim�I�N��?��l��;Q��C���p�++KtV�U:q�$m6ڒ��g�D�	_�����$ 9Z/��B�p2S��Z�0�����<7 i����G�l^��X:�}�����P�������t%?�Z$
 r���f8��)�V�>0���q( �G�F6�syR1�<^�%��¼���<�ܢy�T��PhC��� T7UD��
���P��@D��b�2%�>���1�@�ǾBb�ȯ�ad�c<'��h 9h�7=~�Pu�r4;=Cy~ާ�y����3�
�@6CBM2ў<G(�8�@U|0GJ&S�0�C���|�eŠTьT
�I� �� ��e\�5}߀�~��������^����_�u��}zO�w��%��	`��6��x��������V;������Ⱦ�ݯ�GT��bFa�_�e�N~�����/_�/W.\���گ������r��� �����`8��3&/(�mYal���0�B&�����8X���D:C�Dd76i��R�x����Ŵ�q�X��B�ƫpPf��T)V��nK�ԫ�V��.�B�f�ez��9�ڵo�Zw�G ��R���v�W�(��7$S/CI��� ����A:/�h�T�ފ���4���F�P)d�[�^sw�ʏ�(vx	LeT(2��K�*�A9�x"�H*5|� �̺���pZ�wk��3��3g$h���?O�k5Z^��m���RgHw�RU$>��ZN�M�׸\�V�� �S��h�d�7+4�-�f�20Jp�q`:^*��״�lq�ڡ��Y��"��|�u��9^���8�/��T�񹹹E��.�V�N�}  ;IJk�:�����M�K�K���*�ȦI/�(])	�DY��0�S��t(Ɛ�Pw2Xy�A�������a:2s�ľ��%�� S�*ԩS'��ˁz	t���ǔ��9~Tz+�"9Э��F�!wȀ�ȓ��hxrZ�1�`��78��SY����o�_t��^�s<��b=`��x�  ��l�����{�*��.R��Ȁ�ʈ>%�w���j��U��{��r(�sb�3T*�_�}����K�<�A��R��DB�A"zD݋�͇9O'Ξ٥�<,[���8EV|��=B=J��[7�tE	C�Mܠ�
��B͂�kğ��gU����fT���g��W�j�)gx^�ȸ�ؼJ||�ӹ4���F(ir����e���J%��7p}A,s+U��l	��s���01���Ic`PI���7��؋!b���ԯ�I%$7�y��jTj���U�-�/�V��^Y[�Ǧ#�:;=Gox�Q�1�t��0������/tB�*K��D;p조��_|s�JUJ#���b�y�<��|.C�T������#2���3�x�v(DJeI�몶pW��7x�o�_��~���MQ���������@���i1���	Р�����w��؏��UR�y�q휣����?���Py�nWoDX%�G>c��qg^�pa}ei�?��������v @�����͛7�ه����J;e� �@�����W����~<[�9;�AD�fx�8��ŭ5%(5�4��i�!kɁ�Ap�+cdg��I7n� �P��w���T@N�u|�Tby�ȧX�V�@�.�QL�G��:]�l���i��D�4��Ah?���<P�*������H��ʈK��<��T}��ǝ�)UAj��]LIo���РA G�4��S⫐"���_�;�n���<-/����3T���_S;W�>Ȩ �8-�t��!ɚ�d����5}Z����h� �iҬ*�2���q����ؘ %�P��f)>GK� :|����4�|�<*�@�)��hh�4�(r�� F��>?�W���X
�!�O�d���%��������:l�X��I�L�r|n�S3t��K��:���/��ݻ�rc�^�p��)~�4`�}�r�e�w�e���$\{�Us-�i�";�q?�HG�C=C�=��H�[hss�=K�W�n���;|Z6�O�J����!����;�p�(�9�^^Z�/����m��;4� ã�
�4H{d�5F�0�G�\�J�N���^NL>E��GԠ�A[��4�9�x|pȤ幝᱔�fhu}U�%0�h��F��8H�@����$K� �:���*^y(�WS�[�
oK*~�������G�{�`2� ��h����PG��`�B"��� ��1	u�\7�� P5	����s��Ѻ��`��~�V�Tc�6P Q��tTbj����� $@e�+����k�J�� �#���
�ʮ��<���G*�C����K?�8�C��@�q��q������$_W�;���◿DY~��EWU�4~_
^%��z,�����#��`��Q��!-7�+�M L��%��GA��
TR�5���uW��Sz���o�޳�Ha�>��? �O��kْjŃ �~y��#{��o��C�ۓc�J6#QA���|��}�4��_A�o����{���1	G��I.��~dq��[]���KW�\�b�4~���@n��� ���u����^ۤ0Q��d�A899A��ڐ��3�,��#�k�T,ThRK�7Ao��qd���6<���To����#�k�'˒6
4^W��o,+�/L����i1���D�~���Z�*�(����IYde}����`��K�(���VZ5�#�
�Bp�ѓ��)L�r�al@�&O�����9%�l���&�zX��A�3N-[b�gJd�� ��^H�����&r��J��.��0nM'e��D���G�H)|8%�2%hB�?^�P�ԴeK@����{/�A�Om�%� x@VԏA_H�҄�kѬ��Ͷ�z��}@PU:m��Ǿ��=Ns���/-]��>�����&%Y�H�ɒ����C��]*C�KSav�����r27��2�Iw�ݢ\��U�JE@r����9�}��!E�k4�|+R *��H5��y��mJ1�ɕ��q���A`�n;��p��H	�~��ڋ�(��D���퍍5~6\�����SH�S�ۧO=�)���?M��?�ӧ��?���%�~��066#��p�?�!�<A<C�{��+t� ���τ1�����?|?ML�����#�1����9��0P�؟��a�" %�7 �>�g�5	���
"�zd(ք�m7���MI�K?O��ը���J �}��iP�9�����U<���y4Tkw��9���G��c0�c����7��;H
x����8W�� [D��)]�7�]�ו�'� ������TMш,ɃH�'4TC���^����m�+�H<���*�Td��+R�A\�纩�=x�̴�<5�BJ0O@�VÑP��%��A׃�����ߥ7��q酺��*�-	E�]� ��O�g(������8�HS�k�ш�&��)J$u�� �U�6�*n����Zj/T�8�c5'��G7@�j�����ER������]���� >ڳ�D�|t���1��W���D�~���Ɂ�m��y'�&�v�awUI�oD�T�ln�իԱ�TF?g��b��=���63/��U���;���;oܼ^�r�������o��G�_{;  ��z+
?�A*�J�<77��l�<���r���#���c��|��˓T�9��4J���n��Bf��S6��9#��jU���H<�,�R�����5z*�s�o)^9�Q������O���h��q�	���2�����_�̺TO ��iq��U9��9-�/�1��%7=��(?]ek�v!S;h@g;��c�h)�1$AE� dy!�,�vS�L����@Q��b�.R!UJO![+[ZPq�H�.�G�R�A�=	��� 8� afrF2�)��"�w�矖 Ϡ��iZ�����oݖ`}0�D�Z�����g����@T���c5ȟ�Q�A���;�9�)����q��W�����8���|u��d�2�p0DY�?�9�C�@8�t?��[|̚P�S�L6y��J�:��4ֶ��:��|I*oA��f@�3��7Yc���Ĵ��2�Ęm4ZR�@}�s7BMh>�n���d�.������P�e d�����8���������3������
�����cǎҝ�%*��1�h4c���8�
*����kw��ؐ�����`mc�"���2� b\��!P06>)�J>_��nߡ~�� �-�	x��}�/h��]{�����@��Y�Ko� Uz��!0N3���C���L3,��1�w=._;;��c��H�f��@J$�����er��(��cP��m*���ΐ������e���Lv\d�sZ��� &E��MSh�g �e�\�E�R�T@�J	K�m�Hzs���u%�����_d�1�al
Ε��/��,�*��r�T?(N~@,�r�.����[r�T@,���R�m�y���c�fq[(��8�K��̌�(S|����s����45=��\�n�' Ǝ����1QY"UAH\�q=t����PT�$a�<����#)Ћ ӌ�LJEX���_C�g�h�c��^�� �(�G�����~�U�8��n��T;�n�U�>��Ozw?`��}rM��ӡ���A�h|`���@�Oa�A���$�׶"Y�� Tt$RZ��ҭ[w�,^����7� ���u�uڝ���0����8��	�݄p��2yhvt\*XD7:���:����'�9X3)Hy"׉����d�'����Au(+�p�4	�XqH]��3�zwYdN�/�V�h�g{�T����0��dPJ�h�Y	�ν�a �:��hq����֠LDJ�2i �I��jP	�";�J}�� ����$�TCu�<��;�>ä1��H�;�4 �N���&'�%�/|{��?�	h7�����t��I����	\�r�2`���k� * �*�Կs���m�A��pR�B��2��U����]��xJ0�7a2]��fSI���LuX&���\��Erܮ�H�BY*�+F��՞��x���EN�d8M���5�o�]'jqP8T�qPSp��R�:�MBS��' O�;�Ka0r0�˚�����pxAw���ߤ��w�
��u�4/� 7ybv��Սu�כ����DvU���M�I �خom�z؉��H�c� S�^w@��_~����?F��_�<�9}Z(�<=z���7�&
U�7Ըf+cr�'''�_�r�\>yq�v�bpC?�NMN�R��� ��)��p��Ї>D��� ��G�����ťc{��n�^����~�c����Q�왙����+�y&?���N�@�H�����``��6���9]S�L�~�&�|�����,�l+
�h?�ER8��o��*U�*2ln�i��&�iP����gy���#���BS���E(��I�r�7h��Si��А�c��ʘ�X-T=*<Ζ��{�#\3��
��2����2���g�N��=�:{�A	�x���iiJy:�}J��9��ZR!��
��; Z�s�/=V��Q�O��G��Cއ��K@$��S�'���_ �3��<�b|�Ѭ����{�`5��1}>H<�z��@`�TRB�d�*�"�6����
I��f����I<�z��C���w����l;A��N���Q��4h����lIe ����봧"!�eax����UEr7�ئ0i�ߧ�գ�0?��s�'ǽ���h�Ғ\'}��_�W%�E�י=�_	��ި��^����6���:�_�d25:��ƶ r����n��[��ŁM�[ah��i�-tT�X���~�4�C����8t��}PABˉ�85F��������%����i�T!O���ٶIk�5�]��٩m�T�4@BT�=.`��fQ4�Ɠ{�d`�mwds�![�CYI�N�1�JAf�(��2gZ�T������c�P���̟�c�s��q�ڍ��G�)�.�KS�/�3�*��H,�J	2��t��A�Dy�� ��)�g���M�8.d���^�͠�C7n\�JhfsD*Ȣr� Hڊų�T�q��+w�.����JUB]Ҕĭ�;��R- ��@T²yQ��Z"��x@P�������s���[�U�J��0ޟߏM��� Ѥ>ϸFC�/����%�w�����u=��kT��'����9� ��P2�A���g�?�SB/�v;���Qk����*�iZ>�^�/�ࠬ��2�u�e�5ġ:	�$
�U=<�.����h5��g>A���w�c�=F_�˿�����������w��R���&�D���.襗/���S�op�A��+���zV4�_�A�ÕĿ8x|lnܕ ;���/���J�¸4��b�ݩ�)%����Aç?���s����!z�w<����8)*��'z \������!z���Tʓ�1�v8#���@�*I?�(α�R���)�/|WzEp>�A�����8xR*\�����*6����0�4�Ƞ��s�噆�W$�CȓB��^��e-�����G��4�C_*�����$�EUk�4E����eL��E�J��n Բ�z��֐�F�Z�5���P�<~�0�Q�A�[��-;*$����35��uL��p�N	0F��P-�8�ۯ�RB�()q1w� <{�A�ڟ���]��$��u���) 54�+��H�D!�,��|�LBS��{��	�π��ތD�v�{(R�4|���<y���'�a/h���F�{h`����#EqP�}Nbv�C���h��(�H�v%�0�Q ��NU���s�����G�����/>hK>K���� �JD�_��D�4�")��̕�����^����>��-�_'���W� �����CNLMv5-J��kBz��!^�̰�?\GvW�O&'��[0??O����$ά�{���ʔ/��//]��V��W_�E��cG��DzB
Yq0C`?>>�DM�;��)Z���B� �ԬmUJ�$�)޾d��F9�j(�4��B�O�ZM�놭2�iMU �l%�?$i�}P�Asg
���|[S4/���3հ�Ǚ-?�?ȑ�	A���cA�eQF��X/��A��BN��)M~�z�TM�F�6�T�^�hs�T$@���p����8*KZ|�X@:���%�?l)�M?p0�l�I�z����/G8~ܯ��\�U���$#zz@U�RY.�i���1�v?�)�L>T��ss����@� �Y������e��
��K�1����G�����Ӵ��F��zI��y6���:��g����ܤ�~�N�8M�y�{�7���:6��TӻR5Ӥ���=�j���,�2�,���N�/�d�A���?�8=~�~���~�}2To��?����>��/�jWA#���2=#�)��ǅ8U]�9�F��'�>*o|9��"��KSSmZ�ri�Z��[�f�/�[ss�x��=�*E:u����"�ǳ;=;�m\`����;P�6�>M�UZ(MP� ��'rɨ+ꍈ@M�����w�P��J����@����\�ɔ�P�m$.�4���Y�vLq4t!ZZ�(s��'���Ѩ�H�����%O��L���2�Ǧ�!;��J�.�<��D����ٴi���0p�\Zg�~���Q���#��o��ƈ����8���j|R����$�,P�r��>y�>M�O+��QM�����
�&���y�\��%�c`��nE��d��@ha��P��W2���+�W�>�ˊ{D�u��򘃬�s��L�(a<�L���{��0��Ѯh�qi���>���H�����m��]��=�{ۯ�n�]9�#iﯷAƞ?��۱�)<yoBY���[Iy�m�j�Ʈ��|���z�n����$w��8�i\����Q���C���f�<x\o�o����?��c�>�����}.����� ������˦��#���f�,cj�5�VhB*�sD��xhhB;J���<��H�,�k��;Լr���^X�E�>hX�E��}�k�;4Q���z�w�����2�9؜c ��!upJNS���jk��\L�PsAI>�i�$�j����I�J1��x�N��J�p�(괡�)�����|�V��lg��;�C_ѻ��cm~%�'���u�q��)�d�y�<Po�(g�)wt^8�"
Pf�<8࢟�!��q�vJ�F��ײ���M�ӡn7MKK�T��S>��#�*�=轩���Φ��n(� �o�T�0�T ��e�~1/ZH���"����|Mу�*#�PX\04�u�����cG�>��G�C�ԋ�q@�I�~B�K>Z~�!�o5���±�&���[���=�M�-�Amћ���qp�)�J�*���'>)A�X� �=�������P�u$s'fZP�d�����Tb�6x��:��R��CM�1(Ua4����l�B���?KO=���]���A`��	:ʠ���}�ҋ�Qۢ���������;D���8W�&�|�C��3E G�.��١j��>�A8��t���ei^X8&�+�6���}�hvvN2騔}�3����)���Y0`�K����~Ђ@��G�Tt0 p����}�8�h�&o ��@d\��A���}-m��]5g "���'}Е ��u;=����9�/&�c�Ξ}H@�T;����3 �\.#�Wu>�T:C��I�`F��p�:.2Y~?�Dq�N��2����P�|�@D������D4X�$g�N��M�
f�
ٴ����
R0��1�h�;A?��RQYߪQ���TƢ��x��2���#�A{�'d��r�_���S�F%����Dʉ}t�	}'����	T0�L��T�F�Hy�QLU�
���ܪ
al��%,� �J�U�91G�X���6�6W>�i����_/�= $��$��W1��~��c���~�����V�]�{��1������{�j����<�x�D"��s��u�@<�굫<e�>�S�2�h>����W� 9�^����tp��)�~����<Y��+�w��7�I�u(�z�ҭ�5Z�Z�f�CC^��7k��d�x��ʍ��J�N 	����$l�Nq���5z��_#غ��e��P5'�9���4(7�ѭ+����FT��О��-&�2�i�l_諉�'��2�0X���B'�`]i�#+	�E�Hz!ܸJ�d@�# �~ �Ӳ���R���d�Ex(����ڃ�������E�#���6-/��{����.�D��k��u(�&k�]V����	�@���P̉jO:k�bS�W��_�.6z&��12QY	X
�
�{ O*N��v��	>,eq=���&��>���E�ԣ�}0GCӭ��O����9:�f��\^�:�1A��y$�����DhVg`5�v%+��Iձ�? ]p��t��M�h��9v��tT1ҩ��H�����n�R��8-�q�IF���������<�z����x_����������u�Ќ ��?��x���G�����ibb��?r��v�����-=FSS3|8H��� �CK�6_�vf�|��,S�D[�W(nx�L-�)����$?ˇ�	��l0�)ѻ��.q��y�'��3:|��������bf�P��=�`S�,�0��5����d�lΜ8!B W/\��G����H/3���x�k������'
pxN�@�xK��I d��OJ(y���Be:��c����n���rA��.nmR!cӟ~�O)�e X*�f[���.c�����__4]�C��
Y�,J�EW�O Ɓ�dm�:�P���_�ۛ�x�M�ʞM�L9�k�gƊ�	?�+ĕ@�{Ug`�pt�P�צ���-�&�<����(�O˳h�Q��W�"��s�&�O����*~����b5Q���Fu$9��Q�C��D-	�&r�J,^;�ָ�6�=����$@��#��#�G\݊hw@�|��BE
�]��*�U�~B��8�1����k�_��ݒ�>�w=�8�#��4$�(��������w�����c�쾀'��H�������(�M~��%�(�M�'8-�JY`t��������}�~�A^k� 9�^כ;2��Q�Mò����cIc�^z@��O�\��nmlЗ/] ��l�!sjCR����l�P��)�5�	�|t���e��t�Ñ���<�wp��#�_w��r!�o���4Ur0#@+~�bС+
B%us��*9I�m��ׅ�[98	�.���Ȕ��d�b:��,P�O�G���&�Q�r��s��Ǩ��ØGJ�C��"3�d)-�RX�����U�:�uk�͎S�AW�� �ۡZ�Ff�I/]y�VW��~^�j5� j��}ɐ�A���C���!��2�:�ZT�nR� �Ժ�Y;�P�4�}�΃K��>��oۆ�P ��~W4	<�~�����9�"��g��Fm���P�?�B�K3H%���CҡA���9�$������!��n�#.hd5�/G�^����}�/�s��]oQ��U�z$����.���TN��! �\_�β+����� �X�,�gQ��*;���(pH��b08�B֣\.M�n��V�A'x,<�'�mo{;n_*�rԚM��׿.�hjf��ϋ?��H��#9�&�'�v���ȃ��)��Z�.gأ�zM@L��.d��_�F[�u:C W��l.C3ss���DBY�@��(W��-Rk�_��!G�L��|�p��a8^y�80༹�L�ަ���Y��!��;�N����Y��<�猞#d�''�$��g|�_����^�s�T�R�X��.ɊB� �����X�K�U۠��*�>w�>��)7Q�2���?���ށԴ- �
y?�<)ee{�+���Q~,G��%Ji<�y�!���{��#Xi�w�N3Z�����x}t]��*�)�J��kzJέ��� �~1���`mk��w��+d(;Y���D!L%E�o	*6σ~�=OU�¸��O�U��GY�����Ti%#�͸Ï�B�c%�T6���D��}@�JAM�e�?"�DC*0��DO�5G׷=.T�g��{�����D1T�����ﳿ��%� 췽�j�^ ŕ�W;�o��VN��(�k��c�w�T?�)[{�f�%xGzrHK(oda�������r��+7?���-��,����� �l��-е0�eo�6D�w����/R��;Pl2x��ȋv����(�gP����_�Z���Ac�&G�O)yZ<��/uj��Iui�c�#Ǐ��;K�+������7�L^FC,�d���'C�9��]�!�iSS_Am7>*����d�������0`
bs�� q�P^(�f��!Y<��ŬLQ�� $tu8Q\ �c��@�Ǡ^����!]��t��<��9�l�H��h�������96�3xi��d�[a��>N��2e�	�;B�
e
�8����P��B}}���"U���,��aSs���18:0��W���%��r�f�4]����r�D�pF|�{���-�W�Q׏\�R>��	2�u�!�8u���=M׷�ҝ�����h�Gy�V-P�L������Z(��1�L��{�Ǡؠ�ץ��Lc0��̐,����鍏��.]�D=���X�Z�2xEc��ܬ�^�e�^�9��� �ȋ�x1-%�`e�8��~����?�A�Ϟ�gB�v�)[d����\��^��?��$/c�k�CS�� 6��I󽫤j��H�>�_ �נ�*��#��q3;w�ߗ	��gN+sj#��1���A����$����%}� .��X�79� �:��#Hn��)[��/�H9ISc�I�g�\*K�z[f��%pF� 6T\~�~��|ݼ}�~�W����У�>LO����������?����m����������
�1��ұ�#�<GG�,��gpRNM�1+�ɨ$�?���P��Q��5*/���FE|��j�)MY����&on�<����$�MQsqU�v@¹R�gj@V)��#/@E��<�9���,��L	`�hm	���@�.2ȷ�j�R���<A��J�6\B7��Ja[S	-��b�$�27&�\C�M�5Td>C&rW�/�7���՗1l�J����1U�S$��j!�i��`S�X���ecw��R�x�kU��O�>�o��$���a�	����؟�u�����G;UTu�Ԛ!��H�d�uռ��s����,�&��p�{^�x,�<��������p�ٗ�����G:��V� r����Ӥ������G�6�z*~��寧仉g����#�k��Z���xs}���./�y������'2a>S&�´T��</8��w�>]��h,��x6%�6}���v��O�:
�T\2FFi�̠��*�
�jM�_X���$}�N��&e<���(�s���J2�|K��m��$tL�Bs�L����m�.~"�h�	<1u�V �e�F$�X�V�ǰT3<2e(b
�]��n{�"�h�-=d��ӡ��]�iMS�?���L����8�2��4�>t��SF$2ш
׍;W���-Q>��c4V�.�w�t��D�]}��z]"�շ@�S�
Ɍ�R�A�	�d��d����K�HgP�����m�$�F���`����Wc�akHf��{�~�Q*LVi:?N�����s�T���{s��E��E�F���!t�Be+�W�8p�{��r|S���ԃ��ӹs����/����X�H��ڍkqӥ!U8��F�*E$�,�!�G�����u�N����k7�«�k��~��T�T����v��253C����3���?Nû�R����|3F`U!�+T�.>���eQ���s��������L ����&h|��:���h|r����bC�������4��#q���Y��t��y�ES� 1=V�K��{����*k&e��e+KsPK�m���s��f�r|�L>�ַБc���+����S�#?�c�����������F�t:G33��왇��˗�:�*���� �!�p��<}�?�|�>y��~�ez�۟��;��O�?��,*)�@�5@%�Qf�����`0�|Y�Y�7.�B3~��M��#��Hy����w�d��Ʃ�����{3�@}n��Z��ؤ<ϑ��P�䶺M��Ar)=YܑpEH�;_(��c��O�U�/�#S��*(f��ʪ«%�L�����P�QF)Q�-�q�DD"�y�U�zK�%]�6�W�e���; CL��h�����ھ��^0�Ю��&�E��%�l��2�W}��k��c�=�!{?�AjW�}B1���)P�4ߣ+S���WRw9��Id��h�d��v��-R�Z���uH���'.���Zd|� |��l �oy{ꩧ��rz��I���7���-.�~�Xu����'
�zSw���͗^��������~�>p�:��B�'Z\�P=C�pmm���(��r2�nm�2�A���X�R��K��wz�����$/غ���D�8.����Fl���mn������1����pB��bͨg�V��#����P���ڪ��TC��=�5�M���/�
�uh[)}�fSd�x�ն|�|��넥R�/��Q�ن'�����z�c�0t��:O�Q���)sc~~~-�I�n^���'tn-e�휽<��������C���|ޛ-M������spn�|�2}�3�dh!:���,�T �T��R�?9�,O�v�.��@�����W�C4[���X�&�B9O�l�V���%��
��Z���%j�Ri�\ТD�7hPwd1/�@U$�quaG_U;�%Q��=
=I�X\(C2�aO~�@���z3D��y�yU$vUv��Cq���AqN8<	HQ��`��	���\5�@��6�k�Ik�Df����x1&�n.�хSth��ܖ��n���6�O-�?�Fס�́��P�ޣ�v�Vz5��ݤ-��=�̑�O�ߗ��
@alf80�p �������D�<��շ6h��mZ��� sK��U:˕�P�@aC S�p�{�ML�d�ye��J���uzB�3���&$��z&YFYkS5�>�)#>\s=�i��U� ���]ߡ�v&k����`������O�����ѣr_�����}�K_RjI����3��9��z,���\��h��]�)|~�^���������������fz�?� esQ�2c�*���}/�o����sg��ܴ*���c�L.~���<#ǈ>#1��z:��rVz\�T<t��U'��ۯЕ�W��t�p�3��d�...R�������d@!J��`C�<���!��- Y���5y��Sǎ���hnr�*|<-MG��pA�T!gX�qk��T���f��������=��yE���� �48�z�)I���'?)̓��P�%tqS�Hwx�0m�"7/歈oD�z�ʯ�b���曗��Y �K	�P��7�@�㱸v�Y4NMM�X`���4` ?�@�� C�80����-�<�s|��|� 7���t�VV�e�m���Oz%�'���C��ڜ)`Ǌ{d�X���h��_�,�穪�%N��#x|��Q*�F"ͪ$c1��|����{�Kƈ=Pd��	ʂ��r�3<��85&�l�-��
�:&zw(I	E)���BG�#ͻ_��sz҇ ߏ<������-����L��E���u�cZ�N�#����+��.(�N�����8�����-��K��~M�1QJ����܃(�{?��[%
�?���Vɶ���1V1�[-GO���r��_���+/^���O?����w� ���b�\��4�?V�����C�G�?�W���Sm�.�Չ)�I8^�u�d �v�|{q�(�%�7�h��Ee�Z����Wi��f�Y�b@>n�;9.,z&ZX��Ț�e�>< ������9D��f�f��*���@�����縒�"�L ��Q_���H�p��MLOSy�Ji2��5x����Hc(O��X������^W���d�%B��Ź�? �����$(�·�'e������-��]~��ʤf��~8�-{a`a�҂����X�T�P��L)�K9��T�`0��d�_sř���Y<��DB2U����T����cT�x1n�:u��?L��җ.�%�r9.�q0*&���KI���gY�Չ�S�!2�������Nu$�h��HUD0�k�'���ω��QL�
����TOܺUӻ4l�qF	�}�r�)�*�HTPw5.C����"����3BZt�-_�����cg�Q��&�C.�TnR4����ő��"�fѠte�Ʈ4���g��q��pk�&5�����E݁CfN�؉Ks�"Fcq�2ö���$��t:7�?��y�u.�R��?�:��qƬR.��bz�O�3����M���0���������ex�p����Dݍ�����Ũ�L�!�!��D����������pec�ڃ>�iC���^���������C♁���&NE�кp_z�	��`�=�M��!��^��F]���H_��K7����|��g��تc��?��#B�j����{�9����쬀��qt��6���x�@�}H0�|�Έ�, {-���ⳁ ���+/�D�\Z ��~��?r�Ξ=M?��d��N<�xᅯS�� ܳKc4���O��^oY�Зp�\uǃ@$��L�h������&_�*���Y*�J|,E��)�w�!_JbqX�q���Fo��w��ez�㟤?��?0����׮�5��k��y����ɓ�i��y?p��7���q&���<ǯ�C?T:'}dݾ�	� LL����"+PɁ06.m�m^�j|�C�;��y�.n���Ӕ���t�J��y�_���?�W.?����B�&H�%�o�|��Bbirr�._�@y6�q���%!�w@�UQ
UD_@�WX�yr�X�`\��jT��J�VЬ�OG������e� +%����}<�QQD%�((վ"�O<s��u�1��ki�	5���B�OD-�?���<�����=^����R1RI8�DҺ K�}�s�%�h�c϶��'�{�}$��ۿ�]4�}�~?�ה�T@F���^�����y��Q��
��V�>?���յ�{�]4:pG=�71g��G���թ_�[����t�`�;� ��̦��{ߛ֧*�v��[���S���~���3�O�fG^x;�O(�Ľ��&/��?�C��Eo��7hzjf[v�̙��Px��5��<t�L֓�3��ŋ�0�W쉉	^����j�����k4=3M�K5Bt�C�LMM)gd�!K��Ak�k���,���"/�0��wC�A�	:���h6�R�� c�	��B3�@�z��5�pT�Y�rI�{nϖ?K���h�ccZ�8x�1h�ɵ��Ҽ(ApС�n�!��Ē�����4l~6o����,�	�NM���a@5�N��P�W�_ћ7R"7�h�S�G���4��<���z.|]+�1U��z�2A��q@���l�����쉓497MF)EϽ�%��X��ŋ4��`��	 �l���`��f*�^U�&��Wm��ꉸ�vf(�Z�}���TO|p�+�Ќ���� � V��{�Q�����q#%w��͞f<��1Ep� 4[	2��t�e�>��l�2߷�f��N��� �h��V���+Fs���ͧ-_p[��j��6��5�`���N�4���TH��S<�4��1���8c
�Z��cъh.[�"�s��i���;�������f���q}C��N���9_����8���9$�%��q�8iM�.�r�:��IS�RX�*�B%D��\��&�@�??Ϸ%s�������ct������I�%����/|�P�:a�)0PC����*E�z�&|�VW�O�XŉG�(J�d��D��q��Й�RI�s�я��?�m�o�o��o�4.��|�L?���g����{T�T�`0��5����d�H�Z������z����J��$��1�dm�G.ѿ��_�c'�´G� ~ɼ�h��������'0<�E ������.��qj
��@� Lt��� t�mQ�蘩N��T�($���5�Ag ���%IH���{T��s��9��?��{$�>�g*M꠯!9��=	 n�|Q�U�l���-�r�
|=�83m�X%I!� ��w���:�6�s�D�G:���V�Ai�լ]���4��i��s�:A�LF2�p��jvi�ѧ��$��0��kQ����k��XV�����jl��� Th@5��	&ҽ����j�{p�qq�Z@�jKz�dl�Y¸Wϔ)J_2E�?Ƃ�[T�H�CE�44�(�`d�L���(�_.d����@�_�C%	EB�K��\�S�d�G�V�Փ! 9�*�6})i��{(D9#���ک�<�'|/hx�v�k���ޛۖ��a�����g�<��V�.��%0� #.%6(���H9.���C��@R�S�2��	q*�r��!		��oߞ�<�y��Ƽ��}�so�l,� ��S��s�^{����y��y�74o>���M~��&�	����n��g�u�SE�[��ðM@�/;B��I������_�q���++����+]~��������\�# �g�>��z�֭�3xjPL�V�����pp���[��D�4[��A4���kui�g-Ly��+\t�|��y��5.��߾ݒ������^{MZ���`/4���_�A<� d��Z��Y�o6�P�LvS7�.�_``�إg��͛����H��B�f�����9y�������/�p�>���qpL�麄#���V�g	�fhM�.M��C=�B���_=��u��;lU��޶�$1��Ql3 	�"4�u���P-a=s������I���NR��$s+s��3�n\*-9]�]��[Ed��F�50, X�Sv� N[7\!cY��+}�N��\��A�'���}\AԌ�./�#�]�-���J8�+��d�\d�ܼYH�6��2�I��,��Wh��B��%�cmL���;���0�����tl_���q�T���E�5jW�%r�A�l3D��!񥦆�`2
-�o����pR#�9N&�e��������*5/�J�.��'����p�Ƣ@�U�r"�ZA��wd{o�R�P��C�&LF=��q���&���3�)Ε؆��R�k^�k7WP�H	�e���^�*�~��g<���-T��] @Y�3�������#+�j�2 �Y�y�X���U�����,豙g<%��e`�x�%���z!3*�F�^L�H�j'�0�-.ʌS�?�~A
��l�{܁ ���Gp�@���n�0��"Apˬz�A����.$� Jc�Ws�o�j�2" �	�}~q��g2����Os��o�P5t�C������T��?��
Z�)�oܹ#�34�a��+�ɻ�;lu���jM�?��ׯ�葧諑��`(�u	
�J�7:r������R���
��ޠ�Ap��̅W^~YΜ>'&�w��hh�!g:ό��</��m�Z��чѨ;I q�ƳDұx�|�y  a~vVΞ>#���?�_u�m��?N/<��VWe0�˯�L5��c#(���� ���^/�z� �/꽟x �U���>��p��5q0�h���2�l�AB�&Nx�\��gM����+���*�+�9�t\�f�MJ�'�s��tzK����La���h=������)���Y�	�:n;���1d�ab�����PX����<G��U%"*L�~V��Q0��u��Sڷ07pM��F�}�g1�-?=�{���>Å�pv<�ա���dH���U?�7	��bV)�a�s��#Q������d[D�ώ��s�������ߥ̕����Po<|��2�����x'��.�||����C��͎�M��}�����|�m<'��~�����v:ݯ|�+�V������o���>�Ї>$G۟�v@��?�4��~Cg�K/~텪�8I�Pp���s��ܴ�V#׉C��J2�tR�e�*�g��:ic:�rLΟ��ū�z���~���5�q��|��>&E]D��5����:�"H,��ۻ*��ַʌd={�x_�E�Pm��ܑ{��)?�:�(����R���+��&]���M�]���V��7:0J
rha�E6��
BNH�
�=��G{U��H�陣m�?ca��  C�~�Y�[��Qpѿc**�j1k��!���!:��n?��\�N��B1C*fHp�b�&�lUC?}3`�%V�Q��n��a�\�yd��S����B��adH�Zτ���}脬n���v[���� e��K#JcܓU����b�t�i���Zֹ�L`J�a[���*'�I�Lm_��wY���Ӟ��b����1M#xq?�&�b�,Y�w�$�Z�:#�n�o�q�,1ޒө���3�Cܛ`�kmH�.�ܚaޗ�t����e���_)	�Q�S�*��{7�j�\��c� �6�Y�-!�r��b�Mo"Ɯd��O�J�ˌ_�U���9y���ra�4w{ҟD���K��܂�-.��3'eva�^�4� a.�1���QHYT"��cýˮ�������D�V�3$���0$x����`6GŤ�zD�Y��+���F���5� /;�c��8ń6�c�P��	���^��!�M�F$(�T�*hp�ȅ��o�Ϳ#��X?�a?�KH����Ǐx;~Lv[;$���1�P�Db!��}xBy� ��r�$瘱	��N�!�L+2� ��j �W�8U�����ro}M�}�{	Ԑ��Fb	$TF�ˬ,4�-�}��%����
z���9	��$��'|8���X����0��e�
�Q�<��'�Q��u_���D���?&gu���a��9����O������9����i&��*�	� �f������8H�'t} Dj�we�XR��|T����p�`�󄂾�nS*�V�9=�,O�yXNT�d�2+�s�R��euܞ���A�%���ESR~�lD6�w�翤�x���h��[s[nܸ&���1�Q�j��+̱ ղ��IX�K��I*�8|�%��p�
��V��"/�5.4�[�q}3�r!��S �1�����L�Ɗy�S��� oY�A���m�s��&�����8� q?h��f���p�O,G���}����)"��T���+��p[E��_b*&Y{"��u�JwgI*�>�xr�~�C�յ̱@��`Ϝ�2`���(�q�G�E%��,R��A���#L��x��W_}�c��7�`�v��/��?�����?�����0	��D�RmJ�d,�{�����f��~�:[�q�}�x�h@d�@�D��&#.��[F{]_��O�����t��>���޽�r��K� dL��dvnV��7�ބ�����������CB�TfY�Z`~h���86=����6wY�.j���
��U,�0������$W$���������"O'����I?y=N�9��q���p���2�4�|�1�[���O��Q�n��)��hv}�z�@�7�G_�Q:q}�X�]7ap����~tr�ࣛx��#�P � �2������ \}�r�!���*__��f[�H6�6I��t$'���L Ͱ����� ��-T�	M�!F"Y9'6�I���'�����dY��,���X�,��U���#�d����'��/�a4fZI
����kL*��m��~� m2\�$�BIb�a��2�9�� ��@��:_����=�n,�^בށ^<d��3����c�0"��B�T���R���lw�����|Mjqf���2qM�|i�\�P��ͦ\������tfn^��������	cu�a4���t����,�8z�#XG��)���!0����z�u9�:d�2�Q-e`P���f������'�Z��>vX�`Eo8�v������7eayN��D��~��Q�P`��)�NK豯@4�ϱj1"}Nc�t��2lz��T���͇c��5 ����N��J��	S�� �i�r�4�+� s:�$����U�1dl�ܷ�Qb��[��>(?�#S��|�����\��[�O2Y�9�X�V#1�f�Т72����e)lސ���R�$�]|\��9�1ȝ�E
�FwG��{RG��EEwO�Q��yb�4}�B��F���mX���g��<)�z���'�WU.^�(�N�%����sW��_��_�׮�*�����ʊ,-�<�9|���)�U@����`x({�]�{�w�9*Kgؕ1��<�̻�N^���R��?�%FR�)0���Q*�y�%y��#rn�t���*�gfNg��DNW��X?\�^�}y|�I�l=�* ��N��+]g���ҷvWrSz�Ȗ�&�X�]Z�IZEF��p@�b�4E�P�S%���p,w-F�"K���A.�}$S�6�h]�/ �ⰶ������`����s���ٯ|��n������p0~�"�8+�߇�+2�(��p�%I���Y�҃���Չ7�c�	g��V�r�����l����j��+"ߌ�r؏#�v�NV��%�Z�8mY����K����ӏ����#�P�9ō��O�'�yI�n���/��?�h���oq�<��$����>�s�`�;�d{K�^Z��� ���1�[;{l��4 k���ⰶ���϶N�E��sǠ,%_�|ِ�y������#�}��	H��+��t/��7Ҡ�/3h}��E�hp�ԓo�n���d,J��f�=�l�C�v;--]�Y�v\�����:(YommS������g����X
N�6�X�	�O��p
a1��ՒJy_���QuJ����dQ��J/L�Mտ�Q8N�F�l�x܏�Q.dr=W�6]m2�]��#���v1�\���RʊCHi��A���xe^F�P�Uge^�&2�a�AO�Ar�V`6��t4����qB�dG��O)�S�h<�������>��p>	�[C�4�/��)�`ˤT�xdٷ��|8�g%�s���ߦs�.�8W�t8p6�.�i ��� 't&��6e���kM�شx%�4�H�L4�Ć������(ҏ�:/3�r��&���Ay
~�1�p�ST���TZ����$h%3�s2�����!��@  W��HO`���-�s�|�e���ʬ�:��� <�h�B�dD���[�;�J��+S�����e�.�
�u9Ԑ{���B^f=��fT�(�ko��0�5p08q�ܪ��+� ���-���<�yKKK���dcwUoO���* ��b�J<b��9l���f�S*��}W��� b� h0��:�4Я���`���N��sK&TQ�q3U�J	*YK+RW���ډ�z��@��8�ǆ���b��@fE;[A��u���1����'�׸F�����"�3%�ӧN��{W��/>t^���U�B�^��FpBh	�|Q
��[���ݒGO��HA&�b�V��:�;W�g�<�fs@�1���tl����*e��~������"�q�{@1��˖��Z��^V
$�u��^�-�N���Ο��gu�������2�E f�: ۬�aH� |d:�Z����H���Z��۴j�8w��i�̤�!���ǜmH�PU�KXmX�]�M�ק��P0�'S:G4�my��o��}��4�Th+U]��9���:FL�s5&B����0sZs��b�势0I `�K(hU0����+H�\!8�i�=�\��vơ�����y2�S:[��s $�}ۃmD�J��JSg½p�e�s�
c}#�nYr���`�����Z���� �7G��2�o���ω���#{�am,�'����y����</[��{�=z�q�0�~�|�k�ﭮ�x�W�yw���B�����������s; ��qK�=t�h@��b ��Cu�Ĳ����Q�AUjԓ�^�"�++���A�F��qc�t��T��_�tA��� ����[�l;y��A5���y��P�XY9F�`Q�@[2�h7@Z�d�F���=s�m�B��V��*0���Fuz�u�on5��8?+E�+�!G�$��&c��r2��	����%ϷJ��I��(�a�Ć�!���Z�x�����tvf���@Έg�!���:���6�z��Մ���5�fc/�B�ӜZI�ϳ�˫K59Ƴ�^Sp)w�F��J�Ǿ㌤�ʽQ[N��K]A�N�G�3�1*�������Y!*:��`���YN�66;/����������M��	�u��CǨ�g�k�l��k�������4k�Ԑ{�n	�A�m�b�#Sc1�����<����* Ls�T�m�`��dc�����2�q_>�F�����O�]g�d��v�)}�Sr/쐜]Ѐ���a[���K�r�,e��Y3��O�$��C�4O3>��XY(���jpR�@�NI�)����ʔ�i 4b �1�
T���"\�V�!
�����!	�)�Шp����3IA�S�89��"����k���x���l)@�J^��P��!�[,U� ,� �8��߇�$�񓧍|� 	�`;t 6:���z* `"�D�:�$���[(�g�h�7�y�^�їJ9i�nj��X�\3�@�p$+��23S�8��r��Y�Go��1'��+�`<L�dg.��YZ:!oy�%in5YA��x<�����c$��'O�8&��j#�2���&}y�%�2�o���肧�ܸ���vSn\�)��]����Y�ق�{��^�;Ͷ�.����/����ً:����M�x����YY�wWv�6e��Ke�	3Ð�pd��WE�$�*jF�l�p��u����ު�W��}
В��MZ���f��{��Fc�����ถ�����<w�rU1���?`�Z�/�%y��#z����{�����q^+Ͱ}��Y��	��Gc�᠀ӈ�.�g���ա��i�={��4�{�� ���[�z��$
��
��ft��Wdnn�p>3%s-���w�X��3V0��^C\�@��X�T�����A><���PL��-���cB`�F�+�:XT PX��5�~�C?.�~�{Y}㼏k�[��! � �x�1<[7Lw�����r�_��=�_k�`{ ��Z�^����:�m��~�XS��g�N��yk���o�﷈=p=��*ɛ��NKr������aפ�=�g�T�֘,a�`��IL�����n0l�����_�^��hcg��/��/�r���ݎ ȷ�i�R]��x�����$p{�D��<�M"'|��[�J�n�G>�;������Ï2{?%T:}^�js��	J=;�$����۝��*����瑼�B]����n1�E,�H ��m�p"6�K�����k����-�³�����֍�.Zc�A#�x�c�2~��I�(_#�Ģ�S��	f,�vc!��P��3���E����U�����0�A�$Llh� Q0�A�߫�Ɏhۂ��Ɋ%~&~W�U��a�EH�edx'$ ��DԱ�y�T#���0
���%��^����P�RNc��M�K�6���j��7�.�X$�@��U��^�l�O����@7:ׇ~d8�����M�:FU"1��<�vU���IԀRk�E=q"ə��S�	7�Q\,�{�}}��}:3if���/$&������7�G�:
 C�"ǐ@)3:���$���b��� A&�B,z��l���B5��qY����{䙓��q��`�Ly9�����_��G
��A�lqL�l�:��"eU%�rl��Ж����"a��Hr�~��P� AH�~dR񵫁%�h��],�p��&��=�J/����ز>���$dfC�L�	��ȣ�8�mnl��J�Ė.�߁�C8N�>:��"E�b��� ����>r��3��xޚ��� �ɨ��l#Z�8Nq6�Us�}����#V�)��AE�T��vK6�{RL���k�uS�_�������gt�ҫ��.O�71�oH��@(屠"0�� ���s<P��֣Dc�є�VG��{��w�Ζ���sM��#���l1Eu<*��ڃ�mucU���cl��ْ�3g����Jp'T�Od�ۢSx�yR#�d8�����NS&:��wd��=�V���C�K:Ne��375'7׮�^kO�x��Գ�HO��<�I$"�Y��>�?ཀj�F$���Q����ǿ�r�Ε��.���Q5�`C}~VZ㑄��I��l�J��4TЉ ��;��n���~qnQ��}��q��ڐ�����S�E���l�C"�ɡa�Ǆ�� r�>T�b��3؎��P����8O��D�=p^�S
6��\^������LMN_ֹw"w�>��p��2 ��Hӣ�sP)�ܽ!��>>Ӊ;����S���M ��;�*�9 �e�g��eV���RW�i[�qt!� ֠��86�~_� �48������OIr�| B�}�N<]��ص�p���{Lb]��kq����WA�Γ��$o8W~�>��͉��~�XS�+JL�O,�$[g�*��@0#�|*��ْ�i�.����Y�#���8�����w�^jv{��N&�������_���|���;�k0�u���8�U��0
��`�W4 ����h4�\%*��������?P�W^}]�j��#��N�/��(	#��u!�z�*���R1q]��{8r!�����P��Ì�-Іp��e���Fp��J�V!�	�\T	���CG+���r25Uu��=.�a8L67�.+,F�?�y�p�֫j�����n�8FB74��Ad��q�J�Z��7ڦ�1��hT{$%h$�E,A�"ЎdZR@+N��$�N�EQ������@�"����v��өt�I����b��9y�D�/���&�'&a�ΜS��k��=��_�M�f�c.�D����Y�u`� ���a:�)�*BB�'Tb0F6������cZ��;�g�f��L"��_0��`dXY0PpER?�|r�NF2�&�r16���U���d�]���ވ9TS�@֐>���`y=������YI��.��x$VR� %�~�"���.��;��� B�Q�a[�_���y}�~\c�x�ܣr̛�Z�R�kԸ�<>wZ&�H�&{l�J��.�5�H�bd.����{;>� �M�;��t�ӐyF+^U�tE�|���lԧ���[[ �dsg[�u` �ԩj �R��<À=� ީާ]��`Ɔ�+��j��C(��W�ִ,�@E�7m$�T�J3uq+%�r��l�4������k�R��2J�G0�Ӡ�"��h�y׻�!_���w��`*�{����UF��[S��e+$9P
S��d�Ֆ��k2S��O|�cR�J����ԩ�R�@4�UR9�#	���W�����o�����W6����@�U	�Q9F �X����gH�/V]�=�,��~]�]y�����;��q�T���쉓����=Ӓ�c�]�{�<��~�/KK�z\5�U�N볈:$^p��Vjޫ���-T(b�gO�wkoC�x�r����H^�uMf�5�p�����p{-	K�<���Jc<���.�t�m� �=M�U0����#��Q[V���S�u��j3���o�2-�y�!�w���]i��WaЙJC��`y��ERϧ��}wd������	�9`��n�ݕ�t̼���UIH&U���5�dv�#&/0�01cčI���u��T�A�S��+ ��ʙ��FsK6��ů(�Q�^������<t^�Ŝ�\S%�>qZ��)V��1~�ӧ�o�
&�L����?������ȶ/�˃�I���lG��6Z{�z}�Zñ��z�}=�]�{�	ϟ��^�'�x��\Y MYe����W\�nr�{�l��d�C�|�������I���������Ϥr�!��}Ef-5Us01v�c�r�A�?��9�~e���v#��1S
�k�����S�����U8�x�a��n���}b�¸z�c�tV�t���8
��N_���|�_�pc���GݣV��\� �ֶ�+�^noH��s��Q�N�|N���AL_y���#�ɇ�i�i�s$�:�-�8�.-s�g�Av�h5]h\���,�Z,,.���<$�=�=��K�����u1I��K�U�E�Ѻ�A�j�$�aR���}lHd��J.2u�(@~�ק]L,l��]�m4�A>��P4h�2����)�)huqJ4���>�0�����$!�������\V�u�J5x�$���I\����A�	�ph8�&c���\�t,P��-<w�$j�����J�z}7t_��6�~�ޜ���������O,i����־��\-^J!O��da�?��4= ps�p�B��Qr�=J".h�@�n9�^��&�<�^o'5��1mN��dט"hF{F<a��f�$7�7���qJ���Ù)K����(�$��ۥ�����L���1dmCR9�yKLK�%��+&�J��/a �����qG5e<��<�/�W���#��2���>i��8�����yT#�\g40Y((P��Լ�8QJ�0$l�͏�69�@�-����0"`B��̸W�=#�wz���D�`G���r����֞�@�ܺ�V��h������>h#[^�gfmw�~W�qWJgV�m�h��R�j���B�OiQ��9�B�*v)}R�����E)^yA�����ې����jC^��E9����[�eY�Cڍy̡^�K��q�|ӕ��_����� ���՚ -J;��������xj"�=�6��k_��>�Wnߐ������Kr|�<�h�
�����c���C5؜�ƽ���;�)�Z�كы�S��L��:$ڧz3~��?!߱xA�]ҿ{��i˭�U9��'���ȩ�oɍ�oHK�An���W��±�� q��v��6�3�rRA �۟~F���e���N�����z��~��GJ��#���c"%�`x��=��\<���?yV����3bw���n0Xn)���1�4��1Q��1&E�{���M��o�\��Ϟ�B��l0��?]��_}M��ʫ�N���=����涎��T�Q��}�k�?�q9� L�;F�W�^��/W�]�P�ʹ����d�sȩ<[�L��K�E�FFF�-� T�|�lQ��"KK�mZzf
8BA$��'���f�3?�`U�8/�˅9�6U6I}��Պ_��0�_��ְ�kժ1�M�I>�z~Il1�c=��i�1#��h�SPه�
�[ �É���<r�qV�p��?�I�Ė7�f$n~�}z'5�Q�} ��=��/��k�L(��'q0Ae��o��c�;p;g�31���o��Xi��Z��T3��#��&�s�����n%�Blᆼ��6c�� 
�sC3�$5��AP�Ӟk��%�Ǎ��I����3S�PJ�qHOG=1W���:h����c͜�a�*zA�H�|��������V�|��ŋ;����X����� ������{�����?��L%�L����tE}�ם�]��z�`q����U���r�^tmm^��⊫����u�R��^�}K'�(�T��1��g˃	![�����^.�OBڋŢoL�|�, =�/��Q�׋��_�|�ʕp<G�$W�*a���ݺuk��T['�-?�����zy��~Jg���b�l��|�͢���,ǡ���
w�7�u��������lK8���݊}����'8�C�8���(�6}��z���˩QNJ3U)Ǿ@L���绝�=��#C~dЂWgb�Y�=q,��dn=��8o,��_�Q�J�˘��R�ʶFA1�.�h��g:������m����wP�wۢ�
J�|e�~d�rF���X�l!��<F��.�X(}ߌ"�!�'�{D�քEF�zMPuÍ(§"v������T>��� -��Ҡ̱-g���DL88
f!���F�Qa�y��;��ގ�jz>�D�5ț�Dpp��k�q����-i��r��-9v�4� �P��LU�*��ù����s��AC������(.7�ԡ%�6Ӟ�%��D��,�($�ˣgyI榗�\�ՠM�leJ��9�� g0����.+s������SR������Cy���)噜|�����*6S ����F>�N@d��|�E=�_��sr��9��+_c;��d(�p(���P?$�����h���	����E�;6τ�iT���X��D��Ո-��VMĈа0u)�������L�*]��-��o|���7nL<�C�-�Dݺ}[��gY)����ʩe)����{���QO��I�A�!�\����z]��'��=g+���c��7�tI�+H2M�����<��9��0�|��T����eo�w���ܙ���䃠�����g�� �c��х�g*wՊ��!SqC�ltخ933+[�� �P'>��;=�*x6���r{��k�ぴ7��9L��
wҡ�G]�y��k�h�����tz9u�/ǎ��k�ݾ��
��݄9-5��u�X

"*SE$x�5P��t�5I'�Ț>mG�n0�_�~E~����W��g�X~hZ�Lu�1�7A��A�|8R��)��/�I
�Z7
�)�	s+�x)v�2��!�T�� ��;8y�^b�E��
��S
�g�9L�>\�x#��`;RR;w�r�'F>laz���&|ۏ�* a췔��B��Pn9�+Y�Rx��*�ڙ��ۨ~�`�%�G�	+��³����d �bV�\v*8FՅ��8]r7� ��t�����X�<��_������&c덒:_����ן�ݽ�hk{��"�_~��K�t�t������8�h�K��?����|���K�.�Z�M�����_�J���bY����x2��|��M&g*~�~��I���%�~7vݜ��
A'n�V��a��1z_\�'�I�~�R3�����,��⮂�|��`"�\�ո�8҇���D��.���N�������V����駢�2��ʓ`0���z<55���Y;��d�<;�K�������o�O�>�7l(_�2�$��6K٩�_L2E����}:��B�X�iNfq�V.�f
�R:�ƙ`����
������̛!1F�L��%�Y�qTj،��
�{�}�A�Z �w�Pi�LK����84R�6�'�B��p�0�E�R������f��{6�6���/S�}�,$�M��PJxHF~��А�@-ӕ�~L��
4�fX���gB9��_G �W�,>��4G�p+���?Pr4@t��춤���07;�c�3Ў�����u�CVS*su��k��|��W����z聜<���"&�{�Lޓ�ֶ\knʸ����##� �2�k�c��
�}n�>e���rgT�t:������yfE�)�8���|���'~��r�����|�uY.HU��3Ͼ]�î�[�I�68DP�Be R�
�4xW [M�N`�qp���69S_*�:Β��X����/������������_�����<t�Lk�r�F]��M�fi��k�N�)���4������Q�"sz����Sp�z�����4�ղ� ��ֶ��ݔ�����o{���F"v��)�����o}�t���<�����C�9fK����ݑ~jd�R+���	&�7��SH�J�n����O����0�}�#�Աzb�Q��g�
eh7�uɡ �$r�l��bL�%V��
��C��>�u�U�{� ����Q�2��m���ֱq�� �B�KrC�VMXa���c
�� ����X*ȕ�U�����H�ʬ3�@{(��|T��tc�Z6M�}{a<�<��Ϗ�"�
2�0p�aK��͍5��{v#H�����:�����?�)}�t���ރ�x�j�o��:�9I�5A�2�礫�!D���'�vG�Q���V��$���ah���=�xW��F����o�g%ǐſ��ӿ�fd�r����w�LY0�@��^�8�ۃ�-�8x���V�UՂz\�9����L��g��F��!�S|l��||�����:
�|�%8��b]?p�Ƚ�l�Ox�Q݁@	�r�2c#@�G��h2����#� �D��M?(a|�[���t�m^_���xw}�+Q���@9ھ��# �a��׾��@�_�Я����}�����9�=��I}�E��;�N<�*�%�
�{
TڥRr:��o���;]+�R�~]��F��ΝK>�����;�.�[oqqѽ{�.�W��~�k��of�Z�
m/u 0�(X�04���\.A6�����2�m�9��TS�N�o�8f�c�	���-Q��D�+���R��ueYZ��5ZA觶�	���!��si������f��>(����}�d��b�k�
�Qd�@��''b�5�7.�`���q(�$�L�e���p�M��ⰷ攸P���N�Yv��4��� �n�-m�R sL�(�3��; n�L����L�b�ѐD�T��^�4h`*�g���RZ����JsҕD����$�ס�FШ�(�4�� �2TvZ
44�[8�$;W�"{�ݞ���2�w	��]�Spp�C��V���T��	�
���R��:C�iR���۞o�HG啥9����q�����c&�*�����rY5`��O��������/c�].�M �gm�C��У[�#��t�G��۞y�|��>-_�z������9y��%����!]E�ϼ�I��h@���=��^�O~���M���/x?P ��i�)�t"J|C
�X�3Eu���p$��>�V������˯HmY��%���G�>-�{X�j��L�|��f*z����ob��e˿*"k���^�u��s�Js�}�����w�["آ��ژ5����p�E���sŀ�hG��YH��d3V�c����.�dAfb��m0�c��|�>8a�اlz��	����pD�$|'P��Dp�����U��^�r~F��lȨ���E���,-�eo�/�7��P?k��'�~@EE - ����ѧe~~�.�s�L4��������I�$�~$����Kz���t�,K��͵���J���;�����JBU�1+$P0���[����Xǘe��4���*ƳE.�)>�J�c���@f��"��O����� x�:��r��f\�7'fg���<��^�ċ��S[�Fu�H�F��)۟Rq)H㒿�p|��� ��)N�9[!wƳ��N�S���(�!_O��K
A��(D*���n���T?4#׷�` �
9�G��E2C��$�(Ve�D`���\}���a���ݸ���]���������Qܿ;���'~b�8�_����v@���R[9��Q��f�Ɵb�
��O�+�x3Q���_�msu�A�N�@8��a�(Wڱ-J�uӳmVh�Is�ȋ8Ld`�0�M�Ad���&C��ӭ<wp�k� z3P7��! �|hT?|�[�x�p�U��;A	*>47�Ƹ0Ɇ������y�s��%���qp�F��5�Sr��#GE� x��� ����XitЎ�1���F���a*	M�x�\4Mʉ�vJr�2/s�<�pR���d4
�� �*S��;��$f�4���������D�\��6{z}�
hn�6en�����A[��bN��'t�����M����9�&�T�2r2��du�-��X�E�����_"��T;�J1+I�0��y֦��3`�+�e��j�`���A���{eٸvKv�ݓ��MV�f�f�X+�S�-ʉ��j >%;�  51���b�^#���(�z��@ːC�m��z]����c$7]ԟ'��?/�.=#���4U��d(>Ԭf���[)���S�C0� ��2�h���#P��@�����JQ�Y���,�+d�"�|��#s������̂���66d��=ɧ���G�̥'�՗_��^S.���p��v�8�c��p�
,�@��-#[�CD'z;��+(|&�Уs�$�І����X�00%�\�Jj7���F	�qW�;@�W��f���Sk�i>p���.�XM����6r�H���҇��A������e[���������S�}�եt^^�/�
�~�O����J�5��tD#ͮ�����pϺ
�!�|ocK�;.}�@V�Y}�\�E��_��e��^�<��C�%'����^�H�(� ��3��X���i��)GgH��}�sl�=��jT���t�m�1UX���B���	��8E���=*��8�����^v�%N�L6w�|e-������h�|3:�U
��9B���scK�6�'�fp��hn�f��Nk�y�(���M�K8��b)Ю�x"
\T�<��]��M�E1 U��r��~�J�y8&�B>Q���W�\�4�-��l6�v��4�?��ruzwnyy{���[sss����Ϧ��O��O��������z��m���(���ث
c���N��r�����7��<�TFH��� b+��j2�� ��`��M��
"Y/1v[p��V"���z�O�CH�%;���C}������ipP� �rm�=�`�@����`�)���.57�f�D��[z���΍Y��N�����@��7�'���c��7��#�s����ȱ3r��`&�y��=9P�2W;��Z:'��y��|����Xl�r
�4&����o��	�{�t�6%� g<�"���#`��2
M+T�蜍�kp�Q�����N��#�i@;f���W� 31�fTJ��Xd�H�d=c�-����xk����Ⱂʽ@��P5�;{b^�z^+�S�4� �fcv�?��z{W���e���buN�2���"b~��nP�������`>�lf��T)�~��W/S�Y���9��i��Z�k�-�LW%~Q�.����Uy��*�G����k~�׽vK�0'-��br� �	"��5-Vi ����/�|��JI��꟯|<8�/}�s�x߉�-��]��aɕ�;���`��<!�3�\:��\�:�^Z�!��6�+T�}Zo@�ls�z�B㛢�>�U��{H�S�ښ/!����X_M[����&Oc�	=.�<�� Bc�=*�Vx���Xxt��9ǳ*�5�x [�tÁ̟:.�I����B�=�9����u�$e��d����{m[>������(��m��ؕx�����6��3�Juj�\�3�|�������
��ir�7�����yӘ��ps|W�
,_}�e�Z�G�
m.Ln�P�|kEA` �賂8�pt�1��xjLh������k	#�QY�*L���{���؍Ӏ�,Q��M�}��]�Xپ3��k~"����a�H��'{���
P�wa�� 0�g����1�Mm�mj]�c[]AU
�I3>�YU�(���b���|4��J��L�;� ͐'��pp��jaUHQ`��H���b�\���q���;����^�Tze�^���+�8��ں������������^���:� 9ھ��;kw���}����Q�>�M����r��g��N�n3NlX3�p'�4ԂLm��X҆2YXE�\I"u�h�,�|`
���	���8p!��6.l���Ll�4�Yp�!#��#�٩D̹�Dl�W����n�v8��! :�b`y+FQ�TFR�f�R��ˀ�c2fdt��mu'�C�]j�
]�8s���/z�iv;�S����-JHv�"�m9�$+�k�B��ҊO�Y� Y��Գr�����O��,1>�.��XB�z׾&%�K�x+��i)��ҭ�W�Pt8D�I��������,*e��h'2�T��$C7V���2��Ep�T]�gvD�����wlYҿ-,/���'�:f4(kpy\=Vp�n�;7�V���z�&���;TMJČM�60h�ȕ�z��~u�j�QO�%���H�gC���暼eeAj����):շ�X���lmK4��DR��WKKr��)f�gf�)u��_3U<�6��r�7�2��QIr��%�T�ۗAw�K�@�P�I��
�rb�UGkc�o�"W��g<������1zxF�QӀ�-*�pC�i��+/�LyJ�SF� ����F��ׄ�H��D�O<�X�c0���g耠�F�b�#尭Q'�?��Sc8�G� /�4���!�Js9����Q*����Z�T�����Acc��k&%���
�����U��(`����C^��?�O�*�5<bsB��)�ľL��H{ܧR�zkGF
� �ʇ��3�^k$=,MiHT���c��U�c}�n+0L<��Ge&�1'o��LJ��}3z���E�!�X���9�R��R�λ����a2�#ak��DPAґio�-N<�íO�C��?#���4�'[�E;}��b�h��F0�0H��� �5ȴJ��,I	Z�f�xV��Ȏ	~^������V�^��} �@���1J\:^��x�֩����K�A>_hU���0��r~�r��ܜ�:hwt^����!(��T�f�'N��ި[,�^�*�����o��ԮV��#�q�ގ ���m��ت�8��F���)x	��:�^|�)1=6,��G�I	�ni�Ȁ�\+ѸD���r�="u���� >ӥ����5`��p�5-Bό8K�#˅}9&�e|4�C�c	A����nn� [�sqKD�@c{��R
��m�|$�W���]CD�C��J���d�k�x �P�`��	�i����y�gOG�`���M&t6��#��1��-a����g �����/��"�N�5 �uKҒ��W���J��-�G2�k[�@���ܽr�,���A_
��߀�`�f{L%d�V���*2�Bu��z��T4ǂ�#�=�1{䁦hض	V�Ԥ~�>) zʱ�9���}=�PO*Ueg8�{��K����L,��0��!h��{����^�W�CN���l�V�׈�=H�59���π�u�)P:�ar����҈����ե's�G:̗�?�l_X��y�2%<��������w�Ķ�27\����sK����0�,3�����g���va~�$��kw���;r��蘯��e��n�s���o�u�T)�So{�l��%��G�3�������OH��R��*R�Ya4���rޕ�cK2����},c�}����vZ����1�@�?�9�#L�yhc o�V�A���a�]���d�)�\�"2�Hu���d��ooޔ��Q�?K�3		'�#�^�B��\(��M�n�!��z/C�w��`KjQA*�޿Ib@��}s����;��c��^��u�(d�l��?g� ��<�]o�O|�S
N��*2��긅����9&��$p _��h?�Br�k*� 
�|� ��<4�S��GA�����R��ƣ�B�����B��l1�\Qm%C�X
��<,2?ʍ��}F�ߤ*B
�$ ��/b_�x�k5�$��m7c�Ź��D����:�׵$j6�����qC���~��`8���um�(r�|<z zۂ�d2�ׇ�Zm:�yp���N{4r�ѹs3���g��W�?�}:r�m��v@��o�-���歛r�ы0;r#�5 �u�.I�D�� %����=�	[�})!�S@��T5`(/>��uQl�Klﭐ^�*���~���f�@'��ĩ���o�J)Ayx3&�v���kȗ�gZcE[��{RKr'H ����8�[���!v��.[�4x�y^ƃ����Qv2���d��%�m?�CP'���5r��QG^߸)��<&�¼�.��꒸�-��9d"s=XLے!����Lj��S�\>%���dt��ǎ��&�*4r#��`f�C��Oa_�7��f��� DLu�$\J�r��~/���`/Ҁ��],i����=PK�2R��n�Z"K"��Cs�嚎['�:�Mٻ�.S=.E�g�� s��,(�hIb�=�*ڵ��"+m��Tm\dbsU�]ǹ��F{�NKqАBOG>�����S'��פ��_�^���nS��O�]�
�E�O�|!��i=��BE�
_�&9����6lȮ#�f��J>�d����+�0�t�qtw(��0=-�OO����g��0%�XU�J0�Tp̆l�*`ZX��s�Ӳ{�2� ���9��9ak�7���J�(m�a�&��W�d�0�?t n��O�����=�wC� �Z���^[C�磃�yb��bI�ǘ�Bݗ^?�!N!1��WsH2��0���������6)WŁҗ�ZQ�U��IZ��+JX��]�q���:5��-'��-	�Z�l(����X�X�;�t{kr��I�H�VU �ǭ�$�oy�m��.����8���H?c��9�fH�8E�Z3��;�Qg*�z�=��ug�&!8�`��ME6ɀ�t|��#�*|����ۻ#G$�+f��l�$%R,O˾/�ݾ�T�����l���FE��\&��4��܏}�#����+�w�|ew����'�������_6��W�x�4�헶��"˷����{� ]yG����/�v@��o�r� ��A�x$H�j����+�h��jd�b#w�P��F�ȗ�o:)О<ȱMb��p�ywh��eK��"��������`�M�^qV0�lE��+4�	��4������s,ԾU0��o�Y���Ȝ{����6깾�Y6�禵 g�$�.S�0���̠ �@F�}0C ���N�oH��$�夘'JƸ�il2��t$/�]�go���[b�As@�؉&�P�5�2���D2�a�]�'f�$��$�o�ܐF�G��	ژ3C��3-*,��d�~�T��D�E������X�nɞ��L�@Z4��������1�9�DΚ���7q�=7�s+��E�V������m�3�E�TO=#�x����`�� ��;3��5X��{z���a���c���!��1Z���� }����|�;��k��b�
y�x�|�˟�O~�32�4ŭ�Ƞ�,�ŏ�=��j �c��ˌ��o�|M����6���Zql��2G_��3K'�����֤+�[zl�R�|H҂�3X�ʙ򕗾�{6�� �絮��ٖ���r���e�Ր����?��,�.���I���G�	Wt�' ����D�1(�mN����lJMAB��h%�אc�+i��Ap�H�: P<��~�g3�Ϭoǔ)�}�u|���JZˀK�N��,�h�=r��q�2��tQFA���j'ՆPSp�������C~���#�3�R�d�X���]I����Acv��V>;R�����b�>��%y��@���W��{�I�^Z�q<���3�l�6F���z�+�X*j6�-XhIґ�����S�0��ª�Z>�.�*`�s�Tu���}{��DK�Bxa2���@�~E��
����AV�er�AG�ܮ�Bs-Zz]xa��]�k?������_F�w�ǯ_�{=�r�!����r�mG�َ ���m�����L���32f�_r��k��w�����c{�C�4Չ\�cy�T�4(~t��8%)F�,L�1{�,8I�2R��:���/�Z�����.��qɑo�_��[�d��4F�g�ْ������~�gYo��X$�2aJy�d_.8�ޗ*a왠�:���i?�����_�����]М�5�(]%�.�U̼�fXX�����)����q�� Pl�m�??��r�g���I�#�`��h��G����É1�˙i��Ѱ�
��á�	[[�7��
z�+i`���S��P�CL�Z8T��<۱�
[�0v�g�tuv�b�83���OjP��A�Ah1g�!�g���/�E}�7-H�8/E�nԊ�d�riV~���X f�'�����d�I��#t�����B���؉I��A*���px�4�-��C�A>�@�'�Gt�ե@��UPrgGd�R���it�W�����BN<���T�L5�ڕ
PKjD�5�!�gV�
�A86t��Z�Y>)��aep����Yp�ο����f	[z��]��W��ȯ�ʿ�����> O}׳���Ǥ�J k
J�k�0A� f����ѹ!P�g�J�<�Tz0;nU�a:��J��;Z]��ٶx�V� #���%������^f瑸�k�V&�X��c�S)���TC��R��i/���Pd#��� �.��]l��\��
ڠ���@C�ْ��%)�M�s��&�FGAD��zz���rr��C�=��r�ު�#����I�ӖB�,��)�T�=h�:7vY�C��/���PIB����y�	�Yx��Q"duj��KB�yqj�,2�@���P
"
��)�_Z��Ic}O�i�J ��)��i�W���+Q�^G���8��}�q�H���85�q �-/)r��Ty�Wo(x���7�L��v�mlG �h�vݜ�;S8{��B@�,Φ�>��nE��ָ#�	����P�	ȵjD��đ����[�gdZò����~��,X��:C&��J4g z�=�|N��ߠ�g'��*��Y\��1�L��1���P}
��H�4"[�2!�$���Չ��w_�7���>+�?��!�J�"�ʗc��t!�dM�s@�Ƥ�-1`*2"<>�7���9�3��@ ��M<i�G����z�]\V8���A��+gNImqV�[��+0
c^�A^����A�G��b�p�!�����2�͢n!A41��c�]R��!����7A�!��T#2$X#�I�`d�s��ܦ�����@��̽0�W)�yx�h��ut�xU\%��H�|ʶ�	���5���ke_S��T�1%�^O\W��M��Sd��F�,��M*�!C�@�J���@���<���\�
>z�1�<[gr4,�Ӣ�^�N�O���J����yVM;�GtXOlE��N�U��^��1�Qq��cZs&0����eG�rJϵh��`�T��s��+�ET3��jIgؔ�o_@�q�!�"�BRY�^������>�1�
����w�qdd�b���22pOs�����;;���^^V��
�kܸ��v��J�ҍ3���Bl�Gq�V\C>�Y��B	z��)�(d��TF�ѧ��GVM	�&�q���V��U�2)�pS��e�ޯ�4(��n����ܴ��Hf�c��Jia�r�a]^X��J,M}�F�����2p#�W��J�h��%td�;vF:��T#ù�jxO"�h@�o�s�Tfk�d0TP��+�R�
�e
N�.̖Sa�jV��N�om�l��҇i�2#5�ꢘDMN����d�T2Cw��}�q�3� Ir`xx3��
#@�	�M�PD���.�J��3�VmG۷�v@��o�͍{��d4>� G�t�&��4$��i4�]X�L��R+�
�jx�]� �� ��O��Ǆ��r� {˳%�jY�r|qInmm[z�s ��V�*S��|��~EbI����4�sؐ��GDR�bཬ^|�m��c���x�P�+6$q��W�>0�N�hݻ��b�f�R��l�jG�X�0�|n�2L%�� �� 
R��q4��Y1 �ӈR� <��=��R��Q���������SȜލ�0�O���/e�y��^��\�v��5�l���Z�x�&ȉ����<h�����K�^�u��v� )Q2H*�:�SQlW�����*�ĕ�J�CV*�*%��RII����8Q�,*Z2#F	�D$� �!0f f{���۷���=���AT�\���#�� 3�v�ޞ��<OR'pe(����.�1Bi�%���`0��M�ݲ�>�=��W�]��R���
�
��{����pC{�e*K������]���6\��^i���}��~Y"��į�[�V~h��l�LR�;-�����e���w&]v]�VXܪ�l���4=O��<�
��'>���'O���v��_w���v��-q��=�]]�~ͽ1��	Vl�AJ��ല���`:s�����n�������lk�\+�6_����}�����ƍkn�p�V�Su�Ⱥ���){O_n���Ӗ�l���U�s&��rn���V���p�J��6PS%OJ���i#B� e��Ύv���z$$C�����,�3��6�a�hxϕ��ޡ,�\SG%m��זM���|p>��+k�֧��KUb����������~�����t���a�ٰ;���f�$�������ķ�C�9K��U��l�F��[Y��]U����5o��+���F>�������>���w׉�����nbgW�aJ:B���U���D�_�|j�=3�G���my���x�u�T���c��_��<U�����s ��YN� ډ�.�vB��=��)�~��;�~̵��ˇ3M���Ԡ�{�HL¹��T)�jX�����&�y��I�{�=����/��ٺ��7#���{ޣa~���R8�kw�Bu���ǈq��v�|7��w�Y�m����

�T�sXNܮ�h�n�t��WAYz!8���Op�: ��*7�
w���[.�|p�aX>�ҙ��7D��~j��O´j��~��N铝Gh�C䮞ֻ�Rwk~g~I��p++���U$�C�=vK�0}#�%Yt�����b0VX�	F]b��؉���:���X��Y��)P�ݗ��,ԊT���Lxj��\�Zw�;�}`:q��[�� O�1�|��+I��K�[G@NF>(k׳��Y|�ҙ8�f]t�Q���\��]j�[�u����>QT�0m˼��%ǂϐ��	&z,ւ9
3?lݾ
�6�AM��������ޫ��?库�Vػ>�T�ֶ�:iv{��hwh4��l���O�Y4��ε�-?7w�Ճ[��lύ|�w}P9Z�����'��Ϻ��_q;k�O������^�ʷ���VV�lfDܫ�;�����N��w�u��Gܿ�|�/�]�r��YB�_�;��ۜ�r��I�o+	��V٣����i?q�ӑۼ�7�=�]�奞�)N�djgǿ�VV�s�^w�>����u�� <O���|r莌V���,@�������7����������Ů���������\Wi]^w"��pO��V��4$)Z-Wӊy�Q.�[���[�@��/YQ��:+�V��7$v�L�Jn�^SR���LgD�:W�_����c�M5���ݾ��t������U���$���@������k?������顽��kеs&tYF����Jj,��Tz�zi'+����JP�܎G���d�<����g�`�g���>Z�V���.����n<��i-%ә��W��p:(�r�~�߷�}֪q��꼝�R���>��c?�~���fXTQ��"����|Z(�s���V�ɋ���{��-�hG{��Is^��(s��U�o�ƵM[�H�;]�⺌���;�
�vH=|�ِ����K�n%����O����O|�ce��u��ϒ| �	ޖ�>6[[��Pp��U<�,U�;| �h�x��2ʪ��.�s�_]�<��!X�����y�}����Uj�W*��*��S	�p2��n�w�_�
v�VT}�Ur�3�]�@L�}�Ӱ�:mg-�U���E�P�C��$�ru�`��L�!�PFq�o=�O���N�_��HYp~]�+�P��j��J��Ep�߲}{�q�ou�Ut{p����6��s�>t[�!�5]7q�U٤iu��	Y�i�+yP9���f輈���`�ʰz+��f2�����6�1���yXqUg{ZAU�\���m=>gjכZ�R?�bb�}|{+�e���vfC+��[��"v�(�>���(<�	ϚH�?_��5[̏�Ñ`�+���㚸��O_}�M��mŹ��<%}�1�-���~�5GD��W+�����V��^%_z*0S�͡�5���g�A����!Q���}N�ϻ~u���u�j�V��n�pt�sKK:�<t�{W݉�m�V���m���Otgfe_:kr0�T�y�m��ʤ
ɯ&+�������צ{.U2�Պ~铢�M���!	�d]���v�d�&>a�/���Z���%6�o��f۝=uʭ=z����������5wa�������ܰ�/:S�ם��:-t.��z�lj|�}�\G�7�V�j�m���v\��Զ_�3#U}&Em`��v9�"���u��~���w�������V|h�b��yh"1�l�F�j�$$�;�n��>��~�G���=�����G��?>��~۞]s���YZ_s[׮�.m�Y]��\�l5ng���DI�3��~wٿN��p{����{܊O¶�v]�'ʯ޼�n�,ѡ��:���w��\����b4q�ph�_y�EK6��QC�?:�b��l�*�y��i(����U�_J�s3��2�0�g8q����Ʊ۾yӪ/�?n��'���]��2���>���-C�����Qh�w��+͍)�L6���w���_���?��}�;!�����^1��֠[g�ʇ�q����^���N�f�|T��J�&���<�t�l�A[ET�%mb����`V���E�T��L+����~��$���,ꄢ%XUwu���Je��X	FX�����V�~���>�W8��jQ2���4$<Q�
k;.q�\XuO8$m���-�l�7lwa^�"��ۖV ����A\�!M��Y��,�6cjU��M;63;aYj	�u	N�$_Ղk��V����r�Ú�)��0�� ������0rKbv)X$Y� �S��a4Q�߇��tև�U����y5�$���V�_cK^���}��c�>m��f67#�V�4��<g�5���y�D(�����tV#sj�3�]�ײX6[n���?�ia�Gt-� )�]���U�֪���U|K:f�%T$���x�&�c7S�h�f�5,ϒ�Vh7;�+[�k��ZB�le8�����~��zmK��Фjு�.�&�)����툗|2��㬴�7vvI%A�>���%`�5�9�����M�	�zy*��/�s]���k�����=���jԶ����_qW�n��zb��\+�>�Ga��^�>.�WK}�פv/b�,��p�U�|���gK��G��f�,��mV��U�]���م��Z|�9"�Ӫ�L��Y7�ђ ������QQlu�R[Y�Jh�����l�M|;TI�T]ش@з��:qp�O`J�-��N\��z�����n륫��uG8}h�;��Y��mV�Xh�ĝ��u��Ol���O<��=v����N����>����bd�2V��,�t|��&%9m%�z�}"�(��pvE�Ҷ�2/u���tM��B���.��Y��v���Ѧ���P����[i�o?���_��_s�N���?S{M�)��3��v�{���T����qA����މ�f��`w����~k��^�8�W�wE�����\y��kׯ�-Y�1J�E*[��|4���M�N��ݯ�0�>���v�jM�����lTN�Jn&.S��0�\��H%�
��ܺ�h��fWT�J���H��>�i'UV�������@��psU���9k��
}��X���]����$�%�R���h=3�J0l��(|�/΃��*��f�B�B�,W�!�(�Hp1Ua%7�9+�p�ݾ�+��a����>���}�}��"���M��'�M��I�8��Pp�P�m���9i|�1XiƼ�s&&����|#K�NX
p�VⱿ�_O}_��a�v�E��(������Y��t#ۊzU�����KAf��K�;
���HC 8���K2��M���uR���N��>q�&6�B��YQ�t��<<�
������J��c�i��">h��R�k��ˬ3Wa�b�j��EVƣ�06�!b
�X���w�U��+@տ�B�9Q)a]j��Y�����Y�-7��QW���إ�6+7�BK�$��a��O
��6/Cy��*�R�Z%a��#�*������LS��?'��=�sD+1V���Yv9�zn� B����e9vT�.m�g��rd*�S£�#=^�ܥU�N�<�q��r���m���jw�t�*4��t���_/jS����?n�{��}]~����c��2�Y�Y;����?v�-�wv]��d��Փ��^r���
�:i�-����L]��s�V��/�;88pǎsG�U����s]K�f���.�̿W�$|n(aT)`ZO�N'�[�/�A{l�ķn�rg�u̝={���>��^j���<��f�;�F�Ϣ3L���F��g�cd�I��e�P�v,��5�=�a8�b8�g��U+kulaD��y=���?���q����n���ln��0�޿cz=K2�@��F�L�pNLI�BYjt;)��|�k;���-'�Q�F�.{��/�/��S�������H@����V{���[׮�~�#q[+�q�ebe-:xy�]w�;�$�y��F����
���:��m�nҶ��|2��ҚK1�IF���J�R%�ЕE�S���C������t���λ��Ⱥ�ԉGieL���JMG�����o�+"�+��(�벑�g픵��$�^�]�����t��|'
�%�N�
�Ze�tq�C+���6$/��M��l8ȭV�t�#]���涃�ݦ�����՝/V-�ߣ8�r�)�*��J��0�&�ۮ�J��p�B��y�����AKU�f�$��V���<H�[9�vt�[d�5
�`׉���4�^��swlI�칿�I(m��V�r��[��ܚ�O4eU���X�i�l�4�m�Sݴt���������^���tjgN4�Ɔ��˺Ad���j���~8(��b���F�)�!��uVk�n���gs���.[V��Da�������n9���z)�`9	��P[�5%0�-�u[�Ե-���A~����8ViY7���U��Y�v$�+�Ht�x���Aہ�2�X�����T�V�~S	�{mwRM��j'=���u�p�u�]%!E]�cs%�{�]_���h�<��w�%�����T?Qײ��Ρv��\3AK|�*��T�>vl귳��:��O&㉽���������O"7�;�^3]���Tt;ն�f��&�Zp��J䔤̇>��WJ���{%���J��c�5�seífk��O��#�O:�=����%������f��Թ*�k�������m��O%����p�Wo���n<�u���Y��5�IQ�n[������ݰ��^��#k���Rw�%K>ٞ����^�D.6b�^ԕֹ�v2���=3j��̕�Ν��K[[���0��V��d; �B-$��\�&lI��O��к-�:��,�LM Ν;7���t �	ޖ>�!�q�J^<��������˕u:J���aٍ�xk�0��:nU3>��M����9T��K����G�������0���|�Eg�����u�J, ˵�\�J�U�*��q�$�k���K/��w��b- C��.�E�g�ydt�6�÷vR�
%=
L+W��s$j�8�m?������Ǧ�OҺ�$�"U9�ڇ�H��V�Z�W��S]�dAp�x,�T�3IJ�ֻ%�A��R8��YkWu���rꃭ��Zx�j���J�T:5q�<��R��I,YKm�WZ>P׎�tV.U�b�G��~���y�W��Py�XдҾ�G���pL
,���cQ��V�VU�`��P3;ScmvŦV&�h�6>�nBlg`��d��Id;T�:k��U�ý��49]���x�g�Qf�H%�yJTT�e���5���]s��y��D�zh�{%��5�t�uJ������E8��*��5�QԶ��5j2m���ٶ£Vߒ�p>ȅ��ڼ��L�U� �JC��o^�� ==�c�:.-)Qb���ĢR7�2��ց��ZY�o�M�ٵ���vԶҬ��O�k�ȑ�n��-�1����h>G>��Qz�J�&Ӽ�v�BR�\kwNg�2�`S�-���맜�u������Vl�+��a	Q}�)�W�v�H�p�] '���,Y����e�:�����^�De������ދ���-�����t>bg䯃����w|u�v�m>���Ckf���s��8TZ�n}iٿ�|�0�w�͑�)���-)�l�C�7�{ށs'N�q�n��Gn��ω��n�v`
;=�z�dd��E�>Y�:t������ȥ�y[�gмe;>�<4׎^��w]����Q7��ݰ<t�ɝ�(g������~NF�3`dg���jo�r�E��8�g�Vu��c�3�����Uߦs[���pW.�����������v��׷�D�.�Έi���s��P�;y�Ij]R���QT���=����b���H@��w�����/�k
o��/Z�n�k�����2Kױ��"V�@Z����K}��/͡�#�l���&:�ٱU�q5uq�ت�V��կ�'�Vn���W
���Y*�;�%W�ۓ���(xTд>H�D��
Z-8ʲP��h�|f_(����g<���V�uܺ�(Q(��P��P�a��|[I�J>��xF�d��1jV�U ��J�Uv�v�Vv�����P�G6pm6	��*���֎���V+��֣�d|@��wl��ٟ��_˩���U;����Y����ݧN��6
�uHY��X%7I����ӐX�1���Z[O5�0�{��G��(*՝��ZEX���skij%2V����6�{��:M}@�	�MΈ�z�sۆ��Β��$L�nE�|0�:���R����i8����k-�v���z�^�*�ϭ�g���]='Q�����J�p+h�=��z�M�V«�y�X�-�C�UZ��b�T�&��oY_����$���
���$G���v���A���?���;�����3Z�֎��*�t�a����*Y8���I{�����f�ٱ�`����]q;��p&m�u�Im�_S�J�����~��[�� �X+a�kǦ��S��E��hU�Z�؟�Nִ�<�QX���Cr��Fu#
��'���Yt���g��:[� |@�������Ѝ����0Ǟ%�z��k~6��z�Twv��A�׳R��'����-g=��,������u���u2S�����V�����W]�w|��˒OS7(�n_��[awE�Qܺ�2���5Mf���n;�2f���I���O��g�C;otߙG����_�F�<�_���P斅&΅ݺ8�]ڤ�c�'J#�LjثClV��:%�Z$��z}��P�U�s�5��ܒI�מ����ݱx�f��*����䱣�~�mb6���Z��y����fWa�㛿[nw��1.f�S����w�q�Fy��n0X9w���H@����|�i�;�6?�۟p�?�[��+t��뭹I���Q'�ԭ����X�AHKC��Ҿܦ�c;������}R��������_�?��Ȇ\wj��$$�G�m���}�-vET�T�3V��)��d�������҉���*�p���=Z~�E��tQ������A)�Y�^�ceBZ��}0����V�S�UX��@��LU�����>���й���geI��:Y)��WU�_z�>;0u����(poյ�����_tP\�.�V�|���%Vo%wV�퀮:�lF����.�*���ZX�E�{�9�B��J��DE�����,��)a��Rॿt}���p(�P�����G�q���66�.rubV��g-aP05�ڮL�_W�:.�(h��v���6�-��O��2��Ά!�r�����u���.��~�FI�V�����9A�nf`g"����u�Y]f��CK߹uxK�~��_]9���|�jn����]/��~ּn=��V'$�����$��.=^;���R1�ǚ��
m���z�5���'^ڡ
	Hj�2E���O�u�_��J�td:������oɅ�E���{'쒨WU�uk�8
ϡ�#6Ϯ�O��:�3�oI=�I�2�[=[p\�������C�����[�\�����������C���v.qu�����ݡ%'v����1�Z�\�?_�>q�tԭ�:��U����~��?�ڰD���I�v>ZIص�m�3N%�
��M����~��h}���DxO��ϵP-Z�DM�Qx<i]��F������u���v�l�T��u�I2�dB��[#��:���ݐ��TJg��~�5��>;��e���k�ew���:���֎���[�����P`e�Ӽ�����2$�q$u��n$�H�fVZY��8�
��g���֍�������� ��Uu�����KɆZ?v�V�~��Z9�����qT�85�Ck�č�q8�� �V��jUP%�.���G5��7)0�nUu�"i�
f�W� ��A�/K����}�|[�����Vw��Ķk���es8B})����n��s�Ź�V�t�z¹nO���ܴ�leݦ8��$5�DGa��a�{��)����U2���V1�+��R��ጌ�QT�rHB�����'�8u��է�<�iСx����Ga��$�gX�qU�Oz.�+I�ós+#��A���3*q��Ts������38.�f+���8<<]�t�[��iU�:_%��Ll�^'h��Kʖ=���D!h���up\w-か:��H���d�:��J�v�Xڅ%zmZb��	��lI�%CbU�����R����c5PX$F��-ۥ�����6�S톣8�׺RHl#�OV��Bw +ﳶ����(�ٓuI����[-��";q>9XQ��|�̈́�u�k�}�?'�%�J(�Rs����լ�[�[l��+�c��q�#��:���0��N���~OX��$"Á��Z�#]L�&��O�bK�(��`�~��̏�w����t^��ά3Sb��eI��.GB����{��c�9��W���k��IVە�:��kL�yz��~��f'ՠ®=6�(Xo�ܞ�%	�+���H6%��v벦��v'�������J�GC�����v�ev7�����`f�]����֘!|�h�����F����ټ��C��}�g����BDV�՟I�]��O��Y�*�N��ܒ�貿�j��/���ά<p�Y�q�t�7�,�3�΄�p��M?��?��r��F8�n��-�!�S���Y�n�l����~ÿ���'��=�-���m������<�og���q4-������7�AQ�N���J����u�s6�����U�����l%;�R }�*��������L��ű�ZI�D���־x��JUʬ_��g U.d��J>�;e�@ab��ʴ�p��۰�z��J�VZgo�a�������Ô��n�Iª��P�pv��}��>�C�nN�Tg���/�!��"���G��+�!��2}���S׺�����XeU��:)����U[k9�����p̵��i�:|[w�r�MD��+����0�Q�E�*�O	-pC�gA�J���ReDv?	m����j}�!h��V�;�Z�scI���Ow���� rf�� C%=j�3>(\�;�m��C���S���u�]C�"�NI��@v��C�v]J++��Y�݅0�"�]QQw�.,^cV�4��,n߾���}K�3��4LI���a�vߔ�p���f�,��A��G����
K6l����S�|��]K��r��Ν�ر�=�S�.z������������ܑ^'$hE�$���d��Tڮ�r������mN�������h:	�+��:��wui�^,H�vT�����\# Rr� �zh�J�ey��BhWC%e�~�:e�'C+�����k�/Ť�F�>�j����K�m׽۱k��W��b��PiT��nfծ��I~���{Qɚ>����m׻;y�Y��i9u�ihk��7������gV*�ܲ�ﺦ��a�  IDAT���]jܠa��{�v_����!�9{��S�ψ�"�{�D����0�9*��j����YH�R�uҲ��٬��*	�R;��v�*��.��vm��*Y�g������=�n]��.���^9Ž㡇���:�9f?_�%]3͎���Y�������qI�h�Q�ykH�_O�ۻ�O������o����ze��~�c���m�(����r�Y��~g��l�c�y�����˴��>h�1j[�F;L�C	�Ml+�:&[�iYw�R0�\M��%�^����M��2���+�Z5�U���Bנ��eV﬉iHd���{P*@��}��++,�_���+��'��Ir5�u\֝����4��+��S}���W�v/����mi�����d-�����C�Tk���v9����� 'I��@��^��s�����P��
-}Gc��U^��
mU1	S�GC�'����Ӌ�2���p8��zH���A(C�MK�A;V�&HG0d��;��o[�n�QZU��f�4��t'��L��)��� ���[!Z�G�kᯱn����Ӽ�"��8�|�:/��I'��5(��,�:m�Vij�
�8F��Ϭ�,}���s�&��X�Knzx��E��&n2�,ĵ
���`Q�d�7�y�Uc���I�hw�W�:��I]:g�}��4�r�"��t�Z;@�y�H�y�0�{⯙��n�?�Q�w��.�����*�;q�q_g����{s���Ze{�>?i��1?~��_wg�+VM��ݡO$VW���'��o�P���:����iQ��Iv(�����-��%y����Ɩ����~�u�B�������L���C�|K�:(�UN�ۿ��{]���eM)�M6�DUޔXY�����
^����e�{��c��LG�ri�Φ�z�߼u+��]��x�vwv}@��N�:U���J���m��y���OI���S�N��G��i��.�:uVm��ubWB���=�*�z=���j���7���f���+���w��ʈ��B<�G��$D�8�,v |���9������b�cS��ؿ��D��Թ�L�����r�Ñ�����ԭ����^�?}�}�_t;���Xւ�=z�;~��v4�%�����[����{����,����O�����}�O���M�j�o�h<����݃/��}衇�i1��ؚ���l��_�.��v��;�����r���j_�z=��o|�?N?�$j���Ǐ����r��+�����%
r��s�.^|Ⱃ���pn� |OH@��C����Z�[���2Ϣ���ɴ�b:��V��)Vw�tT�T�bͦs��T����r���忤3�e5OUm?G�gy9)N���C��Y�*��_\.��mu��s��>���k�D"�ke���a�[���z
�|'!(�Ѵ�O�Y>�K��l�J��;��*I}"d_�-�����>���^��N��>#�i��z��7+�|d+��,�OE�|6�:>9�2�}����NV�>/��
�Zj�o��2��� D��*P>��U�p�;9<Z籥�r��-�����b`�ۚY���K׵Q)�~~V'0�=�:��'`Z����{�E¡`u<����} S�|b�$M���]��Ck��b%"�y�ƺ��"냕��z����>P^uS%�P�Z���M�w���E��K/��*�U�y��b� |�����w�ݽ=�<Q�ol�N��b��R�E}�0��A^�\���7ol��>��5X]^v�����>��zF;{aފʂ�������۩K����
l���W��╕[ᐶv3�e瓿��M5߱R��#�����O�����v|��K��'�t777����B���>99v�dy�ȑ���C6}�_�rww����+���ri�Z����.�\n��o��O�����v8~��-���Ǉ?���땺�/�z�}�����<�y��>	�]�\���ګ�ҥK���O�&J�N�?~��G>�{lW_}�]���ѣ�����~���[���[���׊��0��u+~��Wݍ���ڦ{�����g��C����K�y�JOƧO��כ^;z���v����d�b{k+��ߏ�rd툽�������#�{�z-�V~7W.�_
>Y�	]y����ŋ>9٧�h8���K𴋢0m��ŏ�����{�M�+�G��_����|V>�O�=�̗�Ą>��sYt���ܹ�K��(4]�[��pJ�4�ӿ?������V�ۋ/�rɿ��Ү��(�"�����O5\�+K��������w߽�P�}��󉩺��n��Xݺq�]x�|�]�������O}�S���$M�C�k���¼*���i�?�f�������a��9����<q�h抃����N~����l}���}�(�/N����W�V�?�x}r�w��o��s �C����գ������/�����=�v|(��൜�slP�q�Zć{��Gk�C5�>6�u��U���wgڙ�~�*V��T����n6<��}���	�^%�J�S%*���~��QB�Z�j�����JOsT��6n\-Ɠ}����|��_u�N����R����x4�h�^m�J� ҋ/�Ky����vz��K��W<����_}��}t~��G~����{��]��чz�\^ZK�����&T�����e����cc
�e���}�����3s��*�pVVI�׏�Y���mK�����~׭��voT����wO}�s>�V�Z��vy�����J�=���IGc]+�<�>�,���z�j��?���engw������5J�t��g~�;}��w�| jA���?�o�����;q��][_+��������ӟ����tum�ߧ�[⸵��| T'Cw������G������؏�<̒K�NuZY����d�n�����K�Jb
��ũ�P����
�U.t��i��=��{��l���<�0�����_�:�i�����`eD��\�'
z�R<��Y	��g���;;����Ӫ��766�u�v zݮ���	Yٵ�Й�`P2�������v�z����d���s���R����Ãrooo��������v��߅��$�O��'�Q�fQ���x��v��g��E���;,�C��������Z_�'?��v%]�L~�W~���r����m���qA��-�}���C��_z���ٳ���}�?�g����n���I���̓������d�VW!Z���Y1�$�|�Y]����ټ8�/�u�_�������c�^��Y1��d<ɒ��6�ײ��U���Q���U�l�7o�h��q������)ͱ���|�A�.]����~e����ۿvg�;�>���H?g�ڋ�ףq/O{�Q��S��R�t��j���O�V��d�u��mm�Ҹ��No6_�ܿ�f��ٜ�;eB���>W������~�7~���	�֒��v�w?�����'�j�=���Q��_�} T䳑���Z�m�ri0�:�3g�O���/}��:�~P(��v�J�|g?{��p_~�����@��-�L��N6�|<�2�����^��ZKPP���ɟr'O���N�ŷ6o�SU9<܉������w��|`<�}P����ر�Sg�N�u�>����=�fJ\VV��v+�.]8?���?V^z׻�������˿=]��mA��_����?�;���Џ��$�h(`���U���A��&�_y����˿�����_����_��6�r�^�vO�����>����x�/�(r�(z�����\��Μ�������_�/y��|6��ݭv�����N�s�����U�<�������|���yF���Z���J���es>��[�7���P��5sJ�V5��K���/��j����'s��L�>{�֍7^�qk��4����[ݤ�=�6��:����#7߼yk����t�����|�/����VVVutPd���ͽ������իo���p�°�3�k.�������ӫׯn�߿�ů��|�[�|���n������^���;������o������z���U&1���C,꿾݁;toetg�����n}��~��-��s�[+���o}���=�;���Wߋ?v]}�*�xѽ��j���m]��������������g�9�" �W�ok��/��=�Y�����������Z���֏y��7�<��v�D��ǏGY�U��4�\4�A�����{���3��~��>*M�YU���+�'?���\x���|�ʥgN=0��䓮�Ї>]����Ϫ������|��g���IZĝ��7η{�����n�W/�^n�L���\���i���A�W+�9���t��]w����Sc?~o|W����|���?���駿2�ԯ����{���~�w߼��V��n����������޿�-%?��u�����I�up��q>����g{�֭��n�3o��+
���k�����[e��|P�c��o�L��u�=�Q�r��C��盃��-���}�C�o�;�;;�o���֡{��o�����.J�w�㟖ç~���~�+�ï���`��~���+W��t��R �����z��g���]��.��o����N��_�>�Q��mfW����Ӵ3�IՉw��g'�\�/�~���YXڼ���g�_s���	¹;�t�nm��/���?��;���9wn��������?�G����{�?~�t9��5)��K�3���^y��q���}�,+��eݫ��ǯ��%x�W��$� ��gH@��V���s�밦������__�������k����$�/���x_��ck���6?���q��  ����s�~{�����ܼuBs#��S�E�j4^U��,�ˢt��V�t   
H@�?���re�����Ã��vw���cǏ�ռH��&���r���,��   ���� vU/\|����O��/���o�Ϳ�{����F�I����R��g�q����9   �o�� ���W�^�Ї����_�_����W?��t��Y�ǣ�ڭ�g�8~��͛c  �@�䓚Ip�K����   �?D   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     C   �1$     �������N    IEND�B`�PK
     w�O\����  �  /   images/32487380-bef1-4e4f-8e56-19d5eed1120c.png�PNG

   IHDR   d   K   �"�   	pHYs  �  ��+  ?IDATx��z	��u���m�{v�&�F� ���X�$��䍜�8�q�	�c���������`��!�@��}C��3==���Z{U^UK�����Q~����F�]����{_�8Ԣ��H�E�*� U5@�,j�TY� ���ReQ�ʢH�E�*� U5@�,j�TY� ���ReQ�ʢH�E�*� U5@�,j�TY� y�غu+n��'�j*��0DIDYqՆ���=n�����5@�!V�솦�p��j�z���AI�&419y���y=w�wQ� 8�(�K�n
��갘[\�����m����O��1����E�E� �*3�z}����=������5@�!t�"��y�����o���b��i��B�>53!I����[1)���ɦ����ïb0��M7~�]��� �?~���6��.�p-&�	,�l���Q*���Ҋ#�OaUW7��uK�ڐ.��0��E,܈���,�{{�ʗ��֊U��P�%Q�����g�T߈��,��i�8\7L�d�~t���G����(�!���w�8��&b^��"��˘��XP���n��~x=����ת���i*&L������P?��O�:�!8�dYzm|rdgC쪢^�c���x��߼���;�pM�:�l���g�8�Yĉ{o�l��O�.���z Hg�����Ɍ�����8.��:�3��|k���������i��B��e;J[�\\������q�
�~5�~΅�v���=���_L��67m���э��0�R��c��o<�L���X�ѡ3��n�0ݦuH���4��_E�Gs���[�lyd��c���>�/�v�o��C�� �W�G�~�'%��JV�J�޿�!�e|*�0�BQ,��1 �:�:���Id�]Hbm��\��|y�����gwe�j�o�	p����������U���3�rI�l�{�e�����X���z��)��VY��j��;��ii����q�|��7�hJ��ϽE9���:hO T
�������ȤNdi��myýT�]��w����^�����(�\�������M��������O:o�<yC��,[끫���O�����k�Fu#7�#@�,?��d⟞{��!4j^:��a��ñ��WR�/�xw��ft�~�+��.�E�:�Rzu�r�$��V�d��2�iK�i0t��eX_14����)h����i0��2�J�u2���)ϊ�^S���d�U��
�*����z��x�A(����-��}��om���S��� �6y��z��F�����x����<�Qn2�s�(2�8���9���֎��b]�%p:�B�!&nXqֵ_	G����CpM���B,q�A�g�ŏ�}+6 ��>�rr/��\�Ԃ��ݭ��e��S��h�j���Ď�����$�i��D���57���(kM�X& L�V�1�SI>�T�ku����T:v�Ya�����=_�FKÒ;�=t'���w�{���_�(���;Eo)+�����WZPW_�T�qd2E�OepL41������vz�9��ٸ��F��(�������p�+�!�3��.��֋�'��U>,o����F0w���W���0>��[��Gf,S�%-NL�2�y�*�5%a��y�F&Y�A4@��FP'����dͳ�O5O���Ǥ�:��g����]#+*\d�9�.��s"�~���?�t���v��?�ݻ��m_'�3����I�6�(�f'͠�I�E��s(E��+I�ϑbA��;ծ�O�|X��r<£��Fɥcq�*����%J(S�N�M_�/���*��)�ٺ� )�q�d�@h/"�h� I@R,"/E�+�H�P)!��9�J�t�%'��cΝ�f�0�a۽1�6[��]�p�}�O��D���P ��44g���@T������ ��,�2, �n9KZ��8�d��3����F������k������p\��֯g���Z,%&Cg0X:	OÐhog]����x���b}f�����C��Yo�9����P� ����uG�"��.t/�߿I�N�oߦ����aӕ׀����ObM�j�9+������S:��C�X־�K'(s\���ќ	�Ak�1<2^����d]�|~���ػ��$GQΑ�*����M�u�<vn-0,PX�c-Wrn�9L��N�苓���Siu���������-t�}s��y�{���G�Cd�g��������Y�Q����.:�~_��
>i!�*�Ĥ�%]��=�G�<��w	-���~ja�f���G�#�e!�*#(0��wkv�H�9։%��CO��!��ׅ`�*�x�!K�}D3=c�Q�f�о��kE$�\Z����XX��g��_���N��f�����#o>�2]��/�DN+X�A�$���h�MC %ڰ�ܴJŰ�,� K�Uô���	���4B���a�2�Sx�_u�W�\�qy������7�P,N��OJ�+������p��ʥ\N�����+8�W���O@A� �H�*�Mp�M�I�i� xx���0��US2��.ږ�T!�#�Q�~�����
~,�rH�4�!��|�6����{�(i&.��XA]|]k��鈀#���`�(!;'�&��f5��,mCT�8ζ�紁9W�8�lQ����z�u��+���yhtT�d�m���d�8����wb��M�"�J�����4��;ݶ��@U0T��!mcQ�Ėm�/�K�Z�s<g�E�&^���g%�nlZr!±&5M�Y�_�aqr�v���Zsљjb}�~���k)�;�Gq<Q���������9�%������ �O�χ_B���ӋC�xq4���[_C�R�������d�0ZB�:}�If�c��"rŢ�+ن�۶��N`��*0�kZoP�i�h_�W L���)�Bz[�)�?���On���b��O7�r���Y�l�TBa�2I�v�h �'ݤ*�,��ym9V.߈;�C�<"ݽ�X�ᒁ�/���"!��(S�R4~��Ʃ���n�M/��� 3���A�L�����C�t
kISt�*��xW3/�a�8���<�Ewsf:��
��#���9��{���=�2�����xr�'Z�T(eͶ�%Y��ie¦+[��n`�V��S�ڭe�G'p'o߃fX�fmck�,IZ��wԏw��h818��������vy<>/O�8BڮZ<�:�N�T��x�$�2��8��#��kr���G��&+l��Cq��|uǕ�vϟ�ѷN`����&4,�D�h��A�j�m��nq/�&��٤�T��PP ��;3����%�p��� ���]�a�"ܒ��.��%a�!q!]Ćk���!|h	.��r<�诰��0\� 2!�IC�� &ka��j+��%g��,H6eY�)�%�,o[�s<c��Z��w�����?��;�:����6����}s�O�5>:��d�l�>d��q0���R.4�2ޡ<7p|��t4��5�v e�1���5�Q��s�1��#�"iF>.�u��G�DQ�ЗC�?�i=	890�-��Z�['8�A���K1lC�'�=�)?=B�>���vl]~5����0q)��g��`f�8�����c\hm�ᕬva	U�f�:je]�(���-bT�����9;�Е���az�aѦ:�V!���ľ7��W\����C���o����4��E�D�'d��)�P���ěz�T�)�J�C���K1\m��w_ܽ2ւX�~���~<7܇c�q�R;�@Zq ?���lD?��%�6�;����/�yL����Uh��N��d�&l�N�ۇ���ͽ艴b}^"{+G4�d��OB,Q!t�ؓ�307u�덧P�U�gql���i��9Nh�˝��
 �N���\g0�:�4�YZc�����@�gpd�хt�}�+��/~�=v�� ˶+��%;� �h��8I���yuΰ�j��������{Q��/�6��(�A�SYȂ!�8�0
�ͥ&l�=6]�9�G�`FI���2��t�n��i�U�vt�\@V����E�z�DK�g
!,�W�L'��8u૙)Ҙe�Q� 
���GS3xa�����>,92��RXE�# a>7��Y�?��/V�Z�P���ه�T<]�A�aZ�eZ�/#�J?p٥������M7���;deW+��o088�6����َU,�U��d)�D:1� U:+8+���s#��cO��b.Z�	�-�ċӯSG�`hZvY���pEN������'��՚?��S/���%ʳ��`~|gR�p�������@f�4�Ijs+ф�0M�!��X���a�p���td���RWOu��5��&�I���t�Of�%�R���T\�X�P[b�� h�M[�D���]���8������[o�OmX�y�����~�/m�����O������ï��Nv��9V�4�e^p8�
VUزF+M��K�l��w�yNp2���#;�.���b�4٦2gךi�I���.�E����L־Ðʣ��u��N�'�p���"ǇQ �O��2 �%���M�p�����@3��j#�z#8�wy�G?�IW7�}#�i\�7A���o��#y��L�x�O��Cﳓk�b��fT\��Yd�����)k�7��v�b��+�رk�?��9�!�ߚ��	�������m��7[>���L2	����F�1�N,��Z�:�����,���b&�����C�'��m�4	&$��`�!2%����SJ(�q|e��~�F��'h�5K��e:ZW �ۍ��}:ڢ14�w"�"�1��a�wu��"���P���.-H�'�6�}M��!I:�ӻփ� Yُ�����m��n	�����^sc8��о�Mkt��F�AB��z�{�E4gM�t�i�i�1gr��/����+��^u:]x����}����eD�u����Ï��g�Lg4F6x#������|�UDn&5���Ś�!�r���(����u�iQqFN�j�8�G
R��+��~�p����Q��� #� F�H83G�����S�+�ǔ :���[�h�	�ׅQҤ�����w�u1(����Ip���x�<i?\,�f�����.0+[�m��q`\�B�s��������F&�4���tɊa݌�(<�,��t��t���AEQw�8qd�e��?p�F8I����`�+@ls��2�ړ�
���D��BW���n�5�VJ9t�l�w�}�u��3�E��Ѻ�3��x�%��FTY���zPI�M�����+�b��h�����`D'� 	Џr��LS��4�����`��/Z����b�4�#�e�dm��l��R(ۏb<�2�"�f��t"��˗a��_���� ua8�L��\&��ޝ[$	�TZVe�P.�q6'�O�◚(�����tw�@(��������w��#�c�����8q,�d�����4Jy��z�п��Ƿ|{��k���^���cSTJMc���������a4�ppY���*�!Q���4�	���M��ؗ�o���
%)S�h9Ļ�.e�h,2j�<Yn�z�-�:9���F;�:��^�_(��=ȭ�[�i��t�@��e
u3��>�zA�2�NWv1�������?���Q�����)�H#֒���>�'�$F&����нb�w����������w}У}������_������klsĳ�xC��Te�t�<IGʐ�5��`�X�1�$��%�33��T.y\Ǵ��˴.���E���/�!f61�(u�*�����'��t�u�CƠ)���&�f$#'��'��u�,��*#�L��W��Q�ˢ��<fɒFG�.�CG˭�mE�g�=�����ɑX��g�E���U���w��z~�8/o�hX`t}���]��،
��C�[Q[�K���b�?���/�;q�m���^&
�ꇋ��8FZ�H�H������_a74/O�L�j��<4G���irT�A7؈L�M�Qh_2 DX��Ay���IG�f �����x)�%MN�Yp��y	D�}h���l�]w܆����ߏ��s�m������������ G~�k�r�qj�<�=;���W]��Sg��{�� :p�������]�bQ�_Y{dd�/�y��[c����{���o���x�l���:=�����OI�,j�TY� ���ReQ�ʢH�E�*� U5@�,j�TY� ���ReQ�ʢH�E�*� U5@�,j�TY� ���ReQ�ʢH�E�*���$�{��     IEND�B`�PK
     w�O\��=Y3  Y3  /   images/3d684ffe-1f74-462a-8eb5-42254bda90cd.png�PNG

   IHDR   �   z   ^0�3   	pHYs  �  ��+  3IDATx��}	�$�yޫ����gvf�.�]KR�ES�)J2�@��6GQ�D1d;� 	� ��Q���`ٲˡe;�%ˎi٢�H$ER�E.��{���\=G�u��ޫ���w��Hϼo������������l���1�d��h�jh	4Y54���CMV�!�&��Ɛ@�UCcH�ɪ�1$�d��h�jh	4Y54���CMV�!�&��Ɛ@�UCcH�ɪ�1$�d��h�jh	4Y54���CMV�!�&��Ɛ@�UCcH�ɪ�1$�dMǱEo�4#��aϓ�H�{���A\c=�7;�1����^"�Y]�xSSS��Q�����!�	݋Hh�_cϓ����3o[�v��ck###/沙+g^~��v�1����v��|��1��o}��~���
_�q�͛���t��D�u���
/]x�)���0.F[��j��d�<z��?���������7ۖi���糙z����A蚆��x��y޶������w}e��������(n�d2y#��qmQء��H�omn�������w�o��¢X]��#�F��0�Y۶ɾp�82ba�Q��,�����b�3ssO��^[�����S~К ��6�(��G�{����/?kF�ؘ���������P~}�����?0-�䘆�c9v�4E�jt�i������=�!�(4Y��][^ܿx�J��k5槦���8��]��{������	˩.��M�2���!��n�V�� ��(�a��"$9�f��V�h�=sf�r3��7�5
��ׯ]	ifr|TtrQ�Y�i�F�T�f[\�r��J��7���j�skc���Nk޵H��ʊ�����K6�Nlll�f�-,���(nw:�Gk[��Ψc[5�E���@���Q���������q����W�/}��n��e�8����������P�v�,��@y"�����,}��=7�X��3���ju�K�W^\�x���7�G���JZ���_}���{O|���כ���M�A�r���\�	�"�OOL^΍T>u���>����k$��Ì�c�D����8��,��댍Mq�>���=��wq����\(:^�@��Ѳ�T*bss���[,3�7.�Q�u�"F[��Ҳ�i�7�Rv՜��=�C�Q�2�^��;NƵ%Q��r������jL���|y{�2r���f�ˊ,��P�DwIV�}�����������L�N�j��P�o��A~�it��bi8�|VE���l��������d�x򅯯���V�q�d�_����Y���C����|fñͫq|!k��\�V�Z���_��v*��[�a$w�pW
)� ��3��,a�F�Z-�����Jqc�[�gs���|��V��CCFd;nUׅ�@!EQ��9W�զ��"|�puu�i�6���|mc�mX���dM2`�D��߂eJڹNG�����L#�v���ۭ�h���{�~�Hof#X"�B=a�n��ܚx�ȟ�Q�FZ��\���k%?�.ُDA��:��d�N�=�����̪��3���1�����ٺX��8���vgL��+�8��}��''��b�P*/f�sbcO����ć�����/���2�*��J����	� \5�iܷ�B�<{��k��$��ɯ�}���>�P7�§?����Tec��6�n�-h��L�<�����شMǽ��k��hy�7��y��o���k�_f=��?�m5���Ƒ(�-"� Z�B.+:��0B���ʦ=={�?gsş�=ólVb6��ߚ$2f�jht҅d�J�F.3���.-f��q�˕���?��ZǏŗ��G�K��[��j[[��D�H]7��,������Z!_,�\e|��V��ԧ5��g��v��nm��c8߈Bi]��#��m����X�Vkf��������_��5��٣ܟ|�L/�\�����P�K��a���W��ճ�a�xi�_�p�����l��C�©��ˇ����ܚ���Sd��G?���^x�Ϳ�k���Z/Tf+�B)$n��5i��e���p�'���IҔ�H����ˢ�mJ���І�f �#���SH�e�1�z�1�Vf@	*�k2��w��1�3�B��/�t�N�Ρ��0�A0�3�xa����z�(�/}����� )�nY"M�c��|ԁ��.d��W�~��4&�i��DO�	�hd�����z7�?�i[�pO{�ߑ��{-�Èq�^.iX�Ѧk��m�C���e�p��e���Ç�}�C����/Ɲ�إ�3d���>�Ϟx�{Ν=��J{9��P3A��FBb%L=B�w@@d�9�����l��vbI23R�[�<'�U��m�����k�������l�%v���E�������]���N��F�7]���1�4�߻��`���4m;q/�A���^]��]����]�O�]�{��[[[o#�1B��.�l�&�\�+8;	�Ԯ�7m�����'|@��R aNZ�cĉ_|s����'b��	�V*J���y���=�#P_��"�}����lv�����	���IO�|�����!ݧ��'�aJ�4���?��z�H֏%v1�YO�>]��'?9$��%	
�lz
7ZZ���'�,��&3�aX`�w���+#�b�$=B�	�&J]�"P��4�X3�T.m
��oP^cWs&����`]�a�3�:ԹVR�=e#��Df��nw�����J?p��ٳ��υ�f�6�n���f$��hZ�Ӥ��(!2��8H
�q��s�isU
3�$cS��}��~�<�v��b��`A�}�O%�����������U�&�4�]禃J?���r�uC[�A�fu�.Ʈ'+i�92w�D?�~$((m���j	�A����UZ��$����y8h2Q�� �*VL>q�#3 ˉ~_�׮�;�.�M�,�A+ f'_�NZ2��t��]� �1`�&�N���]�g����GvhP5s9�;����ɚ�X�$�!ډ�hKǱ�Ϻ����M8%��Pr�\),���B(Bɿ��uYd����jHeC�ȱ���T�YX���R���{�I�����dO8=�RRa  f�+Mf��^D��N�b�O�SE{Ӑ�&1�a��B��޲����Z��avO��@N/a��/v:�6���Nx�H*ET�;�}��4v�B=��7?��\*m��(���s�~q��:X�xz�HKm���H��`4��vީ�����Y˟�����A�E�蓌0�0`r������@�(�N�"v1v=Y3���2W�7��f�i�����,��O.k�� 	��fi�w�/�`�W�?/N���$	���~�J�<5}�k��Ï��v��=���a�#
�w��P( Z.0�\���vd�ar����Qte�8�<>�Sa�k�{��#��@"lBNJ�� n_O�����U7@��&�E�r�z�ҏ�:u��$p$ǡ%#���@��?��ϝ���y��>l����oԔ7���p��2�U���|��h�R�$�9AB\�Q.��Krr%��ϭV7�����z]��qN�t驘���X �SKJ�P��i�&�N�(�9}�I��~�P%�H+%&%��X`aד�"+"aHp,��ApY�d�D���LVc��A�A����q�/E�w𜴀x��Ǻ�\^^���WE���I�^�tIloo��fff��Ą��ؐ/hN����<ummm���	q�����)������<Z�	$Fy�����Hf^	��� �)����*�H��brr�;��y�ז6�c��+_7f����{>�M��WU�'y�3k��M�Y�����M`h'W�V�ч�iD<�%Y���u����<n��zK�� ����%)9(v��I���I���iI�W_}ULMM�C�Ir�0Р��=*I���?�����~�Ԁ��:uJ���I���ڵk�kc�dffV�����h}��2����Էy����~p�Ơ	o�~�7Es3:�#��)��]{��A�.lo�b2f �B�o �q������k��s�l���� �<~���?;;+?�<yRj���qI8&�ŋ%A����$r���k�|����|x��Ǡ9���d;p>��`���(<(I�5r�phZd���Ƌ�-��L����Q�>�I�ӽ�*�~�6"�Ƃ'm;HC`����s߽�;���d0�MT�.��s0Ya'_m�_N��4���ʊ�3��fm��ׯ_�ǡ�`1�M��0��6�AHhI�� #��1�	�r6k��Al�9��H *��	r��l��#����D4������nL�������~�ˌ�(v1�Y����$p[�=�0�����������;���9�3�i�4��3߈�����R��		��;&}�b1/t:-"GG�
y҈Y�7��q���k�� ����I��0�O�>-���� '������ a:���H�?��cN�Ք�3��6���Ȯ�rKBF< �憓��oٽW�J�ĵ��ujw׮��Y'�E��=��8~���</��b_��و�������(JGv����dMO����)$"LT�� �1��F�׀��%��И�QY����z��ny.�&�Ľ�l h*��kS��(4����E} �իW�g0��-��ۑ6�O,
\V��iV�s�R��A_��8��7��d5�`��E�w�@x��y�X8x@���@p h<��8����d�Z,��H(Н�	�ɜ^#��yF���^�ny���V��`��%�v�/8�1"Ғ5"j^~F0	��9���ui=9rD^|Mԅs��h��Ax�?ŵ���� ;���0���y.�q��}�7�� >�D�08�<0<�#�[7*�]o������n�
�E��3�����h5�f��z�=A�N'*���/�7IB�� �`�sX+(ª$Nf��\.�O�����<���$��T�8������-Aq����A0hLL��?���A�	�X�Ve�������
�  �ڄ�8@��D���x�~�M�e0��I��0��A-���-Zx�V�~�D�Ev�ae6+K�L=S�� M�v�<��cd�V�8�C���{*�� ���<a��d}l��^�rt���>O��3|;��J�m �&�����Ν;'�s}�E�Z�Q7��	��� �
�炼���e��΃��9[��q��3N�@�������d���}�ny/E�
�~~gD��W���Z�.ƞ +��ʨ�"�D*U@C���0N�c��MTk���YvC�C(ǙR����a��6�4�9P:��Z��� ���A���7���	F�%�9Z���ԟ�ɔG$7WC}++J��c{�E��,�����[I�Kn),56΁p�Zb����&�Y�����]���;�^	e�^T�45Y�d$�	s��iw����@���͓�Y�34�L��n��W��8W�E��+�+W.��8�~ �f-|E �cs��B�nQ���˫�-�LDmU��P,�$E?q���G~�,q�wjjR�
�`��R��Y��xW���L&+���0�;��]��Eن�rږ�<ht��ϱ�������@x��5U_��:��8C?f�L<e��i�ۻp`�y<�����i��f�N�d��B8����1�a�Ü�|�����8�j%K�w�}�<�����n��0?Q��`�3��e 
߃\HAv�`�u��ozӛd���?/^z�U�{Y�r�-2@�~�9sF��������\/ȍ�m����</���ؽ���k�,�����C��[�'��G��S��Udu}s#��.�@R�; DׇLO�0)e�@�O��J�D(9�" 	��a�"�����H���uI4�P>����S-�E� �ܾḖ8��4%F�w��.^�,�0 _��o����~�����]ה}�u��)�>� �����mQ�u�� *���+���W�|?�y\�MCe2��mӮ�]�=AV�1�l�	-�h0���,+�&?>�����Í �i��&���K�Xq.�� ��d�P�H��|�����)h?^���p� |G��r �	
rr�G��}1]�+w؜�9Ե��LA��I��	�6�of-��d�� ��vz��A�#�A'`P����-��]����^�{��d���BP�����T`��͡�@/�8���_��ƐZ7�3��:���EA<�$E����>��L
��E��#aB"�f'4�>�<�#�mٯL�7F�0\����t
_'+��Ǡ��Xdn��a�<�����P}���c����+���M�8J�3�b�Q7e3��UDX��D��!�Bղ�z[�aG��]���^2�1�+�~x~�� rz�t96����[j�3L]ԉ)�~��7�M
���Mh)ݝx��
��qp�L��,ɆB�,�/��nT���g��Pӻ:*��t~QZh
|e�-݉��Ԯ��׈����x%NzK�����*��)3X��w�����]-ϻ���Zg��lg�(12d+�����d�����Q\^:���ג;���r���D�������%���YU& �o��"_,�l>'
%ծ�آS'��{���bq�*	dKjܬ��D�reT��nlJ�\(�P�uYuJ�q�U���g榻��M~�0Tڞ�G�4�>LI��IND�Q�x�@�/��x!�su<�[!�j����������j/<ґ�Ƶ�l$��7����z��=�])/op��j�IûK�gfa��g��D��yV5�tMX��v� �²6�s#����v�;k^����" ���$�Z
�y�n�ŋ5�4�j�V�/h3���N�5�YADJ���9Q���2h��Ye�z}9ǜ ��T�â]����ؾ�9Y}�;��{ԏ� �:��I:��a;ݻt���\kz
HZ;B4�.Ǯ'+��Mq���K�4�&Z�y5<G	!g��f$�����r�	�sʔ��v_?8��M_$ó	�� �D���o �Z���r{��]3�}�i���׺i�2X���n�w�
(T.��w��ڊ�v�h���JD��i��A�~�|�5b�A��3��-��	&�"���}v��-}�H췲=�:�0H��+�9�m��OT�st0�4�-n�.��v娱e�:�� O�p�����4���w�����$�3�80����+��yC4�ۉ��Ќ*B�0p �]�|����Z��Q^����kL~�{�=�Y��ڝH��5N~�z����ǎ��Q6��d�v���S9 �i�:����\��֨��LV�3�M�:^��s<0NW�>H(�S5L$&�J�S}T�Q�ZX˦�AfS�]y�����]>��\f���^���GzkQ>?�]i���1xӃ�����1/�]�=A����������1��̗���mj�@h!DKy*���E
\���Kd��[��r�M����r�,�NbT��4��q�,���d��3^Bǂ��I0M&d:������6K���1 ����G�s��p���ms�_�w, ��!װR�X8n ����nq�;���`���$Ħ%2��̇�Na��d�6:��v�T�B,OK��Px�0k��޸0��b���z�!�LB��I��J����Q��]A�QL��?qB\ev�D
[=$�6m9_��:�J��=��TkIl���o�)�zd�I�KZT��Q�=��d,��'DA�7�|ꓧ���tr�� L��R9��u0�9�(�,�ہ��w,$�)�4�>O>N��U!I+�Kq�'3��Iv��B���)�j���πM�1��l��ֵ�:�c�E?t�Hf:�#��FQ]�r��b���8�P��K����	-�.y��I�t�	�D@�4o�|�8����<��Aط'/kN�HgH!���Iaθ)-v�n>?�>Wͥf�DT���SL=͊���d�<�H��Dߊ!<U]m �<8���K��Lsr�.V��FϤ�����N�������9A��G��E��|�A���)Ұ ����mGI�s�^o�5m����ܣ2]���Yٝ�Im���C�y@�Li'G���D�y����"M�)��A+�t�81]��b�6Ax@���
�r�|e:k(J�Xe1�vgP&&gŒ̊,�S���+�d.�P��6�=`Mu}hE���nHM-BiQ�Z7"y���D���8�@+ps���沩_��#\����u�i�Ao6�6k*�ˤ}f\ �
�a?����i^��*�Noڇ7T�ɬCH�!)��Щz�k�t�	���v��ރ���	&������/M�.�Y9 ��>Ū��=_P=�ݹ�=��KcL��)MH�� Qɤ�����2LiG�{�$D��<�6���ck'�G�����O~�>�ή��]��iA�Պ,J/�T�@����Pn��ox+&�zJ�������F�X�������Q�0�ZX�&k;�� 
dDJ����2���h��WK%�e%8��^�A���i��I�U(��:LZ#�.��X�`&�4H_[jT�4�
h�`���Uf�5���Ҵ6��d���U֑P�R��q(�o^2{I�l��W֤�=��
�Zb�T�+�4ˑ"6.oo��'�;�������"��������yE�Fxȓ|ؑ�4-4#�@A'P��Hm�e'y���З� C�P]-�5{�d$�c� �`F� ?Y.�N�pDkma�f��?N{���<�>t�'�I���<U�2��k���`�WJ��L#a39.�=+�������Gծ���t���m&.�9��t�E��h�'-|� �d]1R(�l.#+#�BqD7dQ�f�	���w����~�����C9Ҭi��:bskC�-�rhD�#"��Xr:R&��h^)���]���N��U[T7�d@�$p�I�/P�q�G�$�.	YN0���W״;��ڰ�<�҈�B.	�bff����Ϝ��'�h���Z�N�t��Sh#T���{��J��)��yi'�9F�r�]iq R�tCX���`�JRQ�"�#5'�i�l˅��>o=#�J�R���g�"�*��,��t��l[�tf z���<�͑���:�;yT�C�����?z���[bcO��+$���n9��'�v�҅���Έ���f��}��g>y�d��hOEo�F}��� ���bjrF���߼r��;/�#�7�<�ǰ���3w=��3�͚�4���M��M�TF����8q����ٙ�e:��{��T��f�����זE��#墜j4��V���v���<p�T	�d'�A:����b{{SjdN����hn����-Р5�\(��q�_%rtol�_��9����]3��T��*�����ЀSI��H���b}}��j���fĂu����)u��a�iH[�,�M���b,�C�"�Ly�JD����-�z}ll|��	����a1�i?v���y���.Ǟ +��Vz{����<�!��ٯ|e��K~�@fW�\�$@j�/�ɴo����?��pϛ���("�]��	�X�m��H�n��Ux,?�&����#q~a���O��Gzf|�y�
,�u�F���82z�ԫ�s���q�����ێv7�浳(?R*W?��>�3do�Z�7��;f�-$Է�����z��c0�� 1
���#�����>G}��"�]Ǭe����[���oOP=�߼"�s��?~��h�Z��%��}���Å\΅���O�~�g�u�j'��ٙ�{���ӓs_#3{>�Yӈ�t�Nfcs��'�|�69@�Qj�f��}��c�~�#���~�Vk:�0�Z��P��������3dM�|��
��3���s�/��P�RɎ�92�Y��J�W[�6�i���S��[Z:��w�������xe�4LK
�FԱ�YC�>56���C�e�Pf�Y���[��[�r��&��ӕ��Ȓ����:�f�Ri�k��~�Sk�56�cD�����e�� ��\��RcU����Ha�\�vtδ���N�{7�q_.�-NOO�9�.�A���FGGD�2.5(}�3���b�J�8���������S�<G���U{W����T�z���yjj�97g?��g��{������O������Ct�������Ĥ���U�7V��mb�bO�u�B)�7;�`��!�H�hV7���l��Z����p_��a�ۑ�w���
	m�4|0�@V����XY�淶7��Ϥ�B�y�����s&�Ƅ�l"גB�"җ��瑏|���Rue����;��*��&��������n�s%q�[�&C���f,���ʅ2Q<������7V�����B>S*ܙ�)iF��9��9��qԳ}��g�Z�d��q6�	<�la�ݩ�GD��#rkS���Q2ţv����]��f�Y��,����19XFXL��B!;v��#=71��U�Vȧ��yQ��r���&�������߲��(d��"���3����.���k��~9@��.������?��o�n���s�d��W�<�JV �L]�~�]T���c2�_��� �^�-B��L��d���7?p��s��<�ܢ���ڲ�V�j6��TW�o�4\�&��5�Qq�H|³��o\��|�t��;F�`Đ�4����*q��J���l�Jd��VY�|>b3UF�#[=Ԃ������L6S���N���ܿ�pM�l��V�q�������m��j;��|�;{�,xsT�ah�
L�k�bii��9W"mbن�N�.�
0�4+
q.��/�ฎ��t��LÖ�AK"�-[(o����Qp2�i,�C6��hLޱLioֶ�4Re|��v��	aX�����k;x���h�ՂhS��~�/-/㺖��Fh>��}�l�F���u
j�kK-���xKLo='��ۙ�.��xTu,w>a�4p� -o%���\��Aal��<e��j;�4��ғO~a*h��ll��[�r9��M9���x��ɲ���F
#����Jx�[~�WƧ�N/^��3�O;�5C�i��H���`jf���DvЌ��������Dquu���ȄK��.׬�[bjҹ�a��ێ�B�0���D��x$��9���&*Q�>��,13=�h�����7o�A�2�zy(3:Z�kY���v��a$�X[��ێ�v����X3�ѨuZ�a9*�vɄ6e_Q�:ᇶe���t�����4��6���m��e�(���o6[��Mo*W(��`�m���]��n&'�����&KŲ����vB�yI^mku�s��\q����djj�ޞ$S�qܼñ�c^������[I#M4�;�OMM���aL�0�����Z�>Z.�~�ṭaǻ��]s��Fl���.G>?�0�����Ri�c�ߚ����FFˣH(h����X���+�H�5H��3�����-0E�00��#_ɒ���{ʛ���d��s�i��v��>k~;(w�~�,�mը��kQY'+�����/z��n�f�&K!b'���(�t��0%J�R��b>���ho�5�h�y^P�sǦ������{~�L�:��g��.v����U��fw�z�4��<~�퉨�͠ɚ����(�wj���V�_�z}�����å�|>{�fes�ً��Ƨ\#\$3�dF?z��R819sajz�k�Q���j��ŋ�Eat�<R�����D�tǩ���7B�*���F7�0�b"�oц�u*[[�4�3Y7ɟ��Ds��9K��f3����7�_�2�C����jed�F�U*��͍��zckӲ�e(.��X��VZ�~ߏ������e��ֺ�j�CL�LL�I�nnn#�ա��JVƷ
��w�|�[|ݝN�E�'��\����Gq`(h֬랣������o�=M֛�X��_�ӭ�T׷�9�����������a� r��ŕ���m�\�xT���V�s�]�8�R���Nyr�r���y���.z5o��7��d� Ђ̥�+K���K�h�2�)�-ô}����_ϛ��`*h5� ��F9�BĎ/���J��(��#�}�O�����?&_�ݵ�9�j7�Hs�alT�������d��i_%�/F���{��#]͖����i���'� �Z�V@}��M"��/�V�+���}g����'��?�����j��o`�Q�-6���@E~>iT����.44Yo�D�>q��˫�!���x�D"�fDeLM�	�����N[��+++� ��^k��6�?g��wg��ļm���R�@�#��4HC���"�c���|����?���+���|q���T.$�����8�u:y۱�D�e�u^���Kq���C�H�o���~��~�ٯ��Q2���F���Y��u.ۙ��x�靮����u���/��CԽ2W�YChf��e7��z������|��-�����/?�iw
CLU�U�v�z��\���s����q�C�	M���o��s����i��}G������������9��F�����\x��`�"c��ߌ"�
B��a>��Q��o!�CZ��k˵�{��jR��G�`q��+�i<H�_�X*�'[sMk�ĉn����Ï�Fox�v�}9d�_{�>���~����ٳ���-��Ltdem���'������}\y���Z���4�8v�z��?;���I֙FM���0�;� �"�,�>ݷn�}?e�#7�g(������/Iڅ潚���X8|������xCh�ވ����CMV�!�&��Ɛ@�UCcH�ɪ�1$�d��h�jh	4Y54���CMV�!�&��Ɛ@�UCcH�ɪ�1$�d��h�jh	4Y54���CMV�!�&��Ɛ@�UCcH�ɪ�1$�d��h�jh	4Y54���CMV�!�&��Ɛ@�UCcH�ɪ�1$�d��h�jh	4Y54���CMV�!�&��Ɛ@�UCcH�ɪ�1$���)l|�>�    IEND�B`�PK
     w�O\���|  |  /   images/6fad6c1f-1fec-41b3-8a64-12aeedea4fac.png�PNG

   IHDR   d   3   ai�   	pHYs  �  ��+  .IDATx��Zkl�u>w��&�K."EI�D�a[��M*A�+n��U�m�i4�]vRM��O���(I۸E�v[��h�8m$[�+?��e[�%��{Iqw��׼��ܙ���k�!V����ٙ;w�w�w�sg%hZCY��& fM@̚�4�5i0k�`����	H�ن �y8�	�D`�����
�����sO��w��k�G��r�V���h`[��S��O7,0�g�Z Ӊ�9�YQ�0����.(�@�\�Oq�2���,�r�׻\<��9"����$�����cCU7aύ���8d2[C�Նe�$�|��H_�ԭ���_�x:;T��b��{K���;mnn�s��L� �n�je$f��E!�P�ܲ 3#?����q��V�!�a�e3N:���*8���.�����x�����]�4`1�PUD�ښ��W@A��j:�`��LM�6�Oa���G���<�ԓ�����ҙ�|���jֱ�ݽ������՚5����X<�Y6�m�J&Sӝ��m�5U�~����"�"+J2�<u~���!@�{1̏2pʱ8SMN�q2o�T-�Ǟ#m"@0CAҾ�/��N�K+�ku��� S�D2�5Ƕ/#�;��gd#GVM����ڿ����s��i����`�����P�* Ǐ�s��#0>6&�w���eת}U��M��Ԭ'9*���UW?Q%�N	#�}}��hIgscc��"
��,y����w^���]��W
��w!��Pf��K�U���I�}��S��;��,��aS��X�����"8iI �t��Þ�������m�?�����p��~�eܺ�}�o�S�O��� q�3>� lT�������ш*�cQ-�i�1(W�L���_��Q%�i�(2���R�op<��y�,�vE8a9Bjr�َ����#��5 �N5G����YSd֏3	��a�_��~Yc�"�п�pk��"�'��W�����9x�(��W���m{ަ��K�����OO� ����E[���<��P�y~a�Rq�#���l\�8��Q�AD��,@�
���
���������ש����@��~Z����x�`�ex��3x]}�6O*������E-����|��
]�Ͽ��7�ǯ��[h�0TT�>�(<����}r� �|+���#��<�����c�=�5B��UE,Q m}u从�͂O��� �Af|,~.WY��L���_��S�{C 4$7F��m�ha�
�B/�"eIV��D��߱|'y��#�;��U��'��ȩ�ߵf�ˁ#�����<��Y���+�]���<
?� ���������ʮcGHV�e�r��E8v�.(
SD}?��.w:�X�s����>X �2���H$��lB"���bR�?f���2�Jb-�*8H�V�NV��8,//s�軵��
?��T�9�I��� 1�9�'���3�����s]�$�o��	w�c�Â�D����;���i?��`ee��As{���~XZZ
2 `ff��26��@:��.\���&c[k�����k�8-qݜ�o�;������qe��ݰm` �}�Y�\�xuN�|���:�{k����e�řA2�,0��E���"fI�T�h4��H������(��g,�\\D"��G*̿����DW4��i�2�gt]X ��D	�lG����0�{o��&'�29�NQ������A����tN�Z����ܲ9 }}}0==�#^UU<nq� �%�(k�J���":#�"��8�K�t�÷\�]�T�7�l���L���a�-<@(�("ED�rZ	邢�E��#��T��#R���.��u���!�ñx�����*,.^����x��}��5�@+�֜NߗJe~.����]�	��n�@�Ѿ��������5������:��pR�P���ԋ;E�i�~F8><b����Y��t:���|<*����0<<�/_�ل�-@*�:8�H�q���H$
��i������m���cM�-��)u��>=���H�}u֋���B��E*:�bY&�������NԲ^�
��/��u���8-..u��7�����v$�#��i����u����(����U��i
{*E4�� 1��烞#P��q2.��L�qj�d�b,���¬!:o��$Z,����������s�ܚe)�G�b��!���/̃���w���=Fk#��B(PUQ�'��Z�KX�Ɇ��X1p�*�X<��#
M�g��(>.��|FB "�����aP9�q֐X�t�
`�7Z���� �U���d�1_�ō��@M��u�~�p@/�P�L�+��������0d�b\ܷl)�������ZL��4�V��u��㶍��u�~~�҉Z�P}�E<zVzx���ܜ�o�k���Br�])�>r���#�,�&��X���l�w�o��6}�U��r��|w��$, ���$��^�̨�� z�-4@&''��CYMU$�9����*�`��	�JHV2!�K�_hj��pt���2�o� ]z�l��>�fϦS|�
H�9�����*��x,X�r8͹A1>._��[{���cc(I/�([E�є �`X~�j��N�7_N�w�,��nЋԕ_��&M!h�d�o��(�%��B�㵅V}�� ��-Z��� �k�}F�v�:�]�)�:FZ4hϴEl۔U5�%��FN&5���حw�ݵk�3[���P����SN9P��W��xmy)��^RF��:"ј���_���|d.7+*�{���v3��E�,����E�;:�֖V�{yvvV0M�g�����(
�mr�9�kЫ �E}}���B�Z���V_��Zg�<^�F"Jg&}nӦ�B�\	�m�B�S��С_�8y��z��גo��7]|���ӭ�XR��m�����{������{�qU���EQy�#w�Ƨm�3��ū211�@4�q.��?ڹ���c��ML^9r���.�(M�|+��x)��!6�w.,�lJ��^,��{Q�j�}�ӓ��X\�Y�3�����TK:�E�ό\�x�K�	AI���W�Vġ���/�}�t���� ��۹J���_��o��r�Z���}3���46��J�L�;��;Uܲ�WH�P��ȃU����=8�/�<S���~iǶ~�=�iOw0�n�X3��d��#�6p�ayie�����Hz�Ρ)��=��r</#A����m*�#E����Y�f�^��)$���;�B%5e\'y����o~��w/\��.��p?<����o����c��3/�;���D���d\�DD��H;n1�h�ѱO$�lww��2�#�&��Ȳ>����=��i�:��ֶ��R��uC7bF{-�Ut�x$��R�}�u�^U�1ch]�U��<����%YT#��_J�J+˫}�فeFR4^�mvL~��?�>xn���y�<���|�a?�nݵL�TZ�������}�?��MU7vd���j�2Fbqtρ#�f'����ɩ���3��cֶ����UM�����Q��e�K�8V��M�F�cgɦ���+���˺�R�~HU4ӱݟ��z1M�P(.}@��^EUZ������9$�x���մ��J�=��c?�����t�J6�6��o��Ih���#��~ֲ�&�L��[���8�����Ӣ���9	�i]7avv��-[z�mk�t���*v˭X�s-����DT�VK7�˥~L�K�g���6�\��ʁC��cEAT�`TJ$�Y����:�jk������v;9�tk:~�k;�EQ�(	�O˥U����m��6���]]�Q�L���
H��@�eZ�"�i&,�k�H�6*�ר�҂#���MݨX�g��藌$y1�*5���П�EJRK�:,*Þ}�r�:|F=���W�?y~���9�r9��\�v���f��a��8ϑ��zEj�z�n>�!>����f�����=��u{�G��u��{�Q�������ɮ;@~٭	H�Y��& fM@̚�4�5i0k�`����	H�Y��& fM@����?��3    IEND�B`�PK
     w�O\tX�K�~  �~  /   images/80e9010a-c477-4737-bb01-43c9d75c1ab5.png�PNG

   IHDR   �   ^   F�=   gAMA  ���a   	pHYs  �  ��o�d  ~tIDATx���g�e�q&����\��m��@7@�4<@��N�+�(R!E(VcV��U�L�/�[E�Ɔv��YI�#�(G�\
� �0������������޻�}yΫg��>V?w�9y2���2Ox��{�l6+����Zn;pP��%��R��$��H�$R�V%�NK&c�[����a�(���� �TJ���M�~,8q��'�n����>���8&�K�R|]o�%��㸍z]R�7�����ZM���%�7�M����K"�]���I���>�5.--�����|]���8��J��k)
|���K�_oܸ��-..Jww�K�\��7oʦM�$���������~.^�(۶m���>=_MjzM�������e����뱱1)�<�׀�SSS�����y�[�nɆx/����^>�X�1�s�����'����1_8��s�\sssK\����9N;w��N�p�t��q�3�S*#5Y�v��� �.]��k�V��q���5k��իW������s�덪��ϒ$�k*���؄�0#��'99��e���h�q�T*��B�$7��P��0��&��t:��Ӊ�sd�i=�	m���k�&�m��	$7��x-��Wu�����:�e����^N���lg����yٲe����:�8��u�)�7n��@�0`
΃A�w1�^� (<|aƄ���i����k)��<~�8?�������;��-ȉ�'9qqҦ�9s����o  kc���a�0�x�}|��*��������>�~������JZ�����q+��׉1�B���1ſ1�S��%]48�iA﹥׶y�F^'��z@vn�)%=�ٳ�U@ǹ���0FXą\A�;G[;�1�~���v�^��
7�lY2fubk*�U�ҕ֨�)`�LZo0�n�5$�����xzM�A�`HJcX�f���M��&ܸ���Y�)\Mx/�v��� �q�ٯ���((8����5!����}a� ��^x�k�|�2�n޼�B̓�B0!��d����߅�Cxql��Ƹ�gϞ�k\kiڰ��
E�T˂������Ƹ@��z1�/L�>��kL*�����a��x��1ЎР��ѱ5|׋����aL���ap,��A��ĉ���j*+g�&jK)3G��E�s~��E'Ux��ǌ�1$������G��0��0�P"�����EF�H���i6q`\H;jQ�pѫ�B�V�	��Z�WO�	I‫𠧧���j����4������O}T�cWt�h�1��^ׄ�������?�&r+o���}�v�^���:�/L"��:q��.׊�1����I��lݺ���kn����}��'9����<����#��[o���ٴq'��뱵c:a^�HQ�����]����u��w�]w���a���^������&�k�7���u��ɕ+W���A����3������:�7��رc��n����������Op�]8^�I�͇{nS��oQ[z_��1���Z�0�K���:��j̡��*���W磪���-�(�I�)��T;[B{���D���k=/�^0�7��߸�t��9�7j:@�=?�x�����c�p��3�T&�rC���ٙYy��祦B^���ٛ&*4�i\qOW�����`�qh(���`B(0i�?`&���m	��s��	
��ñ����������x}���a&��5��/�x-/��SB`=�����~q=8΁��5@�p�8.c��q�����b����g�-�y��?�c����q�WA��?�C[��W���uY\X��lQؗ�$����`�Z�0m�N�/��Ó�V1����J���ʁ^K�Vq�ec0?���WB�(Fw�G��oM�#ͥ�^kz�����Rm0l�S�_���`
TRzI���<�С.
Lh#
/ի�����X��S�u�'9Л����/��NJ���c�S�N��������{����;Բx��{�h���LA� @`��;ta�0t��as,�|.߁Xx�a���AZ��J�Z"Y\Z��c�ba�;w�׃cB�<�V���!������V����q��v:|:x?�u�|}�ȑ|��0��*��I#L��l�ܖ�uOO/%L{Z����y�1�Q��P	�&�ʑ�{��[�^5, ���0���f����$�k�������ja�'�T�{w�j�y�LHB�d�8К������>I��xm^Sc�b01	<�LN�*�xL0�DL�0I^�y�I�w�ˈ�Ĥz'��?f�ip� �1���p��z�P���m���ڱ^U���M�S/l�K|f5�Ɇ։�ilA��Jaq��#�����"�( .^{���{������ƿ�stxD�y��T�U��VB��&IR��pQ꽤�I�
&�~���s҉�������RaB9�1yC�LV��o��˕O��OЊ��;�������������eU�Sت�8�?���.��;��*Ɋ&� P��Z�B���㺲��Cp<N�;M�CUд��������X��
�dU�ʏ���^me�-6h�T���:LS��}���j�Y
X�0cV��NE��;	�^�pf�9^���9v�Fl�80p���� ����)N�z'������$���]ja�ʀz֥JY_C�b�e�Ջ��e�#�Yǜ:��;�}'���{P(�HN�˥頜?w�_m�;�9��p�����q��J\3e� X�@��U��HƄ���;�L�3 +)1g�A�;g�V��O��#��P�A�}��=�e����:$��s�@\����#�v�ZL.^���AXq�p���@�r��t�a�Pz�Z��a5/x��g������iL{@�8iomh2�"��ڂJ��u�T8�Q�E	�g��9���j��iX�a�1k���"�KC
�_��0��s�eP5����a�T���:�(��R�%\T�^����8�H�'�R�Y�Eӿ��P�b�y�]�H�hVCz�	�8�Ϙ]�����xͤԯ��]�5$�Įt���~Ef����n�3p}��<��Q��<\��sEH�F[�1��|������|C�?������&��:<�͛g/�ʃ�C=$����O��뇠zm�zѮTj�T¸&&ZТ	�"4~���㚲����C�j5ۄЦa�4q[�h���s^��ՂI��q��[{��hI1i��qdh�T`c�s�ڵ������u7����+�Ϝ�7�|K^��11S.��TSŘ &�<){'p��%�S17%��cu�B.%�.�\5:P��M���|¤f8R������0�ߌ�����U��� -W�3	�5#���T�����`L���غ�Zf2�<P�֤I�8(�����������+������_.NLH����j
�|���-���j�*�8&	Y8>8�q��yy�����A��3��sV���|��	/�G�`��7���u-!~
�7�Nϵk�ezz���B!GMZ)�)p�i�y��NB�H`<6$N[���+��!�G���Z�!l��3�p� Ͷm�!gΞ��j��֭���Q�����z��/H�?du�tw��R*S)q��6��5p�.MK)�C�:taAv�	�yY����.�B��ڀ�Ftd2z��;7,R �Ϡ�0#���I[���^<�$S����vd)�o}�[4S�S21q���I�tFG{���-�
o�+m&#�9UC�-���93�E�Oࢂ�j|��=z�� � �f�s���}]��>�-�1�h�$�iAf������_��1���~;q����qS& ���H	����x◾����	��,��_]~��1b`���NijP�]�������ă�8�~��W��x$,t�1����{��z��-z]����<y�|��rJ�޸~M��=R���:���*��TZu^_^a,�h���N��Kxm� a&1��ċJ���7IOF�G�ʂ�����%��~Y�����Y3<(5�K�*4%<�
^�FB�`��]e�F`ʢV�'��2̑�b0��]ҭ�X%1��\Vi�h{o�@?O�+�'��k���,<{t���;�q*�AH����w�l�2NS����چF�T�m�;�W!�{��?�S9u��a��ڟ�b|F@�c�J��q�Y;$����/�+224ܱ���V-��c�=&���@�t��i�e�1�N���P'����~xO��쐃Z>��1;u�S�q��CR�֘�|��W1#���)��f�:�t�)�<��Ԋv��8
[b]`��k�g~A�k��T���9Xm�~��GdxxT�e�V�lo^�J��!�]&���E�M�KH<��ĥ+�t�_���e�_jJ�aN�#�o1%	����U��M�l�,k� � ǋ,ʾ}��|~�1�7V�NOX����Hm%���&��B霓Ց�ؑ9B�Ҍ������=��^�zM�֚N.B��c��G}�i��ÙȪ!���'�� ���D1�[��UgbTq�N�;d��]*��ԫ\�
�{A~����K_��\ֱ� Y�pb��[�W�c�Z�&�p��1bs1]�ǆ�b��Gz��ea�$g��eT(뵆^�Z4X:���z�z�����z�v��y*v�ՋW�M�P2��Ӧ6�h������nu��3�l푭;6K�� QL5��� C����&��:�EܻK##g�_��{E�{��ܸ� ��.��t�Yg�+ԕ3<�V���8��kx�&D�Çӄ��'?�Ǐ�ʯ3]	�Zq&�V���b"3 E�_�Bz��d��(����CJ,(&i��ҜNdT�����V�ɩ�*����p�A<ّ���C�����e�Q1�>���q��ʇ�T��6>x� �,���[4����?׭]��M-F�����&��٨7i&� ٹ���W�g"������e}����r���'�xJ�~�����]F׬��^{M墪�<���i��aƁ̣2�=��t˚�~��/���(tWW7�n]����"/XDs�s�a�6���$�8sTvl�tT�L�':�p\2�0�j�R�z��j��ݳu�DOVX�%o���j�Y]6 Y��F�p�]�qS�?)�
�w���m�^�l�rꔾ������6���8��C@��H�U��߁��s���T��`��ڵk��L�;ϐV!O7���o׬���V��g��XGW�,//R�`�֌��pZ	�&~tt�Z�s�	��r8,m�}� a���E�y�
&���ŋ��b��>�q�����DX���+��c:q��hS#H��Z���ϊ�/z���.�)�AB��_��<�'娚�w��@��N�����������#y��?�����W�3���P���\M��6�]w�&��![�mf7_���X���f3Y�0�`�.�9��������s���8PT�pa[%>"C$�I�H���F��J���j*U����ܱo\��&u��ʇr�ⴴR!��(���E}A=�O?�@�CQ���.gNM����LO�2ߋAw�D�<2c�p\'��䟨�EP�������\�Єx>�����(g�]0<�ւvv3���F�)Gh8BW�l�JK���"#J5'��.(F!����R�qL`O�.��
�
��BM5KY�sP���v}�:��3\5(���4Or-��b� C��q�87�j����F��:Ș5w��7�X0����㽈ĸ,�w�u�L\�İ���IyG5����䵷ޑM���F�� eqڂ�J��ĝ{7��~R�T���A�#�,*Wp���><0l��H�p�Ȁ|J��ܚ>z���^��Ё=��g$Q�*&�1�1Ob9��b��HM�� <��TP��
h����6FZڥ���ڭEI��X���j����.�L1��]~b�oI�[V�Q^,q��� ����_�"�Z5+�xL)���z��}>TO�K��K_��N�:����\ �������h�!�]C�Y���q2Cŗ�z�iٿ��lڸI*"Ckz��	������B+te�Cq���z�l!o����\I-��t'BP��22)*�0s}�]��Q%�ٶe�s�
64%L>4\��4!��3����Sjoj�E�ZLA�#X
X8���nP�< ��\�x�5xNz�K�}@nA^������Kmq���ݷo�_��r���2<�[I]�Vf�"�{sYB�vC��Q�N-��� ���-�y�W�t�d�E�Eu�z	h!���-�/[�[�R��2?�3(w��.o�{\Au %U�5�(����
ڣ�8r���깕�-kG��΃IH-�k��aE��c����@H�Mn)N��Ay����ٳtT�>Π�E��I 8�u��f�±q�z33*@ ��45���S�R��׮0`�v��7����Ag �.���Q�d�#G�J^�Ɇ�����¤�;N���4�v�����y]tRBh�˗dnfF�oMqQ���n�[4�igex:�F�nv25����&|�ç�tO\&�o��Pft����Ȯ�������
M�ÿ�O�k��R�Sx�.��BF���'�������(T\�vi�x����d��Vu�´+�zܔꀧU��U�m�$���$C�qF��JF� �yh`<�L��t��f��!��
]^Oڮ�JjF���HoOQWQ�\[h���Pm �E�{����ߔ�������<��o˿��J�=.����j����G;6u�N�!Z280��z�bT��������w�ȱ�1��Er<���ɹ���KD�O�x�5��)��8�P�s����	M��n���L�19���(���������������Z/v�@?~^��/��]u�ngVu��Z(�@�)�bƧO�$�Ţ�~��VЮ�"����Lڒz�������,d���IS�T���B�Ȃlă�ߘ������/��|��~U.\R�������l��:B��,ʲ���| ;���o|�II�Ӓj-��̪��
QF"��0R�.��9U�9]��Ttѕ-YU�I�&wZFՓT��J2R/̼aĜ�F����1�ȗ���d%�Qi �կ+|�� .�JT샌�
��];Up�'�����E�d�d��Mx�_������O��ʥ2M"��\�@<��TV�.�bh�i��oc�\��62$K��"�o�&ˊ-G׌���c�}�n< 0(� ����QG鲜9s�1S�N%4%L��i�P@��{�]�L��A�/� ��y/_�H�8眞�R�8 ��U�o���EXVa�:��Ӝ:v� �9�A�V��&R��v+�<��?#�A�Ǣ���E&����O�BhqMW�^��S�{�>�S�Я�˧ǎ�O���Lޔ����RSe3��x���{�گ�EX�,�P�4E�LJ1��򄈈"+������C>(o8��c���ڻk�t�Ҭ,��Y("���������J �M�8������=UU7jM5�'dd���4#H�F�������埾$j
>=rT6�����5A��e
�	p�ي냐���Ȧ�� ���׾�52������u���%a�%��\RhahQdd��:��?x��	k��a$�@�쏥�쏭�s�c�V��W�!�r��M*�Ctl�{�G���鑟=J֬]���'��O���vR��>�Lmi�&B���L�bӿ�I���\�J(b�W�A ���c�!������N�'�B� �����Ó��7�0t�����������I�.��B,��K�e|�v�W�����p.��[����̸B��^�vO�CF�a�&Ͷ��HR�U�مH��7��$nX�Fz�y�wT�t���H�U)�� *ΪM[L�����6J+R=��UUOޘw$����f��ȥ�la��&u^f���G�tlP�`���)z�8�c�ؙj5�w��{z�;�Y)ds�]�Vx�a����}Ҍ(`�<���okB`����3ȯ���Fp^j��2����;��1���S�jN�|h�[S7)�C��z�Y�����߾m;�����d}��k�
�q{0q@Ү[�i�p�!�ޯ�	Ҹ�l�e���������0,�{âL�	G}5a|u��3��~I�d�צ��c�����Tf�7wm�*�������2<��ѡ>�UKRo-H1hI)fjp�t�2�H��U�U%󬉴4�B�5�*QM�Ʋ���$hP������Y8uz�ݽ�QJ�)�v��:�z�Z������N����	]Q������(FYn��7��mٿw�����r�bP�$�����KB�瘃c� �b��Ơ!9����w�g�j��=�c���u�,��g�j�u��T�Ef691c��Y
LN&3@G	�5��p ���*R��&Sm��+�e������ ���g��K
��Q��QZZ^�1�"
}�c�ˇ0O�+C^S�qA�@| �AhoO��5\����s57�S =Y�� a:�d�[�e��/��w�Xn�,gO�T-�@���QG�mD}5���du�ӑU,��F�	P�NV5ic_A�� G�:�Y޶:�iu�O�>A�2��ax� bܛ�M��H�|$�JH��V[r���<Z��uEգ@N��('O_P���Z��� B8���?{N�x�1y��Ge�jM�~��0K���o0��\^2
��|�s�U���:��j�O�|*۶o�P���Nb�W_yE�|�5�0�)�X��x�҄��j\<�ʢ}=}��Y��fv+p,)
�.�k�	=X#V�,�(�6rL:4ޢ��'�(\J�jm�����j�~�q��[)�@��^c��=�Y� ��m`4#j'������\�	�|Ӥ	1w�a߾�����c��zf�Y={���w�J��y�1�I��]��.o��ն�J��(�v�QXd�P���q!X۠��`�=���I���u��yN�|3�-y�1�
�8A�DX��8@<�*��V*��T��Vlz�Ƭ���Gr���ԒJ*��@�	�q}��O>�X֭c����)����u�DtP�������#P�햫���2Ŧ���	����ٻv���LM3� G�2@+���#��+���ϡ/���$l�9��t�c@H�x.N(�m�|�";i�j��3�}y�N>	� 幁��qlw�d���,�c�#+�~���"�ijuj*�`\����'��9��/��L�CS����ܳc�lۼETՂ�z�|�Y�X-TeQ�:���/�3גٹ9y�l�4$[F{��Q' N��䜂�G�T�����3�0�%m�i�Q�D����$�7$˪1�ͪ�t!0�@)RO�45$=@"u��ٮ�"�95)o}zQ���,�N^�BN��r �w]�p^q��x��_��GB�z�)y��7ueN�Yj�N\m:Xs3Ӳ�&�	�sV9W"����q�� �hq�) �Ywe����Υc�TO��Q�X�u|�1QVe^�sde-�R�[#_��H�8+�1T8�,J�V
:yp��[#.`hלb����&0I\&(乱8hϳP�AX�g
�[:d�[��)�3���ܻ|�[��	l�l�T��X/�7��K�S�UHw��-�����&��:��o����#�JS�^�.�fd�� Ed�Zv/ı$OE����[Dg)fd0�	 �0;5'�=$U,HV��4R���o�9�A�I���䩶����K%�t㦼��������9�P3����on�ꬤ�w��z�m�e箽���غU�~��23]]�N�/n�	�Qgg�_yh�|�qR� �L�V�`!8���:p��%pD ,מ�pCc�sͦ]^�.�@Xqn~��Є��3i��d�$�)S�Nɇ�<��\�4�o(Q���z"����"��j���ʃV�.���v�[�V>��#��EA�^%l�+����J�޼�P��µ_���V�4�
 ����e���rǁ;x��V�;�.��˯�#�G����RBw�YUz%�ҁ�׮����b�BFM��h���Q�!<scA֎�ҳ�W��+�&��=��M7�V�i�)�mȲ�O`�jc^nܸ&�M��\��e5)F���� �������͍�]w��;�3�Ы�a�T��?�P^z���z�d�޽r���|a��k��iՠx�~��A���*vu�`�������#�8��g�0Uj�C+�Q��F �.���!�0�5i�z��|ӾeN(]�.
f,�t�+B���Ք]��g�57�FsJǤr�z�i��5Y���/V�n*�k����X�q�5>+p�g3C��*��w���Ği�Ha����Ǆ?p��e�q�]�2�U���yR�vzf��14�O��!Cųғ��[7�O2$�$��te�f��j֨Qۉ/1	IB�0�>���&	?8uI6W[�m��?"S7����PWo<��4V�R����,W4#eՆ�5�91��(�6����@b�Bj��>'_��X#���#����r��q$��YN�&�c�<B��̔z��L��OO/�5I!ܱC1��nNKQ��ۘ*��}��'h��%�JƗ+�۫[�D���܏c�%��dWe֚�Yn�&s;I�����&�z&]�L��0�XQhf�zOO���Iס���b0�?�Ym=����%��<�ҹ`hY��|�$��P{{�"��4%4��\W^�j:�o��w�a��Xj��ȥ�������Wn��;�X����ψԄ|t�"+)&g�d|���לt��]��l���ʩ+�>V�*Ά^{$��bu��p���� ��M�Ή�ˉ��<IO1#a�&m����m�5cc������l��Xϡ��Ӵ�6̄N��
L���8��j�3�g�.��Va|��I���^�����{������^�7����ӧ�!TRo�	k=���#h\t��y[���I�Q��Vʞ�C(t�PFm�lF��A>�%�i���{I��v��@�����`FM`yi��(v2�=h{`^0, BNVSou��.�QÒB-���/�9��`Kg������!�O�S�װ&ͦ)8n�\�6��Eu���#�RK��K*�2����zK6o\c��"�Q��"��Y[�Y� ����.]��
�Zr���R�ԁd1�)Q&V��miJH: ����T��R�Ij,��k�"�����=�6���3����K��?�X���e��=��ÏHN�fY�p2A�8y��ص������Л�Ii����h�:`I�b��0�0������'��,ql��_bzo�#��z�k��4x-���h��2lr�e�.m�FN�bt�癢N
"u0�}�-Wb�rǌxK�LstY%:��t�2֬�xUy�+�i���:����
��k�N�R��6�J�*�Tj�瞐yD�ӌ:<�8�ydd $,�HוO�8ꢪ-),,M���s����*�nUJ�)�2��\7�Y��$je(���U.�j�Ŧ��m�yŖ�D����:S�څ ��ʅ6ڕ4���������+�*	,�����ʵk��{����}V���w�~Š�Zoٺ�� #��:�%]-�J���34��"��r��$i�%ߌlܴ����@�]L|�$&��D�k5�)
���$Z�V���#F&�v��X5���LM�z)t��js�W���i�6�-3ݑk�M��c�b��s�L����yy�
���0�S�M��T�B;WIȊ�N�
��Z)�]9���>Uw\�o��ۘ���F���*���(ՀsSo"�X<��2�Z�UZ��e_��c���Q��8�/eT&a���哏O�`F�<L頡�(�� �m$m��!�
�N��
ːj9&Ȏ��&�P������+���-X>�]7t��y�m��s��9}��1��y�id`:q�	�3�qX�n�C�������$`5/--R@\�9�adx���$��H%�$%�da.d_�.z��D�:X�8s��_i��jqZ���w��Ir�R^&�h�(�Ӷ sĿ-
��r`}k��,&�XM;җ�"�
ՎWZMv��A���~�Tۺ>K�vԼ����r�c�o9�v}��9��V��xo�ߘW�/h�a]X�$�K:kI��;_�Ur#Y�l�)v� ���Q��K/��rU=��b�� �q3�����@6,@��C�
ɪx��Դ�eg���K�`�rER�j�l^.��$�^��@E��5r��	���U��fys"�8�82��!��A����3���V�ǎu�-=g��hU�`+� ��2R�
f&�������-�lR��9 �cr2�#Q�
�B�)�i1��gߕ%	�S*/r��R0��O!����N�X�@���0����A�C�%p��N#�@�0�`�QM1K�;<:*gN����h�h�}Wg�TJ�b T�)g\�����k�h0��$�t6a�#��"J��)dk���e��`�!��8"�>�hՓ����A��3����G�UN�$��s�a����M3$�b�;@�ͦ��0�R#@�[a3���T8z����@vH뵬[�گ���c(���<�b���j0��"��5V���o:Mj�YV�.Rc�%j�Tu2�hA���3�M<�$���-��4���:5��N�)lEj�v+�lp<��ФM�@W3[��+ ��Y]���p�VRXc���%ٲe�8<󹂴+fA�>3�8�No�ʡ	7nؠN����(ػu�&;r`�<6��+c���<����M.����wd�"�]R��'@�R]-G�]'>e��H�X�����hJz��9�Zh�%�%Њ�AWyuhS�4ழ\�F!}B�x%�yX�	����q�`����!̔�L���t*����h�Q}�߃�ЭZ!W앚�H��[�Y/_�J����cO<)/<�"���`�Y�*f����*�BG0�m'��@��@�-��`�5�%ap4���!h6\O�4����+��*Ě)�E� g�K��l2�^;�.X��Bv�B�~������
� p>d�г/����3 '��R�>�Eҩ�w�&|��T� �����'?'��7�!'.�Ÿc�e�<�b�di("/�w����Pgs���Ȼ$�]���:�q� ��.f^+����O-�b-ut�#�+	X�{E,(]���=�Ԭ�.��[?�<�8�ږ�z�L��e�����4@����������&ue��3���5ck�_����{�.s"'.]���8z�c��}�.y�'?a#�~���FH(�zZZ�ź^`�=qJ}I�z��,ۅ�Cn�B���@�FN�`�����R����XV. �'�Y��-�|]���^��|�t�t�g~��< �x	@h.�� ��-f~7��t���B^���DlX�!�q.�#���;A0��āă[��#���o����[��G�|"7�nq���<ڰq�������N�:��2��oD��⚱19v���Ţ4�Mk9�B+#�
�n�^���&��MZ�t2\`,IRd�5QXPo�BbJ�j���!;�m'���<˺ �*��5t�@���j>*�{�f�rsM,��A@f����fj�@_߀<��v=v����F��벸�Ĝ1��<~B��-�9{�Մ)�t�zY��:!lBee�i�h`��=u����[����`��t���Z"��3�z�2q4�4<ƬՏô�l�=&&��R�h��4��D��!I����N|1�l�kA|���`ra\�5�����I#��gس��Z-W�;X����V/��^l|\��m�v�3_��<���ĉKe��+�Chε���*�+ЭJ��}�ѱ�w��NF�����211AR&�Ju�bfc��P]j�u���DE��ԭ4q�*���(>���Y���p�p�l^�'w�/}`�� ��� ����~9�\�|fnF�]�&�n���SW���-��"m�ji�b|� ��8�ΜW���1��H�k�v�qF�T7�;�ڱa��6!��ȆMwK��H,�"�w��������U� �Ϻ��=�#RUA_��r�t��d�3��0~�a��7���,\<vDڴ�7���l�I��7��w�eabqY�dgpld����1d2�\x8>�	��։ȫ�����f1dKs��W�, �^i���e�X�|P|�!�r�z>��T���1��/o���.9r��_�KtQem��>�=���QI1/�
 T9uz�*hE5噞���맣��T��ԯh�_�9T+���WE�Z���
��.:)��'P�[��9ST6� �Fd�Շ��o#+,?<zN�������I�Yjr�S"��B���0L���(�_�>�H�G����}�a��ӟg1=8��;)��߶e�|�_�{ݭב�~msN�9'}�������bh�\����P���rU�:q��n(<I���h���dnU�l�S��J�r�n�T�����M�Ym8�H�ɘ0hbZ�߳y�D�X����́�b�ܚ�F�	l��m��	C8����PS\Li�9!��c��X�p�:������gl�"f�0V؏�]?�|����B�U�hb�Q�9ZՆМ���o�� ~��c��^�*�s�hQv�� ;w�˺uc�<$��5����"�泄#�(%��>�? H/ẵC22:�����@��P}lM����6�.��ң+�GMJ��}�S;B[}z��Z�Hw��m:D�aZѰ+d�\�4�t�N�]�����6�wʭ�PM'��r��:	=)���L��=z)Y76"/^W����ifO��Jtv~V�s�D�juI
�9��� qL�S�h���.2�e_ZGč;NJ;2�P a&`g�%Β_13�Õ��I��$�|d ߦ`�&R�q�ɲ�a
.b�k�}`�ٓ�:��o5��\�-��<�أ�'��!����cT붓ү����O ")%��������ߒ9�._��BA!�O�7m���ܺ�U\D���r��y��Cr�=w���[e�%ć��?M���ժ*ڗ^N�.�*��/������_%nԀx&duׄ��B���Ĕfi���PF�������CU��e���d����^�m��"D8?qA�}�V��B�S��vܺy�<����{��ba��˶�?wB��z�Oɹ��֊t�fy=w�uXM/���^�0���t�?��k�b�N��}��}�~� ����Dhq8+�g�S��ߑ݉;N�m�`Պ5�x����!
:�.A�<n-����L��k��j�ڝcY̵I�R`0��V���c�ff�d߾=���t��Yo�_��-;��Ï>B�]3Jo���߄yd.=���B�g\���wr�,�ڹk�:�w�_ҙ�'�9.�l�^מmk���G�[6�f�F��`�@�ś7%ߝ'}���a!��[K�3RY]������Gٿw��m��v�@���y���%�R	OY��|��j�*��a߶{�9}A&g%S�N �<g��D,s���r���dza��&����=y���d-q>����j�am�zm-��,��[�Ҕ�y������	�G :���U� n9��vq"�XvI��Aa�^bd�IL�7�PQ�̬i����YǗ����C��m��Ӷ-�ɓ�i�F!hA8/�j����,����$X���&�)`�!5l�=�g�]a�[0 �$X�*��d-�?�Z�+_��<��Cүp���(�����feq^=���:�3���?�#��W�*_�җ��0��k����
��gn��G.F㮌|���]�7��X�(�\I�T�#扅S �����,9UxmU��W"v��Y����K���Ȇ�!�@7K�z�-kC�T�@?�ܹu��f�-3�Sj�z�dúQul�ɩ�i�R�@ȷ�80�V��o�#3#�?5/��t�Y?��,�|����ʫ2��)RRn�֨�������@f�P��
6��z|��r�>�6YV���j�͎9)�!��TT��<����%�A	���F����e ��-�������/�eU�.r&t]��f8(�RB00q0��N�=�bW��+�=�[$��7�h�qT���0�qn������'�L �|qZƵ-Q\�����3QfK��	h}���g�^����#u�~\W���3�r�jI�?*Mm���+�W.��6��U�n�G9��Q�NPU+\�ၢDjE�YY��'�MVԲ�W�}���tJ+�%}V����[�
�E�a��u-��m-<�<�uڒ�`| Aca�G%��o�$=�'�K\���#�@�2��r5��_�@���!�P >�0�FY����X����:�a�pD��Df�{�XjТ����jL 6E(/V?����~�!B0-����~��N�.�n7x���ۮ��嚿ZH������ �����t ���ˡ[J&�!�x�n��]��1�:;���y"4�X��~˖c��;�A���V�I�a�s�.�6��Λ�@(��K��euLXĨS��k�>����-y��ߗ^x���p��X�\8����E#�;<xp�Z;]��6fc�3�����Q����`(7�m5Ŝ�Ғj�eY�9[Կ��v躄;6o���n�,(� ���n1ͮ���0���Q�9UI�⼨���=/��te���JM���}�qy���>��8�n��C�W��L욐������t������W��g3`�����#4^��i.�F3r�	#�Y��A��*��	�fk;��z���X��:�n��y�.�����B�a�z�:���B��<��-:R���ŵG�V�n�%��\MJɺ����<�XJ(@hL��C�N�*��lE_#n݅�r�e�A�1e� ���f縘п(�c����M��_�u�����C0�`��O�D��y����?��Ȫg�����*#Y�2��yt�����%��&="#>a�K�.���WSA�5ud�a��D�D!Z߰:J���Q�m�<��6kB��8ȫ�����Ҫ�i���(&}��u�6����ky�͗I޻{�:)��	���ڥ�re�q'fe�`�,��z���&�Q(v[a5R����̦)(���.�h�ߕ�"1��hU�����6������$m;m���ۮo���p2��d�La;�	M1��BlKrF�;VE�����B��IL���6ƛ���!��!
 ��z
��EkpҕX�h��f\��eܪ�b�#<cylP�)�7elx�'��`#mɚ.���k7Hߠ�Pԉ�S�HE5�(��#j��1HZ���2Ԯ�"!�-�aŘ�f�r��=����Gx�����d�kL 6��X�M�Ԉ�2h+�@j:8�8�	�l(�.M�&���
�@�ހ:[�=0�~:w�$��}xD^~I����&{�ﴐ���萪�I���	n��ǌRy)Uk2==��E��6�OS��8AF�K�;C�ҭ�6��[��4Ը�ެ�=�	v4����_�M�b����y��3�Ŏ�g�"�&i�4826*MIZ���ɔ��Wo�h�Q�\ �՞�iV8&�r;d�+��&�n?�'�z�&�ƢB��[��!�t �y$`�nޒW_~EnMߒ�����[��^��/����yE���FŉK�ԤUQM.5)�"��%;���p����PH�ѥh����Q_��ޮa�V����z�H��N6p�t A�!����%0�a��h�*��T����:� �d�������1܃��l�I��su��e�fa�_]���r䣷Q�J�fK!j��ޡ^A�Q4�G��2v]ł��iK__�۶�����s�`�C�g��B����p�8V�ө�t
�|�n*0M�V��$r�t�� 1C�^��3�;`�6|�H�K���F�e�w�K:�z�t��N��b�C��c�@�ԱӒhB��x�#�>"���;w3�l��Lyʅ�0{ǎe����.ɒ:�p��~N�DD"6����O$�0��Z�XPGinAF�e��-�F]uIC@!K��brݍXD�lFĞ�B�r\��5�Q3���	gA�Ts��$��kglLb���.�3L�+��-��r$�'.ɉSW��u����R���j23;)W�\���[�W~�Wd�ν�����w��}筷Hk��΃܇���<ZnoS-!�1m�.`è@Ξ��R�厱�#��SԌ#�f�Q&�H��'<�[�E��Ck�c|J�E3)��.�>g-�Q	����'��-�ϦMm{t��7-�`�]�E�9%IGP[.;�8��ϕ[�> 9u����g�+qz����0*���j�_x�~~��V�o��s�[�o�C�	�[���ޠ(q���'�玎|����m����?���ʭ�W$�KdyqA&.\�-�����wS���	l�S
']�����)ϑH��;�e����I�}�[3�_d#(�P4�P��y�`����
I��Œ���%y��2���<Zl� H�j����//O������.0C����GqO�Y���=*@j�e���u�m*�hY�#]ؽB��ͩ�SV�Іj��r���&BQ��+ �`k�ё&�;���za�:�9H0��U�UI�i��>�g�-b&'o�f� h	l����I��N%j+�?%�R�&��BuQ��C��s^�	,�+�q@|=�ļ�Q���إ�0d�m�	z�!��B����@a+�n��܁�j[���/}�kr��òTF��Ů�-]L�[Bt�ƙ3�IuY��߼1+׮�J���]</hGȈ3cm�[��B���e����P$H�Μz��K�H@�&�KU]	�,�-�3N2 �-��2x��R)�s�g���+r���?G�I<E�A�73;/����L���-�?�p �Y������̂�m�"����¥9=u]�m���,��B֩ޖ7n��#������A�'x���\�n�j�x�L(u�Ь+�]���m-eZ5����tj��v���aÇ���:U�^Vpzz��+`/ߗ��K��`�?Ԋَ����xX���֜��m��$4
-��y��w��������@K^�0!���%n�xHoxhD�U���+�Ȥ�)*��k�����mR-ZG� �z��b�ҙ�[��2�\����\��+7�ة�r箍ҝ[#�VIMzݚx��e;�C��� �
3�Y���*���Y�
I��x�:�8p�k��X)�J�A7R���r��M9}sE��b�fp����2��X����C����'�8cK���:б�<}I�Ku��ju��ު��1;�Ā5j��=��k�مC�4����3�h�ZVǩN��Nl�_i���絻���σNvG���]�6m��^#���oe�ؼ+��I|�G���R�a�3�Ng|&�Zn�ٟ{!��74�
��@;�O\�^GL�o��j�}i⢼���o|��O˚�治ݜ������<�����촜WX0�&����jƟ��3����sj����^�9�t}Z>=qNz�r�uݠ�d�0�VT��Zb�j��Q�a]�VY�8�Y��w�Z�^U<'&nJC����E�T=�p��JZ5�OݺEǢ��`fnY�ۢLN�d�Ԧ G�~��vG�O����b������r�K��LGP��������'	30�s�YS*�M:$V��e {,ٞ������Ԕ}nG���U%r!�n��o:B��,疻`<���1+4��
�q�V���RGG�,q��r�y��{�ұ��Q�ʅ��ݶ!��`�4��8�Rm�l!�Hڇ�ڮ��%��� �Kj��9�k�M)\X��\G��,�N<���h	
*/!G��]���T	�YR�����~���&�������l����́#@'�+j��:��?;(C��
g+��<�>{A��2[ȀR���Zv�5��0g��j����FtQf.Exd٤jd[�@�$4���^�4�����x����86<�$@�³��b�/V@�T�fn�EX:�9�fQ��5EȠ��/���pZ]v�ȵ�JK�\����ܘ�-�^�����P����{.��v��������'v�V�xb���n�$�$����r��b��%�;�����/����n��@�,���T<P���﫢�����}�K�&�Nn��k��7��MپsCI���d��w[.���ɳ�ʡ:��v��7�婚��\��Ӌ�ql@6���@���L���SJ!�,���Au��Ҭ�X����BY��3&�L��,'r�ƒ�]�!]^�ӊ��G3�f��^�4�ن���N�q��p�X�0�Ψ�E\y&�3b�.���	�A@b�a�W���@&�B�ʚu4�B0�]����Gň������6y)�o�'t��k�ڑY�9�$qt��L�m��dȶ��Š��J��w�R&����"�K�?�=}�C�|/Zξi]ClW��Jc�1�uߍ9��.�l���TÏ���S����ma�#��� Y�?)�G�c&	��y��[7�tї������|M.�)��ꯔ�.˥��2�{KF����U��3��47�FT��F���,��JX�5�Q�|�,*f�݁J(LH�0 �s��^;�}d��PR�cm�`��q�S;��!����QH�u�Gn� �O�@�!&+^�u�]���"���q �(�˶�-ҧ��w���� �۰��k��P�]�/�~�x^�m2�wk.>&*�5sg;��e$�6�����if�8�%�sq�F/�Yg�-DdB�1�CH(cZ�F�ٜ��̲uL*�����*@+��vױ�iSC�}�Q���ln$�<���)�u�JC(�e�����dY���qo�ޥz� ��:ߐ�kW���)�=bO'�3�I$�sZ�S�� �����������rkv�V80�2z��G�:4|ʠ�G�qE�X�w:�Kd"1B�i��e�;�ó��B˥f�C��q�pa��F�k1H ��|F'EWа�(��� �A����{0U�f�M�
��w��)lh�2�]:�U����v5rZ�S�:�5Y	��t$�5+Ո;�4�3%1S%)�
��vN��ٓ�L��g�[�EP��C~���5��B��9n��ԫ�p�>�~7:,���@�=�!��Ē׮_冰��c�b�:87�]���5�I؀,ǾRşpl��#(�^�n�*K.�R�^��� q;k�vXkTŢ��^	�\���^���9��L��ŦR� �����zT~ډ�5+���<��?n�k�P���Ia�q�fC	0)����	�d��Z���g��0$Ds4G�[����,������8'<\��q�43�.�ӎ��%��~���U���j����ҩ�H2��YH~�^���xF�Ud���i>���1aT��ڔt1���њ��z2N��D��W[�>�6X#�`�us�;)[�-RhODX�b�Y����~�{1.-�zX�FןV��K�U�ds�\5l>��p�4��S$W�>E���N��\��v��2XN�䡦%R@��XS��i� ^�a��(��4�e�`������߿M]!\pzp��Y8=�Qp��5!H� WѠ_����>H ��.���c ܗ�6\��8�n���`oܸ)����A���Z�����s���^Hql�a�;�?#Wj�vԫX�)���8v,$�9U��	<U�/@�c|v�����H��*�g�9{�lxg(�r��i�]GR��Bܒ$gb˜�d�j���a#,<����6ԉ**�k��(C����t��}��$�#��4M^��k����d]�UH�����)W�S�6�NWXW-�U��pHKWD1�r�m%�Aܦ� ��_����b"z����`�GM��a�����1�;�=��)�G����{��Lc�a֑��)GB�v���W��a,[��R�,=���g�=z�c�B�x���o�H�԰��:�Q�,�P��ͦͱ�A̗B�X=c�b��
k�f�1����|���R+޹'y�<̢$�
�D�Ê)�E���{��p��;�8jஹ�H���U��.�ɖ�x��):g����M0�*/�ׯ[�K&��QY5w6�"\����"9X-�pYA�!Z���Ľ�x)q��
d8��Č���	�VM*�
�س�	LX�C��P���V�>|#lHQH<秘R����C�U��C�L ���7���7�Ggc|���4��+hb���~i-�汘@Z�դc`r�=h�K ,�3݄}$�0l��1
��Hx�hq�Z%�&TB� �9H�z�;ӥ�A�lS�ϔR8��L�&��}��I� ��#�>��[1a��J����ԼF�����[��x��乣���|9R��)͠86�J;-�58���}L�c�B�qٵs�-z��_~�Uy��W���P(���[s,Y��������9s���N�A��X���YF�P��H@�f0'�}Y�w��<K>$ī��zp�8Z픂�*I�|��P�\��PUӁU�c�L�::��` G�`/�K�9B. �B^�`���>��S~�R��S{���m�>��c�$8�������b@����,8b �b_J�K�;w�UH	2�d3��N�,�MS"v�Y/��p0Zn+�s_�H��]�x�^X3'�&�����7�"���f=p!��˫[�2��-sLK���EaN���vZ�8~(�w�v�1�����"\�a|3kݿ��&����]�|M�֏˯~�۲}���?�����tx�æ�8v��fy�-�,Z�T۴LMt&l�%h�&:'��-(\�%yi���!ܵeT֯�$۶n�*���jͫ����z�Aإ?NK���rE��2;��&vNn�)8O,��IY"7^@�4/E��K��b��_|�6�u>Qa����W�B�p?~�X��"��	�����?Z'���²6,=n+�&
��a�ɉ����o��b��-$G��f.�ɹ�J�Z�}|p/��-jwv�����	��;��CTA9�H��p�y-�״֣���S��e��"����o�)G0�HiZ?��q��7�Me�G G�[C�
���BDD�|fv��>R�����;r��YՖ�����r��jwʾ=�ɺ�U��9+3RP�W��q��[��1Òpt2*[98z�Z];XT����f�8nr�V<ܶiH��F9t�A�Pk'��3���Uo�`�vvQ.M\U-vL���$�3���֓ :�r-�d��^F���ټb���}7��>y�ynp t�� ����|=~�J%�7O�oׂ����y�b�{�x��h�{��m�����B�����⚒��z����Q�������d���F�#Ǧ�~�IPt���u�M:�quINjٶ�0���vBD�}}�A��&��w��^��YZ�ݣ����Ȋ�L��..k����V�)�
�O�:|�a���'H��������ҫ��eu.�J�2�� gϟQ��S~���X�9/�T٩�T���R곭oƆz��ت�ծ3^�hD�d�6��B[\�'������դ�g�ԛ]*�P�.0�E
�@�]�a*#���3��u�ٶ��<�����sRj��.T��vC�Շ}Tz�����˺O����~��r����~��Ơ¤s�?�p��ˬ�m1m- ӮM���[m�>�45��/ȵ����＋��ͷސ�_C�:�ؑWH��� ģK�j��=L��)�
��6�x��"���M{%��M�|B�aLXq����Ve�:�u�LKX4���=�j\4�Ê�)�ަ��;������UN�tҧ���>����6F%,�K���Rkw�]w�y�����v5`�|��,�-J&F��y�L���}w�T���{ޮ��-í;
BH�L��h���Zy�XiuX��dK�0��V��Y6�Jǖ�A�$�"�S;����|"�U��� ]�vS���W;Rm��t$�T��ͳ�	(l�43Kr�{������k�Kܢe��BKA`����蹍�QV28�7}�d�Ӛ�1�	Ԕ�AC���z����s\��u�ò�oh��J�+��C:�<���v�ѬMfZ��_
�Hqk��bX(^!7w�j�4���� 7�rdn�U��ُ^,R�ߠ�,w���z�igѮ�Љɥ��&�WJ��f�}�o�.)�E�Pw�٥󴼫Vg��r�����O^�����1��u:>���F���Cv˺�^�:��[���iW1��VԄ��eN�$�(n��:��(j|�w����o����N	�9�N �#X�'�4�̱���d��r�ڌ�\�i�N8p]Q�2������?�}�w�CO<F��u}���K�o!o�0;C'���'q����e;�Yi7���ve�q���v��`A Ip���4I[�\�U��x��U�TIJR�H*�@�~�S�����vTId��%ڤ,��IA�H;H�f��|����4@p��,`fz�}���{���^��̈ߡ�� ^�_�b��N�o���1��w���,bG}P�ڦ��\�sc�@[{��L|h�iOxQ�eZ�<�L�4Ă���0����4~C��D�Vmg6ؽA��1�9]I��D�Q���h�Wo�P��f�ay$f�=!�6:9&��;�gN�K/�,û�eyq�4�rw�+��O�%O�8,C�Jn�M�6?J
P��@�qg���b�E���<��2
r5L��o\s�.R|���K�=1�h�:ډ�5�D	��w���3(��/O= ����2��X�吭c&��c�չs�CA�M����f��ay��W�_�3��h����(������iv�1o�Z�uq�;t9��˖`��HC���f�����Ia�;A�lXJy���� ��y��T���O)�*x:���|�΋�lf��ز[k��\\���(Tb� q�,Jb��K:������˗i��{}�2B1MNu���!��G#B�N��"9�����%=���g�*�n����56&��Ưd��4?����eb��[ϟ��O��;K�֥�^�R�<a�.m��"á"��1:�<��"���p�273)�����ؖj����E���� m��&�pqK;�pj�u
x>�Wz/_���yT6 ZP�}��'�ԩS2� K����a��5�%���I�5��V��3<�ŖFcة.����P3��TY�`��v���)��8@�Ft΅��bb�Z��f� �=P�B�F�Q�[��		�qq��G۫�{_�q�4�4�
�*�{��c�h�G8^�
|���$�i7o��[��Q�X[�����?\$ ��+on��m���0e8#*SU�Dz\�ʰ��J�㺳��k�E���7�c���G��鑥ŀ�8vD��k�e׎^���R��B�&̤���i�գ�	;𰗴��Kͻ���l��HZ�wH��o�J&2� lg�q��m-�B�YΣ`V�
"иD���s�ضo��K�̬�R0bF��>� a;|��T�޺@%`x���~�����w���Ƈ>��{D��.�믿.O>���۷��C	)Y�1�LM�����L��T�f�jP�H��Y�"�D9�,���m���S̆�|�R|/��%+��a��y�F��;�a��4)�R�z둜w!��̜_���Os$����|4{�m&c�%eqƃ�ӟ��s.'��ب��|�9��]�Y��ԪU��7�.�\�����3��<��!9�wH�����/� �ۀ2
g%R��PT(��pp�H���dJq;� �k�ur!��)�xݫ�y�XBd�m̧����������ʓ��A�w>3Ӊ����ĸ��?���z�e,������>�l�؋/��7�h�λl�N�g3�e�f�]�!��9`i�������#���N� w<�He��q���L�h����1H@ �����4�χ}��m�m�c�F=9��ˇ�
�H�t2���Q$�21�AueM�p��259-"�D�5�l%���Bn*g���B,,��X?၏��g��1>=%C;�;��Rvgʝ�O��]������C�s;��5wb�'`��"@'�ի��g�ؘ���x��Y��Ua||���C�t59}^��$^���}O��+�8��@����l�;����m�N ژ�1?����_y�iy��e߁�e��y��X�Q=!Pgי�}��{M�zU+	ncv��m�U(������:b�~n�J� B�3�U29�t��/�_WU�½ߐO���z�ƽI�Z;�qc��,�J��m��6f;�wZ]Ӕ�t�(r�̢ʦĊ]���_�,��Jb�O����VZ
rK�H��
<����������e�άLܺ)�>���~D�ɺ��/��7�֛d�ڔ]�{H�^_[��r�q2ۘ�<NP�DEXH8�r`�a��6��:z��Z���m�U���-�>X&�c��k�":��Wd�������eW�����J�e0��Y��b���'乯?/Ϟ�!^7�2�޻��%w�N��3΋~��r���|5��a��f��/7n� <:f�C_Ô��=�ƞ��*�g����"�1�]��>&5�P�	7N����Uv�`�sY��|iÿ���x��F��Ռ�#��zVSq���:���FC$D���&��A�xR�U��� x�<�$�j��/%\�Y] ��<I�
��wy�+_�_~E^x��|��}�m���g��4Ϥ�r���}gk��&.m$E]IÓX��i`L*��QPz����.��J�����\���إ�}D� ��Q��KB���43�ew����
U�G'�ey�A�����*�_~I�y�aT@�:/
����=��wr|B�����s��vl3�k}�g�
"�!��֠�]���E&h@?���̹^o�8-\�u�L��:墽�X[A��|dG�+4��bW1r���Ν���@�F�邎-�P��9�8���}ݕ^Y^���U[�aF�`;�$PQJ~Bg(k��F�`�����Tjp�~(�����|�G%�O����s�˳��7�������z`Xο�+���-Y]_u�Ms���	Vשl=��Tu;u�=�T�0�o���Jҿ�ds��$�&��UM�e �l��e|���'�����A ��9R����ҥ�,NC�\���T����Ґ��%�ƹ�0�/z�A��9QA/��%J�mK!�3���׳��ZJ�A�>�h��d �C��k֏�(ī��R��<Y;��xo�`���a�Ɖf�����^�ٰf�*���<=5I&4N�_,o���7^5?-�C�ύ���ŉtt0)���������ݳG�]��0�����7�3��N���-�ӛ��
q����û��a�������gm՗�B?S��iJDg�@�^��:Z�.�_s���$�m=}�����	��q��,XZ�&�R��2���ȭ�E�����̲�Rܡ��:(F*�z�M���2��Hv8�R�λ��z�ɩ/����qշY�'[���m�h+���P)��*�n#xVC���f#k��N���%� �㈔��uc�aL����$�1Y"��Z��әOQ �LZ~nI��qs@�S(���Y�R�#��\ˤ��"��vd�-��_��l�Ν��L@�_�����Ei������#��������Y�ѿ]����&�[��ʲ�����L��ˠ�qD�v�#�CD��� 5�?�P����Q��&������qf�
̋��d[�N�)��
���:.u�݇6ò49 �2�z$��f��+7䝏� .�6E�R�
�D��={�?y�J�W>�"�3$'��� {��Q��;���w��,s�͒`�;���ڤ�M�F�m`�%�%;��:�X �˺��J<<2צ3p,������^)#�SH�=}�!%C�݀��p!���D��.��ч79��@����}{��2��4��o������һK;ɪHm<��_�cg�M27U�ì ���7��?��?���@@��̯ʇWoH�K���2�r�o��C �B�R/j��@�Q�Z3`� �=ia~�-����.�Z�9�5)�`<���� ��ʺ,��d��������'���a��e�ű ����r�"�җX/�����~Yq��L[}�fĊ�{fzJ��`ۜI!�\I��Pp�2��XmNGg�M@e�a�����2�v}�*@��l�2��0
�Ѳ3i����T9�-����$��*U���HA����w�0ï*r�f�ܛ�*@��7[>���P�]˻s_��}����E����á�b��<r��z���wf�H���)��C�����Ne~�!��Lz��?~T��J_���G��!��F)��a�׀��:4HC)&x�����QXm���lS�j�܇U}������ܺ;���Y�rXL��Rk�һ�B�1���VL� s"���i����N
D ��yl ��Go�RBP��↎�i�oe��n6�~VF<�<�HU� F��)롰�I%�C�cM�F�����#ik[%c4`H�d	�#u�Z�u���
��+˘6X�ϑg^��W�ݜ�������C�����5�W>\BiFj�������+�
;fo�;O�5�0}�dh�^2���ޔ��W\�B��ZN�O��{�aٷ�[��$�Խ��n�� � qGх��;W$��J�ZK�W�MNe�@�^�qD�~<"��]�%4l�DPz���
�Y{Vk.��.T��r�J��Iĸ��]��RsqǬ[���t219E�$���ǎq���ΐK.���e��2Ļ.�E�nV�f�����X������Q/���k�� �Vs�I����������D�=��D��P��������(�H=�2�|V�N�;дh�j�Hu:�~�5����n�0p�� s ���!I�9�S{�qٵ{�|��i�� �����������*PW"���Y@��-�7�]"���Srp�N�?< ;�ܽU�k�=E�<�X�5�i{��������c@n�B��4�q�^iqL�.v�P��=��Ȯ�E,�*h���=z�m��JtZH��'��~�.�\���;w�mLʂ����������Zd�X�(���e�x.7�V���;7%?��A�R�6��1:zSR�� �D_U�����z�A&�?3�\�X �(Öm"�Kfk�#Ϩa��V)G�M	F=����,�X4w�b
�D�ˡ��b���E~�)��3�Z��c�ceE$m�_����q�y���nŻ���A�20�Z��>ߒ��E�^s�y����B*��]:�O�+�Ζ֝+�*$���U�{bΆ̯�e��Q}6��&"UK��4�6I�"zS$@�D�m1	g�O���9t��޵�?�l�-	�瞓��s^��1�T���?yl�ڃ�N�/�V����f�M��'''�E9�;6L�B*{rj��\~�m��=�X��#�� d	�"�5�S\��O��,Uh�M�8a��F�m�R{�\�xj_���5 �zm����A��ا##�<�pcfw����ʑ�{��S'�݋o�����D�C�%�-�,߭LJ�҄D�R�J)��(q��B��J߃���yٝ�kR _�h:����q�5#��(��-�Tc�JE�����td�0�+����%���z�o6�I�Z�ߝ?/#�^�׳�%*��yЖ�������K>6�gj�e�si"X���e$��{���d��;%Ո�~ԯ�H���G]��H#1q걬��Fӣ�ُ���?l��[����{��t�.��*���ͱM�k�`�6�G$ hb|��A�b��410X��fL�r���T.L��hZI�/�ي[E������δC�v�Ha��.N[b���Pj�T�̴4�qg�k�ɒPFg�T��ȥ
�j�8 ?x�7�I�z�)y��<a\���{��>x�/�Q�8�>\`��>젾Ӭ�g���k�@�� 4��H��T1���v[�Ї�һ���%{�-��Ԉ���{�z��n�$�gڨJ�iu�_�#s�N���������[s^x�1���3_�_��W�K9��lk	0e�^�n�! �k3%K%Q�C=9��{P�φ�[=��DC�ԉ���_������D)@]��Q�L)����n	Mb�d���z]̰ȁ�[�V���dx�0�,a�8�ɩIY\X �u�<P،���2Z��E��%��Pޫ�J`m�r,���2���6x�-n��zՍ�Sɒ����\�$$n�"��\w�F��{����<�b�4��%���W��u���$�8��3g��^ ���jx��YxRk�yu9
��J���h*aC�rQ��[T@Vc�ɂ0@3� 2����P{�S�Ó(�d3IKg�ee�H�� Jڅ	��n���+(��ς����2O&���x�zz+Y/:o�f��n����ȓ��:͈7�V�y���HK6B/L`ԋ���R}�m+��ѫY}ֶ�|�Y����U�6��k�9����6��\���wg�G��a�-9��w ���`p�y-}������Y�t��� �^�^�~eh�TM��w�K�{
��-�Pj�D�$��4*)mGP�$���[���cD33$3\4 q��+?gB��r~�'(��{>87Of#�퐤�_��$b��\��jy�7�
��yc݌���l1����oͦ�q�Z�ۦ��N9������=��GMa�Y��;�s����s�!'7=e�=���D�"��R��-�v3���һz��0�9���M "A�2��肐M.d{�͉A�L�� �X�CX���}��nb��S�h6��hֽ!�3�i7=��>2����|>�� �-�-ف����<W��f�M�Yi����Øg�Kබj"l�쳬eT<��cB���s	r����=� V����zG`�v�Y�q�i��\�q�aౙ�����@��Zl�J�eן�����Am��m�i�؋n�1�!�� 3��('@�Fk&�I�v5T���ened{�}w���ez���5� ������&��Z֊�{��B�1k�+��4R��km��<9��a+��nܽ�t+��y	�9"|��Blv��e+G���/����#�t~<��-�%�~a�T�UT<f�*��UW���)�&^`x>I;��}v/��]G� �����Q�C/9i*�*>��\�@@,>I��"��T��1����(��٭SXG��^��~��I�e1�_��e8Osm��uh�YF��� �,o�y:Bl�xH�yO{?~o�]��,�W��7(�:���043"Y{�ͣ��0�c��FQ��l��>�f� 0��O��㴃w R=�3��?k����d��hP�*����'�ط�� �(T�%���(�9�1b�A+�4�����ó�kq��-�v�l�Z"JQe�I�e
J�1y�}[6���)%7JP(���佖ye3����I�N��g�C���{,�0���ݸڛM.5�����W������^�3�n�r��gS�0���L�`^�B���l����A�ц�D�{�
>֏=�@y����g����P%������f�y�kU���_8x��J�?}�4�a�}vM�o��{�q�
�#{���7�U��`�.
�fP7D]�رc|-�c�@(��=��������	D��7^Vb\�k׮��_xޏ�b�T)��9+�k��(P渹���o�)6 �q\�|�3�����F�^5���A����5/o�a^ڒ7l�}���<��m��y���p���Q�`�m��w7���O~_����I�]
!u�y��ǂ��v��N�F�c���1���A�� �6?/�4��׌{w1    IEND�B`�PK
     w�O\ےtR�2  �2  /   images/6a650d67-2f6f-4705-ba20-a1e007a57e5c.png�PNG

   IHDR   d   8   �]�   gAMA  ���a   	pHYs  �  ��o�d  2SIDATx�u|i�]�u�ÛjU�*�%�&4#!	����؀c�1�c��$�+���G��g���W'����86�c@f����,�J�y�z�p�����ާ��'U���9{�o{8�ݴvU����R����R($�}�,K\וR�$�m��8�y�ݖ p��'���q�plQ�<�v��JY<\���6�K�j��Q�DB���� �lVj�y6����z������T*z�r����8x�o~~^%�sZZZ��[($�L�\O���p�%�XL��1��z��?y���y�}V[[�c��;^������h}�w=�N��6��<�7�wRr������1\�J��,�_�%tn&������MNK>���27�n��@xSX`��qL���|����P|�S��x����ֶ6���;dŊ҆�9����
Ei�OLN�g������;@��{p"�8ojjJ�\�"Y��/c^W�bZR,���oGG�
���Y������y�\.����ͱXl�q�������=��挲bL<�����T2�
�J�%W�C I��[�X��͍�zkP�J�Z��"cr|R5ײm�Yd��R� ����%pS�����.B��x�q,ޫ/�"�;��qA�M4���F����N�9�d������ÿ�h|MOO�x�8�ݜg��D�ttL���
��9�ܗ�S�����ǿ����	�rI��w�&T��K��}yn6���aiF��u�>�W�CQ���aŠ���YO3�RcC�$b	��b�(��:?�-�x������
�3xF�8���>�����^�|�:(W0PO�,�8O�d<��sc:pN���p�"��>� ����T��X��S�qU�˕R�DF���F��ٳzU ϯZ ��}�����>-���=rL�]������vu��䄤�4nx=
��rB�B�o"�N�h�1q�)(�;66&O?�s�����N����w4@���Z��s  �	-Gof+.�8Я�B�s0N`,����?q0)Z'G�Q�ǛZY��[��c�f!#E�1\�h�z}�6!��s#+�^� B.����q�e��
-��s��?��Oĸ�E�z���{< ?��$�������^*���ŁYg�=Ѓo�~�	XHMҖ��'�F�|5-�E��2K/H���X(�Յ�B���X,L�R�G��I��iY1=�-{��Ge���綾��ÇŃӣ3� �Lպ�[tb�N�Rl�p~�%��m#q�rB��w��\X�	��Ò�Œ��B��J)����5�Pഈx��y�e˖ɶ�[eӖ-��?���o���桷�Ȗ��"�K�k[����x�S�6��p ]��β���,��H`b?P��T
���~���wﭺ�oz��U�pXhX������T��α:ʃo�!�Μ�cG��o��y���u�36>&O��gʪ��7m�$Ǐ�
$Ph0x��+%����7�;���tvv�'��W^������S5I@%�(�*����������(�Ч]��:�7I]S�tt�d��y��L���O؀�6�"�[8^X$��1^�K�n��x�+��!�,N�'p�,��4��|NM߷]�c�N,�����Qn޹Sop��9��)�����(j+a���LLBM����f߻�*\P�n��f���OKo�Y��N����|���W��ky�}
s�B?�>�6�@�S5)ٹ�f��?�Sٽk���x=��C�ēO���ۿ�����VT���A���TY���s��3�ʑ��Ŏ'��?-ǎǚ:\{($����8�_���
��ʫ(j��P���ݻW�l���LM	`֠��\�[�P�W�����/��s:��p�o�$���'e������,�?������/�v��L����5@�s`/�RY�V8Aj_�U� �����Cj���ڄlذA��[�4��_�X⡏1D=�e7i�[w˞={$�q�����.�a%�� ���ߒ��z�J�W,#��M��X���>�---�r��;dbjZvܼ�ȓ��Q��sO�ؚ��,�n�V����U��n�ѓ<֞�t�̘�������t�v�6.+X�D֬�$����[�xuV��(���_xQ�Z�e����w/C��!dm�~����?jx`�~�e�.ٶ}�����������1���&��իW!�4�nr����Y�v�ZӦ�eqW��/�N�����J^Ii���ke㦍2�k��_��g��u2�wB �Z��c������%e>v
W-Ee�kѠu���� �k����C�~�/�/��'���������&y����O���7&J؂�uz�����[�RF�9D䞑<�c�K���4���{nǞ�ǟxQJ8&>51
g;%g�o�d��x[�L�$;�o��W~��288(i,2c����/|�r��Qy�_k�B(� ���SSҾ�].\���A9��e�~+4	�����4�4���s��$R	�(5w�ҥ�p�qP�y@��ai�v���4��sٜ2.��~�nYރW`��4��{�l߾C~��˱wO�M{o�����V��%��g��|�����ZE��>3J2l�;(��5Ȼ��O���zq��� y3��yhLI`&�"��"�]�Xj1�ټܒttw�#_yD.�?+��ò}�y���[�%�@��(zN��oy啗�)�W����T)��=���د��VSA\D'<::�>�L��بaEX�/<��z�^����+
د���]E��σ��eTvs����E��RhU���+{��r'0޴j�!�*����PҘ����r�d�t��Y���_�{?w������'�O�
����K�x<_�)���WT�!1�?�5��Ϡ���i�j���-�#NhPm�l>��z�Ia��` �n�EvB��._-�.^�A^,�֒L�Ї��K��+��tA,u��������viz���ZX��U���À�^@����456aA� ��RW_+7����	hwZ��`�E��[�V}�	@�r��9�|�2��cJ��D�{%�ӟ�>�����B&��:"�	��u{�?�]`��R�ӟ�LښZ$?9
�O�Mׯ#�Zd'5'%���u	���P�\��@��U��������Z�B)-Dׁ]�2Y$�ܪ$�d�2X����Z[d�0;3+%�o�i�$������N�_�~�,�Y���C��T3����Shq����Z��?%���g��k�Ms=.#c����+��O��|󛿯��X�؆pW(�rHc��c�����/��H1�'vlݡ��'��ahp$L���0ׯ�I�>���Q`��y<9��i >�gm�|�C{�7ə#���k��@�3T�rZ\��8q�.�	J���.(	|�{��i�Z�	�S�ţ� d%?�Cå���s%gw��c���X������K�<��V�f��g����L�qt ���E8�U���A���>r����������5k�`s�l��MR��g,���ʎ6,J���i?�x��kI�b��<�'�y��'g�*�Y�D"��2�.����F=��n��kM�0.�%�>�K~��z�QP޷����&���� �6,݅��e^|��H��"�#��19��R���DT3��̂�pr���{��c�ҫ�%�����ld�k����y�6�lhߣ	5�b��AOL��w�ר~qw��:Jgj&��j��hfL�̢i��k�G?3�eά��y<�¬���֨aDli�����dd�6�^���n�䡘��i{�A�5�S3��	�+ʀ3𭩍K(�,�2US#�We��e)I�g�r��1ٰ�6�-�-�h�<2�XJ85��+jZy�T:��0=.�s�i��TJɅva!_�<�B�L�1y��=��
L����#wB���'���פ�j}]���LAP����/+�/Wv�H�0��5�	�aP�|��� G9h��)(=�*&��A�ϚD�T>�L��X�}��s۲Uؚ㲙�4�G0W 4j�CG`Y�c>����ɠ�տ����gO�>l�l�t�|����ȁW���7䕃'eò.�w�6�
��ʰ��+H	R�}�jW����X^����Er�H��qQ&����)L�b�p4�.���,��O��)`������K
�{�%�C ��۶��?�y9~���K�ki}1�:=;�ME[�b9�C� ��\@�Z��1A��
p��2�JA0��-�a����[��Z|	�j�ح�7R�'��岯,��N9��0ىq���h.�ק�3��V9�0{l���ދ��b��җY��7^; �^;,kV��|zJ�VWG���3�:ټn�4�7!������W��PF��5����4h��𮌍�
�5p�D�Bj��ڌ�5�nb���g��*~"�:;���E���;u�1�xI~�����d6ы��0����_E��Z��V���4|�
B����B`����Qrܪ�2�#��%��D��Oj�P��ibI��mc}Y�;彁�t�^���k�W7I�@�Z`���a)8&�4�`�o��;�I�*�����K�b$�>��d ˭Q&���b}Y��X�2:��L1.Y�,�v`��Ā���4��B'A��p��_�/_4$e% �������۠�@ap�	���m$��c������1H����F��0���g4��J�)��6Ag�}44�Kܩ�{�����'k�t�Θ�^̆��kꕾ-�k&U�}f���3�Ψ0��BSߦF����e�նM�^3��`3��\��~knq�찐.8a���Y%����dQ����W�Б3���n��"oʌd���LM�4�k���
Dk-�I�3�p��i9��>���x'�1Y+��15����B��q�����HbA*K��dr���뚤��^����v`�N�1�;�1�S/�MI(	�ecǰ��	m͸~<��4-B�y��:eV�B�D�VX�3ǁe�׹x���Y$����f����{(�Zs1̐kYO�ɲxc�b�f�M2۞F�����/��H�|�88V�`v����j�\���V6y+q��"�'Լ��:���i}���o=���l-�����^׊���@�A?P,Ԫ�^%U[�l,
R.���TSa��E0[�i/�0k����󄴷Րߨ��LP�sM��*�*�g�
�5L�o�?��<���7��S'}N�bq��565i����EK�]�X!�#.��`]���$���R����.</�ۢR0O�_��B.SL��&��g�_��LNOย��E8�M2R0s��Lͳ؟�`sp�s���>�aY��%�N�i�Hk��h��7u泘if��SG�JՙNa��m�#�<������� ���ӂP�B�>���JK�2@!�@?)�����7b�
t�Λ�O��O�(d
9C}���{�ʷ��-�aS�gAIE«��*/�f��E֘�z'ó�g��\�a1����W���@��OܹQn����7��)�X;Ǆ�f����˲�`��{iJ��L!E��Ͳv�z�_�ChI�򚑥�LM� V2�z�b�n�F�V_{C�c��X+IP^��%P��2�˘3sOt��5�j�� ���EIᏑ|��5��ha|����3�=M�5��C#zJ�%Z[1׬T魧uO6lX/_�����%�r��7����&a��ЅVqfv�k'����}�GJ�ˢ�:Y�٦>E�K{@�h���a��%��ݙ�&8+�$	�0%S��[>�s�lߴZ������g��J8��������W��Vj���_���L�K*n�ʲ���䮻n��E-��Z�T��Oa�j�VaycS�2Hih�������>��ւ�5�N[��hS�[-0����'T@,��@"���R�G3�aF��ZeQ&'�4���!�۴u�|��_A\�Z�uJw�8~iq0�S�#�e+RCc�|���t}�RV�|�"D��-��F0�f=��@ߢ+����`dC��.]�ZJ�n�x"�$�`X���I hٽ�W�n���_ɕ��vG�9���r�]���˥cqh]���s��	΃��a�K�'� ����2�����M�N���p���R�%j ��wfdy�Iy�
g�e�(�������(��a�Ͱ^�z`8�jj��d���`J��L6�9#Z(��$�s��]�U���5��c�lL�~��`��G�,9@�>���o�����^����r�7H#Y-�,|DJ<�B k��/���^��߇�3��&�ՏkJ���edǖuҳ�\��W25=%����g��|�����1y��9�&>�qwGR�{'��Yu2��0��tb6Ο9��G�$֗MW�eš�)��q���Y׈k���f���U�ʴ{[�Tf��;����7�n��JO�䵾3V��g}�޵��#W��V��t�<��%����r|bB�}�Yٲm����c��2+�pK������MRgM���'����
�Y *�!&������9q{�vJnvx�Rlep.ħ�qл�,m�����5(r`�7ݲS�����q�+k���ٓ�$=U�b9RQ�b�T�|AH� 3�Œ�Hv,&�Q^��L���,WsR�c�2,_��I���ni�0�q���n�ÆKa���i9*?T6��&�
0[@P��q�4��(dz����b@�\'S��6�~�����Y�	(�\����8q^n�amǂzS9|�I�ol�Ȕ�d�v�Ҩ�;�/nc��8����wX��$�+��vN�������8��dE�*�X����]����U���+�7���^O�r~]\�
��F���Ki��`�@��.K����)�H�RP�`y]�&t��;��K�el�!�m����xLsIJm˥j�G8db��Ě��O<)_�ʣ�۵Z��ojjn�|��d;�k�P�0�2�>�k�a�L�̧�Ҋ�������EӨV��y+8��^&���`=�-^)���9Yт(������������fR0�)篎��IP���-K����U��Izl^.���m;�+=��KK=n��U�haq�j6]�pM&�����([�n�b�21�ᘗ0HK�F/�xEՒ	�bI���eF��;�:�td��{%�����V�L�Y�(�<�
�ma�U�g���:�G!��2F�l��b�.YS+gϜ�2���O���Ř�@��^��-B�7膢W�t�Z>���8�H��g���(��nG�"I�u�nK6.��[D�j��2�Ԍ%/���ep!.�%������|X����Y���;�#;�o�B�����K���A��y��X��m�t����K���C���_�CcZ@�o��<���~y���I{{��ݻW� .c��EyƎ� �&�ʟ��	L7�f�5:g'�������?@Kz��/��m���ʀ��gÆv��:wFr`~��;�������LMLʹs���楈��C�*L)(��@k��l*����Ro�I�j�8����	)�	�0��ɢ�qȫo^��׆�[���A��w�+����!�m ,D�E����'������0���FON�JsK�g�KN+{s�i흭!���	�h�da&�EV%�����y��&�0�V`󀘎]tXV,a��j���~1
��O��hI�.�@�?{J�~��/K3�x�`�D%	g�7��v,�4��821W��o���K��J�<a�#a��7��̹��Nb��7,�pQ�I��m��oedxhXҙ�\�2%�.N�t� �,ܟ�FF�@�&M��e"ߤF������4�+�i��(�wtc��������J��l�&�{!�a���>���K�X؃�|�J��=�4[�V��K�ddK��f�@���ua�p]}�:w�W�\��ź��2>�98�_��Y�`ߺe��,�a��KCa�����z���V8kX{ɒ׏^���Cr�dYG�$�Q!�9�
�W쳔S��,�;�7ȡ×�h_��.�l9�f�XH����m�I�NG�8?��V5,�Uf�[0�e|@�þ\�ă����6�(�>�����:�5��cZZy���7�wQ{����PYm�05�'��Y����H"A�
��N( �Եfn:�կAp��yy�G?�L����&M��؏���~V.^U�\��Ͻ ��K���/O�|Z�>5(��ڥ��FR�eJ��-x O��+��[�%C�+2ŉ���g�`���@*��N��U�eِF!����p��vdp�IF�a۽:A	t��nj���ǀ�w/��+�ʄ�%`/sM�y0o���[��������F�N5]n��.?l64U=�˵eW���`)�c�X�N�m!I��$�wX�ϙԌ�ᥣ??���1����o���!��- �I"�L�(^���Ɂ9흮�i�W�~%l�&�� pq�<+���	���VPZ4R��	.[~�Y 'v`���U�߿��L��`R��l���u���-���9��|��!4-OjZ)��b`)���ƹ��mt��f&5)!k���v�#�p�p���e��q���D���XI��Jz*;���w����
��]-G;aG>�x��El�2F�aF�*�f�Y�g�vr�
ǳ(�d�eĘ���WjL!���2Qf��0h[r�AqJE;ᙆ�4�cY1]v��~��E����~�i�_�HZ�۫�I�zD��l���]*��k����1<wႬ߸�v��+N�n䉻�vh��|�,�B
�G޾����bht̔�4}T���1�M���h[���v�0�Ln�Η�w@3�9-t�_���IeP�"ZPcY�JVV�ǋ"��2عh��p�*���$C^`{�eeX�,�p��D�Z%�|�

v�M7��ݧ{'a��V����[~��U8��m��%��I�"�FQS���bG�Ӛ�#��ָd���`4��FKÎ$;J�O1E��*}5�&�S�n�V�)Z�m���a��~�d����QYL�͒\._m|�����)3cʢ?+A�i���_���Y�#+��:$�?�=y��}
���k�2S���ה���H��cR�p����k�zٶe��"�+�-�gK\�YO�G���r�Ҕx�J@&�m�,�9#���9��K�ʃ>����c���A+Z�gҏ���ݺ�ߡ�R#[ۛe��*�_xAn�{���mW�A��W���AJ��D�e�B�c���4]�pc�����
�֟�����E�4*�YN�'���}�Z����B�GsO�PL��������s������o���8-�()�]���)��l|��^	�) �J6]�����-��g�4��Uʀ��e$��蝗�����k�%[6ZIlL�W�h�tu�<���͛�J���2�2�*����ĲY�Q3�TCOE-hU�j�}7��K��'�Ѭ�n+L@�9��d=	��l��5����Y�5�n?b�aÝk5Ȣ��R���n6����J؟�c� LF&�:wKji���ځ���C�;�B�g>�y����}eW����#�7�HcCR!9� ۪kTB��Ε��#b�)�4��;^p5�b�������ʹˣr��&��N�:%�˽R��$M�Z���cK(���F���,+5��<1U��ÿ,_�L��Ľr��~9��~��ƛ�P	���~�-��uӤhM��)M���چͨԴ����j��S��L/��
˯��-CխJ�=e��T r����\F��?�/ٽs��B|T.�b�qy�|����k����x�Vh�)L6�}���o�;~XVv��NwͲ�e3]��H�L��+:����o�M)x������)���ɩ	P�L�����6��Y��"�0�MrA[�N��������v�u�fٿ�u�&v���m25w�6W0uh
���],f���Z뺦�ghy�׶��"ٍ�=��������O��E;xM��QN��Yp?���3�^�X��.\ꗁ��R̥��5%?p��y�Ji���͎��b�y�t�䳦Ϲ����n�� 1�B1=�TB1_�&�@��o�/�/m�
�١�7^������|�����F9��ۦ#����������bmT�g����5�������d�߭9��N�Wt"4s����uL1�� �jAQ��̤�d``�l=��>}�*(�5]/�j�L��̪n�6T����n�Uk�!�H�mw�)��3���E�9X'�����ׯ�2K����ú����m��=>Cw����QzZ͐Λ�nPQ����@]S��Y��a�.��=�ުU���-���9�j��(�8
 ��n�驟=%G��������{����"���l$`j��.�֫�"L��e�En�����ȿ�4��Uy���k>��yllR���x�Yq�k�M~d��,� ��N�ɞ�n�����_���ֆ� �<��J����݉��S��o5��|ĺWF.I}[Yڄ)W+�DXnm+�U�m�`W�Nꢐ�h2Q��_��lܴE<����ڽG~�̬�r#��������ň6��5�9���[��c\i�6��J&WP8��hSȗ�äҽ0(��z�����9'�nމ9z4�^]m=<��������e9�_�x��*݊X��o�>��߂�ڰN>��O��|�;ߑ��K�5ɍO>��b�[ŗ����%���Q�+Z�9Z܎emb�y �؍�� ϙ���}��GtzqxF��3 y��@7~�{���`�ᮻ>"�bQM��9N��{�0�g+=���Mv��}c�����Iէ+�o45���͘�u�*�!5�1���'�`������t�������<�K��7�ؑ�q/4�pK��G��8'�G���{����Js�"�o���ѽ{������ej&��V��Ђ��/)�Pk	3"x>� *��f%��-��F��u1�32:ȳ�ޒ���R�X�'���?���qM�'�˗-��z�,��+��n�1�����Li�O�BY?�v��l�Φ���X�h����H��Kn�D��ت�`S�c]��qXGN���M$�a��]�������~<��069��?��`�{
���3*���g�X�eInX,i�˩��%�,��6K��2�-�0]��P� &nyf(��y��(o�sY��K�����8���k_�i��ԭ�#J=&?11)�2��B���)�?�r1He����;�E�.^G�	{��E�ݰ7�^'g�Z_�'[-�>���bp7��9K���Y����a�������,d��������IB��6��ظ\��� �(�׳�*�+�/_<*	�Fٴ���wn/V4;s�z�x�r��Ny�Gq��2�p���dV2%Gp�p�lpc SW�,q7)c#�2�K�tvv��{>�qF�������D�'���x`rzVV��R8d���%avF����Q�#��{&3]�������d�[���,mX����[�<�6R��J�����<�7��g>�i[�HF�&$�����N�8x�e�rn0-?~�Mٲ�S֬ꐦ���5`I���!	j��{)q3v��]=*ih�¬�3��F��QXdO��w�=�Ӱ�ѡ��;%?�i�W>}��hQ�n��eJ���ב�W�"yk������RJ|��9}&[4�1�eNB�7���'F��2������5KKK���Naܙ4`/��b�撫~��įf>�Q^�hy��r������%�d��z=kU�8;���c%uh �͆⺺�.�1����p
��hGI`
�L�Y���.w�LG�W�xs��2wŧ+p�,����"|h�L�D��5��������U�z�7�u�k��>d�=/?��&}XAY7��A��&ihs�Tݶ��YE�
/��؅;p��F�lF�Q�B0W���[��W�Y6�e���dye�f��7[�m�T0�5	�q�u��oi��W�X�,'з�_

�E�y�����'�x�@_x��:xUK�L�=zD�/�WM�-����v!�2��BQv��Ξ=������g���/sEZB� *sJ4b��#����Ml������wT囬�O���W�"[�nUE�5?��J�y���QC����ڦ�y�'��{`6���`���Ar	��c*�p���Y�q<��+���Uu0�'��}B����P4IC���Q.+�.F�n�)��Zo��(�>'K�+Z�����ߠ�����mU�������D���DA��c�����?0p
���}C4��׫�k�.�{���g��e$�ځ>��Mpֵ�+a������yײ���G���DQfu��"br<�Զ��/܌�~��pA>�s�-|}�5���NU!�S>���)j�{�0�=_1��-}�b�[��M�GKU"����5<�g��)���9nS�2)x��po�y|�ʁ;�,��h�L�HBJkjv��!v{�tD�'ę�2�{�����ωZr"���"Z���P	�_�0�uիuk&���b?�^�%� �+jK���_HL�A�!�+([�����o�~��`Έ=Sܻ�
��Nkk��%��|E�CԈ9܆F_B��ӏ�J*=�3���)q|1���}��& K*t�_��YE�:\��Z�ʏ��^�b>�p� �����c���/��W��x�cA3;��n������FOq5��
�ݒ�>2I2S[�����I��f���    IEND�B`�PK
     w�O\��_oLM LM /   images/a65aebfd-90e6-4215-8cb5-f5692b012cc2.png�PNG

   IHDR  �  �   ��U   �zTXtRaw profile type exif  x�mQ[� ��=�8�iҙޠ�/�12�,����_ᡑ��\U�$2gN]�#�1D�]�oP�*	�2�%��'����ʩ�z��D�s�.�\�#۽P�B�,�[�.���tT��b�9�g��'6��6����V��J)�U�@D2꟱�\d�HJ��˾\��chZQ:2�B�r9΄�0[zc'\���q��v8�}�������G��svo���  �iCCPICC profile  x�}�=H�@�_S�"A;�8d�NvP�8�*�Bi+��`r�4iHR\ׂ��Ug]\A����I�EJ�_Rh��q?��{ܽ�f��fOP5�H'�b.�*��"�!�0���L=�Y��s|���׻��>��P
&|"q��E�A<�i���C�,)��ē]�����o�K<3dd���!b���r���G�Ê�Q��sY��Y��Y���������:�1$��$R!��
���U#�D����Qǟ"�L�
9P�
�����n��̴�����zw�Vö��m�u���+��5��O�-|n�M�.w��']2$G���E����)��kno�}�> Y�j�88&J��������=���%ar��#�  viTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 4.4.0-Exiv2">
 <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
  <rdf:Description rdf:about=""
    xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/"
    xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#"
    xmlns:GIMP="http://www.gimp.org/xmp/"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
    xmlns:xmp="http://ns.adobe.com/xap/1.0/"
   xmpMM:DocumentID="gimp:docid:gimp:af2322b1-529a-4b8a-bb63-8a16a68440cf"
   xmpMM:InstanceID="xmp.iid:e2ccc7bd-7563-4995-8bdd-ee54e5669374"
   xmpMM:OriginalDocumentID="xmp.did:abf57cb8-2880-4205-bc1e-6b7909543b7e"
   GIMP:API="2.0"
   GIMP:Platform="Windows"
   GIMP:TimeStamp="1716065832663280"
   GIMP:Version="2.10.38"
   dc:Format="image/png"
   tiff:Orientation="1"
   xmp:CreatorTool="GIMP 2.10"
   xmp:MetadataDate="2024:05:18T22:57:08+02:00"
   xmp:ModifyDate="2024:05:18T22:57:08+02:00">
   <xmpMM:History>
    <rdf:Seq>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:1c838011-541d-4cc5-97cc-1bb3eecb47b0"
      stEvt:softwareAgent="Gimp 2.10 (Windows)"
      stEvt:when="2024-05-18T22:57:12"/>
    </rdf:Seq>
   </xmpMM:History>
  </rdf:Description>
 </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>B#3A   bKGD � 0 0*�IS   	pHYs    ��~�   tIME�9
�ML#    IDATx���%�u���{�qo>�����DR��Ȱ���O$f�F�Ԁ��'5H�!@�?ȲG�D����w��>"�<�a���EȐH�� c5�]��7�u�Y{-aŊ+�?���ӫq���!�i"�LJ��2&����r~~ngg矾����`]�+V�X�/Y�`Ŋ3�={v�s~r}}�_�zUb�OD��8����)%j)�*!T���K���A��Ӌ��B��������X�bŊ��X��_?��O���Ov���W/_r}}�~��x<��DN	!�@����**��v�����躎���?{�w?�w���?[WvŊ+V�wŊ����Ϯ޼y����n�n��>��ۛ[n�n�#!=x���9�톳�3��-!��C���B��R3g��_\�����;;?������+~-<{��*��d��<M)%J)�쉠�l�[�l6�~���s�bŊ��X�ێ�O�������ӧO���@)'^<Λ�k..�����?��o|�������05'�%WJJ�Z�Ry��%w�;��޻�_\�Y�u�޻�����(���?�J)=�a
!<QիR���	��""�}O�u&"����zj�b�
º+V���x<~g��=���f�����!��~����-/^� ��Ç��^\�|o,��ȹPr��
�f{ƛ�WT)�Z�Z��w�ߋ�?��j��'�����榼|��]��H)���13Bѭ�""�� ��������3���������X��+V����W�_�z����5۳-~�C>��0D��vK���n�n�g�~K�ju��*"��QP�r~q���~�~��p8|����ͧ��ֿ_յo?�?��㻻������憛�a��X0�ηg<|����s����J�i�9g�a`��]������/?��{�����p�ǬX��+V�V���W�^����px|{{���������򒻻;��㑔C�����n6<z��T��M�a!b��Pj� He����+��=���գG�|�ӿ�����������6�v�Ov������8��R050q�v��\�����b�C��vZ �SfG.�/Ǒa�����ɏ���o���maŊ��X��7wwwO���x�ۑs"��n�q8���K~���x���p��������vKL���,`fNpK��7��q<2��4��~���z,�JrW �������'��׏w�1F���9;;�x8r<���00�������K4���[b�Dt]G)��ϟ�՗_!���>�˿�����?����[�b%�+V��M�˗/��ݎ�~Gɉ��7��w�{vww<���~G4%�)|�����J΄�W�Z*Nq]Q�b e������哟��G�޷W��ۊ/������7�}����O�Rk����8r�������%��Çy��������l������M�C�qǉ��k^�|�0<z���׿��O޼|��w��>s+V�wŊ�����{��g�?y����;�4q���������4��R�7=}ߣ�L6�R"��4M���qU���Spr��ЩB)7�<���	�>�?�����_����p��˯���͛7���qs}��r{{C)��n��vG�����25../x��9����]����C>|���9����www�\_���+�a`\\\<~���7/��ɣ��_=�+V�wŊ�I����x�����=~��)�rʨ���c�Ja���G?���"���� Q��\��T�)#!g�<��gg��l��>�ُ�wvv�������|�����~������������kr.t!pW+�0.�yRş&J)dI��a�勗t����K./��l(�p{{���9��Q���������`��y�X��+V�&��gW7�7߽��~���K�q$��;L�\3}�	
B!F�k�"N8TZȾ8������OD��,Oi�&hɼ~�%e:^=��׮��ۏ�����i���kKE�b��{%��4�m�SD��%�S�9SR��LN	B�ݰ�n�϶�Z��|��:_�+�>KG�P��C�{�M�!"H���N3�ץ����ߵUf�.�,"���ȧ����<>}�������׏www�|��4M�@�>�T��z�'"B��0���v`h�"����813�͆��3�_<���t}����Ͼ���k!Ċ+�]�b�o�q��8�z�q�������*�tLQ�s��Z�䄅�U�zj����BKk6j�0��F�x฻���s�<|����./���NP�I�����"!b�T�#�a�T����d���4%�8!��@I�������36�@��c)��aV��\i�Hn�'��rt>W'��;5�/z"��LnK��\\e��u���꺦���_>��?,'�⊺�(�	�������t����33���������n�_?��O~_|E_��nC�bڞ�po�ў)��%�j[�\*9��@n%�=@S���J�� ����}�׾������VwŊ��X���>~�z|���Gw7׌��}�;���x0�ET*R+y��Ƒ��S�z"uԂ��Ȕ��T'�9���6��H0#M9M�G��~	]�K@��m��w��I)q8���t1rqqA�:����6P��s���
���rº�������|K�_�S"uW���>��]\�R�+�uQ����VTOJ,�F��*9%rN'�{�;n�n�=��l�l&��*�x��3�k��.���j���{��\��?���q3���_~�����f��l��j�=+b�)mH��gTd.\�`�����^�����>��W_��O����Stx�쌾�]d*C��E��K�<o�V�91M��R
�41L#�⛵�C`GR.�V1OUx������'��X�zW��Ǜ������'ww�ǻ��n��R�����;�qX��Z3i�G�����;'�3=���fMMM�T!�	�HS.���p<�4_�����B�|{���9�J�@�@.����~��Typ��w=�ѣG<|��"iI�H�F"3S)`��b�`h���[Cp�>�f��������	�z:���Hh��E�m��/9�^��S'���{=��Z}�S"��R2fN���-!vLSbGrNH�t��*���]�P�,*��/��̵��S�����:�4��x{󩚩�͂��7o+�o�S�z��)Ͽ|�͛7Ԝ	���"c��AQ3RΤ��:B��bQ�7>��Ï���y�o�{�6�[�����?�������Σ?����[W��ƪ�X�����U�'������'���Ƿ7��\�+_���80#�q$������z<2��B@C<�9�[�!�L.�	F0�
��Lj6�\����	�L���uE]K-�2�p�㭥2�#i�JEr&�b��\<��:�vK��d�\��d��(SF)����=r�m���º��d�uZ�6���B��"ykSm�,��F�|���Vj�(�����zOMS�խ9�:�sFf�C(ʔ���%7ϴ��SPU����Ϻ�t�/ţ�r9)�3��36�3��ʂ]��[	�Pqo-p<���cww�t� !D��Ȕ\	$(�Պ��FpE��h�<؂Ȗ�0N�S=�Z`�DW�U���y���W<�����|����X��+V�k������4~���������^>��W��������4L�GZQ*����Ԃ�E	ZN
�lL�)`;"�T麞�0LӔ��\�'64���`!.|.v�1�S
J�&?"��_�ӀE'M��o
L���̃��.ϑ���V`�[Dԇ��{}s*�𕓷x~}��OCu���IqmkP�`UTO6�e��N��\�������q���D���K�-��S�hrr��A3L��+eJ�q��\�T�X�L� L5'�q`���4���n�P�ﻞ��xɇ�] �{�b⹵}�Qkel�BP����l�b�I`,�$P�B0B߱�6�,����'#�r<)�c��M�a��w{�
q�y��\��#�Ñ�>�������'���|��JrW�X	�+������8On^��~�7?|�]ݽx���g�oo���2��5�))1���⵨���1!v�}G�������q��oS��@��,BQ��a�"ҔOCMQ;)��������Pճ��R
A��F�
�����@���=���E�׈�)�A����`�;Rʐ���Ŝ�G�������{���]��O�f'�*S��q��!f��dQ�k�G�ſVU�P�B��j���T��>Ab@jX�aF��,����R���Wl�JΉ�2�0����w�=ǻ�q�ljYQ�1Z �T+)O��mD�Ԃ��o�X� �����#eڀ(��X�i�3D�`\<z�ˇ@�Pc�Ӂ)M��N��b@��\���Z�tǮCM)r����nON�Ϟ��������ܾ��O.�]c�V�X	�+�U���������;Ͽ���au��%7o^0�n��H>�OG�s���ZFT����ɤ(��t�۞�f��I�00�9�`�S�x�@4��)S.�D�"�17mS�g���Ѵy��Vt�<K��D����x�XJ�:�8�n;��w>���N�B��^��|m֣u�a����X��|�L�^�����Ikk[sf�nQ��A�e��Tܓ;ǜU�Y��2Z���u�H)�rRr���^-RHŽ�%gJ
�T��u����ǈHe8d����������׌�e	97;Dm$��f�X	�E��BM���o��'"d*)�Li m�~�<1�wT���R�)A��8#��H�!T�RJ&%���9M$QD|-�t=bڼ���H�H)p|p�?p����/�`��o>>�n�l�+V��bŊi��۟\���|�����hw{{������/��~I��h)lcG��Gӹ`�.ܬ]t1RTɪH.h�7u�tt�����u#���'� �g�tho-��)�)eR�H9��g-a`���K�,�i�6X����'Т�r��H�HJ9��^���wy����؞]6[��Ps�ֲ�K~oS���2�r�uʜ1Sn9E�Յ�*R� �m�Y����o�EϪ͛���X�D��}�f���\m�Wy�R1qB[0��5��Vb͐2���p}���+��פ��9e�V���$�T0q��]|#| ��K�0Mdq�;S�f�40���ra,��xd�P
��#)�!FO��l���`��B�<&FPT�S1�6D��Ml6g����%��9LǑ�펠ᣯ~��O�[�^�
+V�wŊ��x��gWw���y����non��}�9�/]��ӑK36g��c@Ku�)�G�3�`��������3�3#l:�>��UdP�Q�9���p�B�-I ��Z���8�ۤA���P���V �fO�mٲ�j���i�PM�%���8�v�Á�����ѣw�x�q{F�o����RO��9�v�Q�O;efڢN6O���@1'K�5E��F��P��K)u&��~Ѡ���Ȥ�l�uIi���`���W�n��Z<��bѰh�>ej���Ȱ;p|s���k��_1�޺2k��B�M�`��e�L�`Ė۫�
�0M��J!����y��8M���T
S��O��+s�x<���ns@�ȹ�Rb:O����%�A���F������ggg�]Oґ�p�ͫW������'�?������W��b�o֘�+�-��?������Wϟ?~���~����@�Wa����imC]�Q��?��O%�JY��ɘ�Vr-hľ#�*���8��Z*�z�XN�M��Q�� (�����q}{C��������S+��g����V�6�Z��5>��Z<�5��Y��J;�/.�|�ۋ6ggl�h1[��z�B#�����60GOI�u��{.[m��sɃ�S�[�ٵc}�zΞ�:�z���� [��.Cz�j.�`Bl*.8�k	y������P�����_�aws�ݛ����f�-�ZK��Fqy+��3gc�0B�����ke�cNL��=3�%��qL�)qH�!%F�3�)	(�h0B�������������zT͟��&�-�X�l6��_pqq�����GJl7[�����{�_\�`{~��������6��X��+V���W������擗O�>���~�����RبҩЫ���SSngնQ�{D`L���eh0j#�S�L��RSuB�rE�a��B����+�SΤ���H*�c�����nwGS,Tm)��F�=��3sg-W[t��!4T�03S���+��PS�;r��·f��l��؞oٞm�b�>d��.FB�r���*��,�?SkŽ���%X�B ��3mA������昮h��,{DW�l��j@p;E)�km�v�E�y���{p�ib��i�vR
�q�۱���p���������vL�#Q�ؔ[3E���UN��چ�D��a�;����Aʮ�N%{B��7��S��X� ��p&���1%F*I�$�$Np%(b�@ՇC`�&J*���q�=�kf)�b<'Z�RI9#��}�v{�E+���m1���wx���|��u6���?�_�hUsW��7�բ�bſb�>{~u��~��������~��&r�EzS��B�bRQ�
����x��uѷ�c���l&��EĴܼ�k$ X������
�7	s�V�C�RJ"�%M>�����u�h#���"ˑ�p��5���9P���.`-���:�����g#ǋ���������@:L�=�lB$����Eb���!�͆�m�&Ĩ���\juK�R��W�.�w������cԚ�a)T0���u/n�Й��)MA��d��u)���A��ٸ5�0����iH���n��n����Ȱ?PR��[�b�jfk6�5�I�Q̇ *�T C��ŝ.��M������7ѹ D���7��A��5Ω�'�?�{���7��8:�7n�)OqPo�˕�p$G�݁�fC�^ ��8v�=g�.�^\>�7�����o�۞m��{�����X��+V��DM�I���i�GK�7.7[6A!'j� y���*�NĈ��������S�b�%�=SI��Wg�ch*�S͒�Lθϴj��R�40��fbP�)�T3�
4��
��y��D�ΐmg�A#�,*\�uSjr�;+}�tc䚩ZZmmb�Ry���
�#n:���3r�Ġ�`8yW�ѱP�*�� 	���c�,��&��BpK�X)TQ��HnKt��K$j���1_��Mr�L�@F�7ܼ~��掻�w;��4NH�!A�J�u>��z��l�[ETZ���Gv��:���y9%P��m�:ٙ����U �6�q�(l��\Z�n.��A�k��2��)3����r#�m=�:�;��՜�{L���ݎ��[������GW9MW^�ן�����������+V�wŊ���9g˙-�NߣQ�v�i��B��wXS^���B�#g]h����̶�;�4y~t����֎H���0>%;ζ[��M��`f��VW�,�,!�D��)%�)1Gj΋�W�kfK��������=ES�x]�ez��Ơ�t!����,'-�И	>4u�{��]�e��L�)O�cA��g�qv~���%�f��5bt�W��AP(�s�G�2���	]h���zxA���� h.Ly��޹]�)ݳwJɽ�SˆM��O#��;�޼fw}��k�05�.��ڲ�s��$I�o�\�ۼ�U<!S���|bp��8Q���kO\B��.��	�3(Bh�}��(dQ�*C)L�8Y.����
�8��Sr�4�v���j~��j�8�)��F[	����T{7/�~�|����v�ݿ�?���}�����7V5wŊ��X���˙�VW>K@�Y	
�fJ5�ؚԩ���ɬ�->VW`sNX��#:tn�2W6+��{ζg��P����:Kv�E-L�0�BN�R�:��� ����KAL���y`�L�Vu+si���WL��������U�bè@��^Z�kgn��@N�x�l��
*�8��up��0����Ͷ���ͦ�[�� 'Kf�t��2��%dUR�13R6��^Z)J!My��%�@Y-�ó��%�v�#�ƣ��    IDAT80�����Aj%G4':λԚWو�j{��6� �b1�P:�\���\��U
cI���5�t	��XPD"���c���Q`�R3X���Qh��-�C���Ua�ڨ��b*KS^��հ��ڽ����~����Ip�����P��JN���n��/��\�������j��z������`UsW�X	�+�)�S��	)���;�j��m�G=wS�������;�U\��a���ء!�8�Yiu�q�o�]�Wk����Ք�L%#goɚ?r5��.�e-OU H�7�K0��,�bc�P������1�������y�*�"�PC:W�K j�tE	�I���MX�4 9H�PJ���[�B ���F�}+zh�V�ק%��%����2P7�.Myft!4,�q�ל&JNh����}�/��_���?��m*�fC�+�a:P*Q� ��L涹�^<��-)ZÚܕ9���HCE��s���@D�蹖.L�C��J�<%L񶶜ȓ��\K+�p�U\�W%�yp��)A.�)�LM�%>���qU��L�C������ݞ�"��k�R{�?�����Ǳ�?�~��O�����X��+V��(�=�������"m����Љ+�fޚ��ٷz�I�s.Vb�0�TQ'Q%���7=A�4M�44����e���Km6B����:����T���`���6eA=�e���USm�9�u�G���!<��Itm~�l�=�R�҈t=�F���9a��R�QcJ���j��⥊�T2�z����ܞe�t������*�.�Ҽ�]�]���i8��()!���7�9�����\K��Y74�5R$0`l1vE���N�(J�S�j�{m�!����,���$DY�H:b��ٽ�%��7�[!��ڠ�v��^�2��[|�Kb�_����ob�����){�ok�+)QBX��L��!�)sR�9N�FD��-*�,�J�ʔ
y�'�|��۳��1Ƶ�lŊ��X�⟤��D��)J��S"��$ּ��"�,F����Y��Jˬ��Z�$`��hC���D �!4��j|=
�I�'��rW�b%c�`qBS��Ҽ4y�)!x��
ڻ��B�4���KZ��#��������a�.���'�rUկ��b%�a;W\ݴю�����в���D� _��9[6)��ښ���L(��ה���������3uar�km�3�H��!���Ä6r�m͚ϴ���cm� o-b-��}M͙<�H�D3B{6�q)�y�gB��ª��W�q}��>�םmy��1F�vw���1f�R ���Vs�}v�
R������i�BD��ˇ��2SZ�r�	J�.���t斜�ho>��g5W�]k0d��KYN �U��Ԃ�ǁ�Ϟry��.���������p%�+V�wŊ���[]�RS"�	�b�f�T�������.��䅤Ѽ�RY��4	��ڱm���C �	,,��K\���fIަU��������'�Ee3��j`�����W�zZP��3��+�i536]G�w>u?M3�q�ܼf���܈V[�@i��jB�@$������Y͵f��	S��u�:+��C��Ɓ�єx~Fh�/# ��`K�kM�)��d-�A/����{�����U�[[/��h�]���d�����	s��[jSciy���]S&��jh׳�l9�n�bGJw77Ԝ��nW�
�~C�o�@�i�T2�z��0�*���Z[���%͒�-g̷Cj�V�4R+���S�	��y�٣�Z�C���d�����m̀�ݎg_~�{�wu~v�dUqW�X	�+~]x׫���ג�"UZ*W�B>Q^gB�$�+�W���@0/\����g��z���n������Z������)��Q��sf��S.K�k��D����+��l�9.��UJX|ħ��爛c��:Wю�է��=#Hi�
9���F\��y(����joɖ�늮�[�X�ҙ����]"g��:����=�8Ş2��-yI3�Ƒq�<Y��H��E�[C]m�l�ng��|���e�+$�B��C�%I;��K.� �P���
�R3A�FG犲*���UcQ�ؓrf<r�Hu���7��~ՌHi�����bٕ|k�SjEr�����Gkys���ZI%-�,͎��PA)d�,���b����R��:V��Pre��~���N+V�wŊ�/�_7o�L��1ÉU��j;�6�y,)K��+�A��rL+��U�b������.ت4�Xۿ�]�)1M���O�5��RI�D�G��HŽ�f���PDH9�o�z��L��X�۳\�]���G^�d �M�M�vr�o)� E��}�lS�#Uka�`��5W�g�TNW�%�%f�/�ǖ� (]�
w�׵�ku;�~㛕Fʆa�0���ڴC�ao�4�����T�|���-�҂t�A�Q��0��`��P'�45B���[.��!������D/գ�B�S�i�xؓǑR��;D�I�~��}����NpYr�U�bM-�6�V��#���LɉZ��+3���B̟ǂ��/��br�X���S���j�E���N�ˮ�{4���5������?�<\+}W�X	�+~%�R��ٕ��11/P����X@�,�驴�R9M�������L�m(�N^N��k��'iCiMhmk�c��		Z�P���>)5\���k�J��"�{�mh���2���D����s�A�I
�r�����j�ւ��R��Ii���L���!�k��Zs�.�2{l�-A�.Fb�˽�R�1<!Bnf!F���r��0�j�;ے�L�����ZS��kK㱩̺x[��ՖDP��[4FB�U���H�^�Ԋ�@���)�w��U��Cy&�rjy�SKKhQa"�m6~���Q����#O��t�mG�
���a������C~S�3��֟��t���4N B�b;I��vE(RQ-�%O�3�i$�dJQ����^_[aEɉ��-�8\ݼ�^m
+V�wŊ�*j�>�J��VϿ����6rٔ��K�'&��ԅІ�B�oDKq��9"jΐ��[���z"l�0PN�	�):�t5"8ZMid��:%�r¦��.�yhD�{TZ�Z�so-~��	ʬ��lTͤZ�h��Va�dU�drM��?�T�
"�ѵ�slːS�/�,$*9��7�=��B�F��=���1nч�H	����8pmȫ����.�ŊPL�mh�4���Z�[)N K�e��AR��V�����Gƒ����fC���և�&�0���l��hrb���i��<��B_������_��x���L)����5�]O(�~��~ϔ�u��ؤ�8y�j�<�a��\f�wh��������C۰4?�\,mC�a�ŨWIPR�x8p����զ�b�JpW�X�k0\Z��t�j���v�<mǪZ�/��Q��.Wo���$)h#�,�R����ߥV� =k>W˅l~�^sr��J#9m +B�Ь�d$M�"i��,����u�
�{y���������b�jI�y"⹳��d�)	)O��k\��p/K�4Xik'���h�T�sMnJ��ul7[���y�mo�	���QK��WQ��7�fJ+R��LJe���ٜ��P]Τ���v��w�8xC��~���T���t��!��~K/�]\4K@q+IJL�HΓ+��#Z$Ği��)Mng�{6}��^0����ش�+�hϡ��;����E�r��?#�E� &��A������ꚳ�Et��?F"s!Gk͓��k~rAS����Ư�Ǖ���U�� 81�On�?����gUqW�X	�+���{����6�[�5��j�*'�<6��_Bø�guO��	�/����1`��ȭP�Q�g��܈լfs����Յ4䜑v�,��a�!�K��kk�櫝�reQ�KjG�!x>�8�K:@m�w���;WѶ�>L7�Omʯ���j��M�JJ�^4��>�G��}�����$�ɱ�Oy��2JK��R��Dijqm6���g!��&D�~���ٱj��ĵ�AjK(�)��DL��l�Z�@i�i��G���p$O�+���҆���d9�ŞM��6=��S�0��L%���;�6ol�޲���nS�0Nt}O��֔y�-4�.7��8y6pN��mXि
"s�3�Z��G��)B�ԇ��*}��qON�����4��MaŊ��X��W���y5�Kn~|ZsiǴm�J�k{�UBk�j�ڹJ��k|���BO\�I����="<���*��r�y�A��4v^g[J��I�6�yV^UѠ��&�T\5?�֦�*,ʮ�?T�G��\�ǱY�3s�ZK0��dJK����y|_��پ��/��Q禲��KFMZQ¼�~}K�F�a��D]5�g�h�v��h��7R�{�81��+���@�X�l�[B�^�1+�f����yNRi_���)&3;4:9�\�Ld�(fH׳I��x`��3J��o��li�����,�d�D�U�t#P5�P�
Y�b�&b��[�qf����Ԣ�愄��\oH����s�"�{���?g������*-Y�T)�`�p82��ÐןT+V�wŊ����yp`[Tܗ��U�'hk�b!c�;��RYF�OUM�lN����}E��}W鉡"��j%5�k�R�H9�'5�+T����X,�Z�9�80o�reM�<�E�Aj+>��Xi�sɃ�,𵤐�����NCgs�U��_���#Į��ч�R����gJ���\�U����Z�1{߈Ӧ|��ʉR�^p�����H���g0�g[�-æ'�¦���ly����	�EtJmٯ}���W���o�Z�8ϛ�}�;���:L�!D�Ñ�+:J,�1ve53'������Jr����V��,WWY�*1$t�r�r�t�#��8�%�L:%����6��x�O��l��E���AGiCws�R6LŇ�a ����jŊ��X��W�6Z+���Y]���s�T��"B+#]�^cllۊh�s��O]�l���-R�����db!��X�RH�l@kCBTO1Г�V��մLT��mC@&�)͂@#�U�����be��	���hf�O
��+{�	�L�U�ERy����J\ke��H�:΁��N����Y,!Z�nMh�a��%W�l)�s]ot���y�V���gg>�W�_�E��-�sgSM�9 ����]h�2���PV=Q`N�P����b�=����fd�o�����J&�@1a,��xd��	Qz��!b�`퐢���Xt_�)��}�b�d�B�H�5��l*B������!�?a�N�����{�F���-⛢a���X��+V�j����J�ꢶ��J�m�	�d��ĕS��}��w��ZO����;KW~��-`�\�o�xZg���ʚҧ�CH+O�+xEN
휔���6QI�}U�J�7|6���4vo0�NĘV�,����Z3�_��[u��l	�=ͭf��6�{r)���?J�����M��Y/o���B�U܋�B�B)S#��յ�(��f�i"M���������+�!zD[N������7���!P�ZHuW��K������M��,�V�Z�Z`��rv~��͆<��[əq��,���U�ɽé��ڽ1i�x������#g-�LQ�id��Q�M.XX|�:�0�p�*��=�=AN��D�	�VQ=7$��8N�)��'Պ+�]�bů �ZD �@в�a뜚���gͦ��<��quEoQ���V�����,�.ٸ��H��2L�fX�WQ�4����(���i���}\��ܗ����5�ڈ��T�Z��7���mUɾ�-9���Ui'u�4��\��H��{$V��{ʲ�(J�%�����T���V��+�u�y�`G/+���	3U�
�O�Hj9�AB ���)M�:T4�*9O���U���n�[�6@j��) ���z��͡\rO�o��s��*&J������p���x RNX��<ac Ke��E�-�6[��Xi1i̻��\5B#��g*����ɷ���^Njmٸ,>��*rO��噞��gl���B���#O������w~��ي+�]�b�?���WW�pxR�#!�Vd�$xi�Z�a������}�<[b��o��5��=dj��`(�4��E!t����㢢J�֪�sS�����,V�.�L�9��.��"lmA�\�_����RZ�Ui��>�7?���a������Wֶ�����b�y	�D�2�$�W�Z���G5���4��u.��u�ڨ[e���zC�����[��E�vt�#�2�"f�J52c��l����s4��jU��eB��r���^�����ZrSA�Ek5�-61,g�ؓ���xS��.z�]�����fq�6��*��r� j��/���u#��(�T
!{�C��Y\�\��W�%����-��-�=;�Jk�-�͐
1F�P�^��$�+V��bŊ$��z��&דt��W5$4�U�tiƃ�[�2{:O�v&2�fj#�������YYW�m(��@����y:������W]gDm�������l`Qcg�l.�p{��rp��.J[�۩�)׶�v���-���'�;{�����~��clQ�D�@[�c�]���	U��Ŝ+�&,\.�Qpm3P��@d9b��km~U�*�Z)s��!FĚ���������8iT����[Q��d���#y�.�.)@��������R��oQj�\�q�dg�Ur#��F�^T���W|�������l�8����%�7ϟ|-����55�T���y��^�򜕺T,��l�bŊ��X��@-��G�R��m�	����6Ϗ���S�����S3o�8H��b
�ŋ�o;�{kp����|"}��{$s�S��V� ޠ��K�OQ�{G�o��
�J���n��Y��R\Jm�K����P���Eu!,�a&6��iN<�kή����!-B*Xp����^�z�6���+�g����F��{�%ɒ�HS�9Yl�#�3�C���S�fD�{?++��+#�� �̣���{mh������=j�O]{8�j�F#ZEP�R�Q|�'p>p>N<oA$��ե���pU����z�M�q�u�*��E�;������ta	Ό���%�1Ay[&��`�]%2�wi�S��Z�Ѣv�3r�ψi �e�ط�|�G"���o�0UeFS\��(�سg��{����1�����UC�:�� 
���5�QO�ͧ3Z:xpo��ᮅ-v��%����p�aZ�@Q����WduS�3��i�=8$�+��i!)�Ru��E!�����F��X�͂ukÎ#2�E(�/�Kֲ*V���1>���X���*˙G�+���b]��,��x6�J#�������b�,F���K;G;.�D".��(*NW~���MD$õL�9��t}�8?�^t+�7/����7<,�S˨�C!�1�'���L���g^E~c!�1CZC�7��Gi�!�Mb�/.��Ѭ�%ꂥhM��Oׅ�*3� Cf]�g*�a�ѯ;~l�=[��ٳ���#!̢���;�� E.a��/�k��)vW���־���8ψ.x�ASR��g��ٵ����q_O��ʬbGCCk2[��e䑽����U� x.��v���85��^[�Q�)�G��m��Z��( �����:¦�����m}!�������!���Ŋ@AD�b�~O�gs��Q���������M��o��l��D��S-ѥhg@�9��� ����jW�)R��#�ñ�n8���Q,�y�긵x�Ikc����#��2��Z:K��Z֬EF=�ii<��pSh���C�n�=[��ٳ�	\$d>@5�u߸��p�DH��u$��Y�k��Y�9���4���cJG/��Ł%��� EC��U�lR�B5��2��{;�SR.\���p[��=	�F�G��?��=]N����4Z��t�X_ID�B��Z5�m��ZT&{!��|A�U��K�1���|}G�:h���}M!,ɀ �wO��li��8s��h)#�|�9�+3���8ζT��QQ�#o@ɔ5�8=^��d#��e��A,`qt�ѓ�{k���4�	B
j�� �Œ��H�y8���j    IDATK䷣ef�aK|�y��/&��g��.���P���wR&�;���������?�׽h�g��{����
w��z������in	�r6��e�����K	��rΆ�]��'���< 2
�,xѐ�C�
�t,ty��R,D��V��>�*f�&���ю��5s��P�p؎��m��J"RT�C���G�31j�tV?W�,��MuY:kAHg�K�&d�����6�l��B;Db<����)0M�'��[�0R�Z]p��G�2���'B˱�u�j�r�,# ���H��������cq�ȇMd�*�)��bb�0^r��[�aȦ�ڇ	G6�	@,��\�S�HpzWʆ�c�˅�Og���{�^�塡p�hM��7IaϞ-p�����������"b��%�*�S���M��R�Q�+u$�h�`o���pY�B}��q\�
���[`�R�*��A��#�x\%�Z<R)�3D�v���Z��⾌�z�qtnDWX�/e��Ųز����9ۤ>�}JJP����3e�yq��.z��}HǜrI����xH��_v���<�(Ԑ�5��3 2wI�?/D���>��hrdA0Na�,�0IȢ��
#0�)���J�3��6"@ �Í�Lf��.���9X���sfB��#c-�"�@�����E��H 6��xj��k|�\(K E���)B�ǒ��I
{�l��gϞ�5p����ۉ�� ��P8dp�&����k��_�>�D��y.#�h̬g�κ�>��L��q��I8�P�_���+�8#
�����XUS��C�³x�8��h�����%�Q��'O��	^�"#`����E3VrQ�)ټ��'{x�iL�B��e����J�k�A2\s���!����f�2�b������{�u�e���g�8�u��6������@-3�ZG��$D;�)Ў�I@���3���e�!6�:!������J�d��)��Pq�{�*6AcYl���\�r6�-�^����( Y/���ٳ�={~G��Ir�<�`�Y�jds�/m�to�s:��fh�?W��/�Z��T X�E�$�?��q4@��+��,�N��C��h.ʃϪޅQ䂪�6�۫���s���2'�MB0��~�q�f8�k&�P6���ة+��C�Չ��48��f1�Q�����/*~��:P�n9d���Y�G��7�r�K��ā�ۅ�12ܼd���<�^��K[�P�o��v�@e�UG�  #�4*|��})� ���W�-�x�$5I� LЈs�+���h�J����03מ�{���wϞ=@�2"��<���u��v�����ʙ��c�� A2b8qO�ϻ���42��
��ђeV�3C�7$�O�SL	>���Z)�
�Up�*�`d�����ʥxf'8��=�L��V���\��dm�y��5����^�j�����̎B��@ �)�Wr���O�B��P����<ٹ��o5�����w#-,a�B}qo��k>.���WT��@CW��Fm�eC��2+�׍n}|�����}��}"_'gn��aIy�!/|��:xu��n�IK��e]��[��ٳ�={������ga9
��s"p,�����4��D3�?�}ɦ��.��n�0�o�U.����������'�u�:�]"�S����uFrO#c%Hb�pג��5D�W�;����8�Ξ}k?��w!�r�<��>5�c�>�4����q>��,B(�5���.�R��>��F�FFC^r��m9G9�����:z-�ЫĬ��rOq���r-��리�����r�� q�`�\���J༢p����&�s�m��P
\׈�H�|^8Mm�A,ܥ�n��vp.��xNP�_&[��{V���by�.����pȱ�F�Я����GkϞ-p����{���5��n�z�o�LyLl�"w8lyd<���L X����M��Žu�4�zG)o�/\�O������V�B������Ɯф���E.�#oOz���Y ��������oo8� Bp�Dz�'�����]G��~���?��h��x<��q@��"�����}��J������E�c]���)�缎�G�6o���>.�e�ϯ7��ݗ;�׊��ʥl�"�s��dq��� ���:�b尤uDλ�`��v��O�!,p��@6/0d\���/S%.��gV��!��i,b���Nn�1ˈ�>�kiq��s�����s�={��ݳg��;���
����J�E�DKޑ^�p	px*�����xU[Z�k�`�@�ƂUqo����N���}�g�4��Y3�"�'����g�����?>��sT�u����u=A8�U�z_�p��$�j		�h3>q���x�W|m ��03�1�����,Z���4Y��U	ĒI^�X*s�#�����)����[��j��1Enx)7��	w|b�x�Ό��"ri9�O��C��� �Y1L�r)^��[9�"`IZ	{^�iYQ�Z�>nk,��>?�(���v(��. �{<�?��J&����[�q�4�5B�����ٞ=[��ٳ�\�W�-)@)��s�i��ୌ��}�Q(���u�\b��)�KN/w�)Gځ�pa����_���!�G;؟�C���dE�Fk�p��V����x�dh︮'�������F����� ��p.(5���o�[n�*o�JD��く8�s
��%/�[u���t�x�o�&�"Ć��+,�e#9��+����#wy�d)��Hg��I�(�r9U�)D!���Ʊ�q��,D�� 4k�`�t�1\�r^�|0�}8�!x�M�MlR��#Qu��#�3��y
a2���1E>�d�1���b�C�l���ٳ�={~o�/K���oջ�uA�'��G�)kj�
'�.�u��U8d6�<󩿡',t���Z��@��p}ۅ��� D����8�!��G�q ��э�륖U����_KW8���l�4&"�U�����0Ka�8��jf�9��8*��ځ�P���8�D<��"<���g`�~u�i)�X�	���!�ц��)i4���[IZ��`���&-0a��B�Ƒ�s^x0���`O��Vl����R�G�-�^<����ӲN��pd�#0k�\'�`�����.F�����sTX7�c�7a/���2�Ů�H�?�3'<���^����Wꅙ�=�������?�����]��g��{����
ׇ�'��U���7�_��F> �$�ح7NVj;�B��I�m�̓ze6�h㞬�O���q�H�`3p���)!T33<����C$��iҷ�[�����t=��t�.�0�,4X�NN2��\�,Ե����w|����`����,X ��kqy_�j(�mFJc)$��ڇSI�}$$�u�!gS����[�#t�Ak��J��]ZB�y/�'6�$�*s1�_fI��C{�w��U`�X	s-� .��2`w�v2���,�H����;�5/2h���ǿf�G��\\�SQ�����K!
�u��D!�K�Q	��������wϞ=s�^jwkpG��"����77����J�7��I6��B��AG.��.�x�_f_�\/���q���}� �<ӄ���Jw͜j@����B�bP�R��џ��"C���@K�+"���\�F3��\��a)��цk'ٖ&�zV�b@��?s��7�l���}����<�^?��<,}{��&�p=�e\�TĚ��	h^���G��/�̓Q�w�"�fyQQU�05����#nA2�����"h`h�H�[���x�yA������D�e���3�� 2+��U�\z�qG9	-����b���ٳ�={����h/[�rD�Y9��Kp�ϣe�l�(S���CG�@�GƆ*&(�Ռ9���EhXH�8���<����|מ����N��:� -���p��ϟ�׍�xD�����3�S�kj
U��fF�����|s��tp�50�Q�j!k,G�pVg>u�]��;�~��e��ʔ�o�٭\D��0��E��^�����	^,Յ��n�����+
³��������TE��tz3;k���G�6�g]#���W��߷�l�x����é�����8�(np����;�k�q$k�ͧ��V��h�g��{����������A-0!��L�B,�.e.�DA)���\m���,��X�a|��!�^|I�E�m<H����L�rk�*0`%.��e��"	Я�ϟx�����p�nh�cl���p
q}��1��{M̔;�&kVUq���afM�d#��5����4y}VFC��>�ҕί���sQx@��{�ۤ�+ �a�,|ǵ�����4�AX����wU�����ģ�A�F��sF*ƒ��R�WH#CQ��� �=�;<i!�j	�n�ҪVU�~C��Mf�Ge�Ix�>���A����|F���������rϞ=[��ٳ�w��䋺�?3����\� ��M��'���j�%�t�2* j�;��2�����8�q���	��h5[�f�!�<T\��H����2��Jp5<�ğ������af8�$�l K,�,�5���,}M��1���:��8�M����Bt �XhjGdH-%�u��>]R"� �$����`+A_5�<�W�n�!�|�<X�>\�E�y���BqY&�L'2�kC��1�,�R��_z�=.����x�p�л����ڈ�B�=�g�cQ�2_��-S�\v��֍��i���c�w�7�u^$�|l�ߛ�����mϞ=[��ٳ篈���wb��+�����;��@����o�LG�4QY��5���:�1��ଟ�Q&0���q~��le:�Wڳ�aiƪc�r�8�͡���`���|���gf�Ȩ�W���\K�Gɖ:�GL��P@�_f��p�S�
3܁���nK� �E���A�k�yD�-h��,�b�C�YW@-�ǎ��y&��2j�[�Xs�����;�~��P�e��.4V7q�׋�'��b�Ԑ0A���\O��q~�8���g���Zf
� $�{ܲ����4��������Y$�=IK�F�W�b=Y���J��d����7wϞ-p�������o�F�T�q3O;�A����?�����a���S�1AQ
�̭}��깍��^�\�\��A2�@�0�;��C� �s_g!�-.%!K$�A���k`�ˈtU��Sǹ�̑��{׆v�,�X1�����[�O��:���0�8��q.�=��%�!��>�G�V�GT$��$�s
����^wR-��Gf~a�PG S0
*n0	������{��w�y���kAᛸ�b���b�ދL3�"e�r-��"pO�&��%��q��CM3�0��-Q��v>qe_ᚗ�>�� ���m�,�I[�K��Fn�^���fTdϞ=[��ٳ�i���?�	�����/	���ܓ�[J���@yA�@ ��A��__�_ϱPŏ3�s��+�U�O��Dч��n��(E�%�YHP�Q�KKL�u�R�f�lA�[;������7|���ֆ���?>�Z�E2�}w��A,h�`�h癍V!�z�!n�Q-�@�5|T���p=�x>�qaP�m-n����z����v�m8�Q��o������n��;�G�K"?E��7�w��R�Q��^շ�l�����qܯ���zXt:�PTW\�ˌ(4΋�y�0�kBX8��1Zɘ�P��X��I���"G�]��Q���S�z�0� k����%�=�G��TcR&���tj$v/�r���)�ٳ�={~_�������dc��D��j"˨
���;�g�:���`�����p4��Zh��	�*����Tk.K!�����lD��5�<f/�X�����*qk.8ؽ��������"��� KC�'��A <����	�DZ�~�c��O�7pqU{���}�X���w�̌ϯO<������;]���&VX1��v�Q��X ����ы���d�	�l��*
}�����V����Y���Я���'�88�AɈ]Qp�΋��8p�WW+��g�Jc��7B��D�1Q�nTi��hp\E1G��P�by��t�W\[.�͚��P��1��_��z�w�HD���r.��l��g��{����WǦ�8F}e����̀����7�{�v,p�y[f�u�l,o-!h9z�`��f�^��U5��T2�JN g��{Օ����������[5�p��������#E��y�]��b<<��`|~=ѵ�Ue���%�
�z^x~~���Y��������5��M��z��n�Ì掼�J���fea)��3s[��v��ֆ˼�;��%��F���YA���Ⓕ9�y�~>��_EWC;��;�d�j�03��J<�/�l��(��Q��*�q;�qd)H擳���N|\�gS�ӞV�%�R����\�v���5�U�3v02;�2�G��A�(�D�%�]-�A�����ٳg��{���K3�����+��-�DB����]SJ^ɄA�B���5jM�8 Pkp�e'�Ǐi�k(��4�n��jFl���=�fK��{8���=%���qF�{�����	�������'�[�GN�`�3C�g�tQ8��n���}+
 D����h���8�$��9qX�w<����p3��p�_w����3R��IZ�1�e����_Z�u�Q.�n��6�=3[���/���W���g��������s	�,���v>ΈRTc����-]K�%,b4M��Ń���d�(^��%/t��q��^�ͽ��(q��3G</0<O��-VÊ�]OH���b����ߞ={��ݳg���["8O�\�b�}���jAK����p����#� ��0�3\$�� � ����^�"��-�/���M~�,��K�Ki�E(�+��P�R/�1���"���pk�k/8>?}^�׍��x{;�$���S8t J�k!��r�u������	�p�= "8[��X"�a]���u@-��р��!h�*���E�x}�"�4ْ%��t-�PK�o�aݡ]�Z.�G�I�Q�Dv��e����}C����_����3����*��	�d�|��8
�)�t�<+{��!Z���d�YM��D����2"(v-�{�h�����h4���kQ�ʴ�,����3��V<O����ۼݳg�={���yM��X��h ����b�Z�%|؃" �8�wa�I_3�@k 9 j�����-�_X�e�Vxfn7��`;��ײZ�\�����B7��'~LZ��8a������'�??q����i�x>��T!?��������Nm޷��p�w�fi����x��eRX@��|�a&Bkr�0��hA�����M��Z=�>#��r����5Fd��+�D�v�r�Y�#P�W��ݪ�+_BoPkh������1�?N����`C#�B�#�	���-� ���[�8�҄���g{�=n"��<�`��I�v�@'��@n,�BZ�7��U��� OM��j�G��1h)s�F�h�����ٳ�={�����U��|�Y�AR(%DA�@�, ���j8IQ�CHq���c��������j7�\kP ��m�H��%�Bn��׬j֮��]o��=���}=���7���<�	��/�������|||����� ��������F�F�A�y�y�|{$f���X8C�/o'��*6]>J�kn{6����M+"y1��<���P�?���mq�5];z�`D�� T���q���󑤅���:���㎺渓��w�g��ZA�Q�z��w/@�3z�qD��*�h/�o/�ֺ��B��$��9���9HJC��U�[� ��r��S��^��h
�]Lw�^H{���wϞ=i̅Vg��M�N: !!��B��	?�e�}TN��$-~-w�j�H[X��$����n�� Eu�^!��=g�    IDAT��G�fRɄ���������w\�?�����}���_?����_����x��_�˟~�ۏ�Rt�;ބp<�DM��Q������>aB��7��R��r\���}A��NK�GW!�GQ���I���6�l�M� !ގ��=���6Dݨ����F�!�x|�
S���Z�/5����7`����M������G��ęA(�̠0�[�ٕQ�z�/]U�k��<KDx,��{�h��x���e�h�Y^��D��y��-��ٖ��u^��ٳg�={��ա����?�Z�Z��j�b�*�q4�9k��($�V-SIB��ȇH�)}9^�\l�0$�!�"��[�-pz:a0�8B,=��U�.d����j���I-�W�-ך���~�8X��_������~�����_��_~��'H�tC}�\��m��j_xpkI"��8����c��ج�uz �8]����.ԥ#�p#���\ T�d�R�ۨV�nc��#���ᮞr@�#��wk��'���s��`X\t@8�|����p�̭&#�
jmf�ᓉ<.��$�T���ӈ<DqC�6̓����	�d��B�)r�r\~sz9D:�r�2:�54G�Ǫ�d�/�z�գ�Z�1�1�[��={��ݳgϷ���������_�����W9iY�P"e �J�I���a!&�3v���LЅqK�̺[�[yf~}��?'�X\K�q��9]�̍z
\P2n�D�� ���df�G�����Kͯ�ns{���w�����v�����@3��B�}���¾Djp�S)��\��|.�=3��,g���2��
' ^/�f,�� *{M������!����.�zf��т���X�FP4��l���O�n3,i	cɰ^G�!�'�������0&kkM��.8̮ў�1�v0�.դfB���M���=b
���B`'c$\�z�EZ�h�#�g����ˋ�,{X��	S��B� ��ݳg�={����+\����:���FNYÕb֣T!,���qr*��n�/�V�B��D����	SB�ճ�.܌�,~��Y�qu�O맄�Q�༺�h���p����|��| M�����5۲ZK{ɍ�ͧ�T��p��F!������2���_0�!l�i����%�`W�W#ۻ����{�*W�o��i/#"g��X�r�<u��^/�\<x7xO���v;bAa���T�ۘB�w��x�������pp�"`A ��2�R2�.U"��^F�;��b��v8��R�j�v�ф@��Kvo=�|\E&0c��^	����מ=[��ٳ�o��Zp�y�\��>��I�
G7��r�YO�XX���E�2(�[B��r�'�H��4��:�凸-kq�g����r |�|l�e!�p���5���������8'�v�0u��������'=�&�:���׎Y��A�/ܟ_S�Բ�4pk)/��D���
�ƾd��k������`�bAUq=���Ϲ��Z(�����q;����<5g>5۸����bt�u�(��-D�3kq���`�@:�"���]��p�a�K�2�|��E�RP
s���Â���C��u�:�,"9���D�0�&>����r�!�%�Q�񌡃ba������e�˵g��{���[㫕� ��h2:�w���lm[n�3�*�y-���b��t?\�p�k��)s�g~m*�z9�]�0�E,@|��D�]���q�|;����,
  �X�9�BxR2u����;�^"�`�Þ7��~�=G�U׹��}
����Ĝ\[�X3\|fRi�Q+ۚKRϯ/|}}�_$�|Qh��t-.,����G�oy��o�Vw@��է�)���"�j������̌"�#��ȵ����׵$_g3��y�b�3��g̋�Z +���7�xH�(���G����c�COI�m�kB_.$}ppG	K�]a����O�������kϞ-p����..~�b5��*�W�)\"��R
���F�Wm��M�.!ٸX���-�ռn!b�]Bf�[�������LF�`�{�kB,���kǁ�8�^��s�R���ΣAZ:�p�}�2�w(�!��u��z7Xm:xy	a�J#'k�!�8]i���
�X���`�a=����ӽ�o�jA��^�,ed��N>��bPt
DZ6�a���f���yԞ�xk8��d��j��}�F�0������w���z���);�{�V�����/Biߺ9@2������^1� D��4�[��*���& /H�.ua6��|6�a+X:�ٗ�={�l��gϞ�1q�ү=�{IG��H�+�o�kl�'�j��e,��y5��Kza��.g�x�KBėj�%mZ6��F�p��<pb�X��.�4��L�k8nr��-������%��8юZ^��������}��nC�jW��!%2*d�N�]����@]���,)�$hM ��e�ZM��
g��X�ᠵ��p���Daтe�V��рUž$0</2j-1���F'4`���;��aw����o'PH��8-p�������Y&y�� ,��:�2����ظr���@��\|Z�����@��+������Ј��z�`�m�����x��ߊ���Z�۳g��{���ω��SM��ڲx�V���~��j�S>Cv!���nI�y>��=<�z��4��F��q3��������"�K�4�U9L�Q���p� #��v���b.�������#kK��wT�U,�Il�®��ű��_7T{j���H8�,CdQ.��>�>����w��&<�G�й�6�u_pu0kh�0cw︮�5�Ԯ������EnEp$�F.�#{K�툋�t���1) �?��>��0	t�Ԣ���	n~��AZU����Uw�j�u=��
���c�w�T�����j�ˀV������FE/s8Ҫ�"cF��au"1��|�� !,�7��-�f�zG5��yG��hϞ=[��ٳ�w������j�>Bv�����ߑed=Z�T��k]�e
���~��2�"3"��,�R!:`7L�p��iCV��Y4��p1�	��E3+a+ !Ǒ�h
�Ѫh�"��d)�:�����5��z��z^����5˺�ԢvW���8Ѥ�eUr�H�0\PS\�wdF6���"E��x��5`�(�ȸEk�t��a�q��A���McE@.;q��T�Y̠&�;��a��(b;�<b��u���q=��啖"Z�=Dek��=��6c*�XC���
��j���.+q�b�����%�S�{�R��@ϭ�k�--p�;��o�&�m5#(>/"�.�Ó� �Aiϙą���	
{�l��gϞ?*p��]���5��Y쾁�O��32�o�5���t`�..�J�ѬD�G]�D��M4�C
�o�v}A�`��*b 'ǵ{,q��̗���rh�H�(���8:C�	 ���'�G���p]_�3��wG�.�����[��&,Q	{'��?�!�ܦ���<��o�ȸr�k1�RWc��8�h2Ut��zmQ;{��>5�3�Dୡ=c��xG{<���\�b�D9�Ј���[���3o� d	�&Aը����ڥFh�#����~A�>|J�6|��v�83�K��gD<9�>�<8÷U��SA�`
?Vˀ>�<�TG��y:��y��Q��B���#�c-�U�GFk�kK`˥��ƭxH�E�v��*Ǳ	
{�l��gϞ?$q'3k���b�gT�b��Õ!� �=�q������@�t�xކ�󤋋[9ZIS�<�r�ڈ��H!�L�FK���p;W��� �A��:^=�8R��@p���}>��=�_����*ȘǢ��B)P$*m�"a-[���q��G�q�r���e�mUk-]Q�>HrxǆT�5�c량p�;��(� aH��8E-M�qf?]� �u���;Yd���`r_��c:��A��H�w��_2 
~<��d��q�=��zY��m��bb ��DPbh2��U�:N
C5�!���P�	�y,�U耀��b��$�afP�|wO�ޠ����qr~�f��P6�5\_������o�=[��ٳ�wg�ݖ̤�ض�m���b�!��!oo��7@��EwQJ�����E)���2�5�)p��?w�'�kh����}c��n�}@�=٣�B�S���:����X���Y�
�|�w���������q��ϟ��_`�*�Ęl��$���y,?�^�T��3�9!���-����8�<Cgym�X����DV�UႧ����A��+�{f�󂄆��]��y��BF��-��p�5T呍g�G�}]Ac�8Ϫ��@Z��FAT@�!����������a�P�z�k��e�� s�Q@e�3#����%��03�y�L��K�O]�%�m0���7�yu��RŻ�m�=[��ٳ�?��V[�ZF���r�<B���3i�AF�þ��=ĩ��1�8��-YF�j1ͯwi �R
���4:3�=b1ǲ�����7�)��J�88����k�A??��_���y�ޓeʃ��儧+m��5ڱX�*��<�Ú��N���ʹ0W|U,{���30T]e�q<���Y5+�Pb^;�y
�7��`�A�p���T��s�0i�Q���(�XTtDMq��*�����>�ō�'HZ&e��l�=���0�K
�u`��à���>��l���/�n	ܸ �!�׬� /���	���}*XV�L\^:�≙��j�Bo�=[��ٳ�:�i���/��E��ڴ��{�Xɶ^���'����60HR����I ���rt]=���پd%�v�C��`IC��qK����G,G������y�~>aGҒ����B�.�~ǲZ�H�3S
T�8y���V�ثH�z��SnѾ�W6~,��D�_�����U��A��&�����GKg��rH���ݱDJ|�h�����|�E(o��Z9���'�e�q����e�hI ����zw����B��)��j^`���|cϥ;�Lm�#�B>X�47��������種���d�"�%��7��=\��%>JF����A��={��ݳg���]��1�;����2�y:�|�X�E�2�mb�py�b�dGdc{dm���RE�ݫ��X�c�e��Xp��2�[�n�����s8�]a��7���[ѿ��_�� ���P��4�-��ˆ��� ��W��0�շ^�`~�����ؼ�f���I���R��~�x~}汶��3i��� �N�6x��1��u�?���(�W�
���ҶL�u�U���ȶ�F:c�fY�S��d�r:��nh���s�!j}�F5���_�������ٕ�(���V��3�x����Y]���I���H��PEY��z���a�����={�l��gϞ�_��8�� ?jy,�S,���l��\#[I�_4�H�;�)�|��wE��B��pȁ&-��ߝ��-��w��� �C�a%x{ �p���w�E��C�������y��"���hC"���U~u���q�g��:�"��U��^��h�2F��H�ȭ���'���p�'���?�Ym\���4�����p��{d����DΥBJ�=~]���Ơ%p�t-�q�SY���é4 ���=a���m߰�	>G$��D	G���$�҉QE���\���X�qS��]�TS]l̺�QM����c�3>��&Z��-�x^/�;�ϱ�ջgϞ-p����G�DT
�:f.�]��R��0
k�c��,�Z��X�,��N�u��s������;��O<��	y�-l _�<5���������
(3��J�kf}���`�vE������FI@ B��/n�̓�Y���/���������eNsp������eZ�Hc"�Ѳ�+�	�~��*3�*@��){]���8_ �6���qfO�ŮJ!�)n/���B���Fr6��B���H����pf]8c!BQ�kn�>���c�Ыs���N�Lg�Zf���<�` �K�,����T]h���E�N��t�M-��l6�3gm���1��{Q�^�P�{-��CD���������՞=[��ٳ珌�f�����Tמ���Br���7oNU0EhH�X,�#��ǴX�FyX���t�=oܷC����(@�
$����󉯯/8?~���� �����&�@Zԃ9�Ij(l�18�qj���21�`�bZ���{�Ȝ��E.7e1�E�tK-f�&f��㾷��Z2�I-�<�f[�%;_��`��*�V�M��͈��t� 8������aIY�;>_3�rwН�Kio��=?�(�O޳� ��-��Z=옮vf��4���ǎ#�c��
�,�%؃��m,���ۏ�2Z��X����3�=MmL�/��Ōe��'��?������ڳg�={��!�w�1����4�P �S�h���W�K����#P,y6�Q��z2I��p%�9��ь \�������_x>/0�`����������;��O�?~�Ǐ_�_O<�+���^Ā]C��i8/!�"Y0��H���Z,�q!Đ�k8����Z@�x��`�X�+!���^�S�� ���F{If8�*W�4��|P�B��X��ן��@e�IS96.vi#��\���[d�m�1�t�1�d�x�lic���m!(�k� M60$�d�O��Z�`�j
�@�5a8	�;8q�2`NP�J� q $Q�L���(�0��>�<�ж�.�
lg���z 4�š����y���ٳ�={��0�l8wqĭI�l �P�2?۫�W��`�\)�-3�z�(_�o�Y)�NЯ'���K�_���P8��F�o��q�'����x8���7������	�C��3�3�]��啬�%p�S��M��an����(f��9aZ�/ի�D��F`�<�64�s]� ��ا�9J 0�X!����L^��'�fcq��/��lUQ5�C��^"�~M�����1�*n:@�*��������5Qj�~�wfgE$D!�u��4�(��{�ڙ��vh��''^�r���3��:G����in>s��m�Z���&-�D�7�Q�i�(W��y���pY\ߩ�����n�*»�lϞ-p�����-S��i�zo'���gdt�n��ƑtZ��}�:����I&�OXB�!_OU����S/|~}Ắ�
��pa7�4�w��Xp��o�x����vw�� 8��<#C�U��������8���oi��~=὇c��0,ݼ�臲]c4��H����\^#l[3�P��0<c����L�F�!�<3���۟"�EZ���Z`W��	f�k���\���ĉ�{i��?K����8'�1�ӹ���q�qb��6���`�;�n������a�j`�e���z2�#�� R�&�Z;�Ӑ4M7��F�t=��ؑ�5zpj��@�2g,�g	�������&��yP�;��]�����v�ٞ=[��ٳ�?7V������ی!�Hafv�B�5K	�a�N�7>��x^�����p�=��}3ԁ�5���o?�D�q��!o��8ډ�8��������r4���,P�Uю����]{
���6���_�O��q'�ǉ��;�[
��}�����{��9|�uO5����0!�8��Tح�J�nF�A�A���-�b����0�+�P���⶗�j�[ZKN�^|O��=1�b��\ѵ�3�h�c�h'�S�t@��S�і���gJ-��d��t�L��!q�Y83�<�����˥� �e#�z�k�E2]^Nn^ 4�����-����dq�>�[�a�����<ЎcCp���wϞ=tT���^�崖e���Z��B^0X���ޯ8��
7B���*n��鐦hw�f�K��C>��HV�\ADx�ox;Qg�%�J[�q�8�s�Q�1�å5xRbK�E��	&���    IDATn�,���uI1s��G�f�h]jS6��ؔ'4��
S�����D�j��9Z�,�g��W���\�YbPB�_����'��uM�xB�a}�W��w0+�c�OU���+�Ve8W!�5�ˈ��f�Q�7s@5N�5��hD���%M@�81��.�����,Jb�<J'��X�k/^m,��逑�
�<����"i	�e�y!Q
ŀ.���-tϞ-p���󇧫�S�zqX�����l�B��Z�a];����Ԃ[A�8���P;Ў ?�Kம�-�pJÏx�} ��%���X����p�,U8�����&ӂ,��
8�8)��K��.�e?����&>I���~5�kk�+�lH�-y.�-��"��`�J�'E�,���|��%�������b�ݲx���k�b̫�vJ��h�b�XT�7�-dW�3����0QD	3�}ݰ��[�q1��Lq ����!dq��̅4O�NC�xI3�$K���G�3y�3<Y��q� 5X��5�_?f<B�ݮ_���Ͽ�g=��X���={��ݳg�wp���/4�8��=���ѳ*�������[����c�=�K,�8�퀋$�� �9�������"���%����f�[eK9
H��ʋ �_ˑ��
���|i��Q.R�+M��0�Q-1�w.[��
_���/�W��]n���x![�hc��Ʒ��j�{��U����H�1�
#O��V�?&L)WU�䎶>Oy[�~�/S��jCsS�u�h/7~P!���v�IkH��
o)/6�8����U/zBb�,.�����/�g�|�,٣,�(�jL/��^�/�x�Z
s����LkS�?�t���g��{����#¸�����HQ^
UP�Q�mWŕd�SHc��'��M��q8Kp�UwO�e�*3A��T�e�QJ�7�E�W�W4p���>7�Lt��W=�貈O\�]:���Ą��c̣:aܞ���������;t�t�^\�Z��Z��<�j������c��^�\�"�t竚%��1M�O)��=s��9���⛛�:�Zh�К[X���~Y���fׂ׸}�0[oW�u��+�'�x%U8G�^9�x��ܺO��GÜ&����"��r���	���@Đ��!�����p���Ͽ��wk�	�=?��ALh�	0�+��	
{�l��gϞ?,p١0P������'��9��+�vH|�͈�I���5�9�rA݁[;���y�@u�Ꚍ��8��!�J��,(�)[ Hk����T@U-�ȹ	����o�Y,KU)*m��yV����	�1�����R�j�[���o��$*�3dnK�6�\�*g�Ƽ�q׿w9,�K<#����rZZ�j��_B������r����{Q��5����[|c�0T#�dP;�f`7�:�ED����F��􆚢[���IQ���V��ܲ���2�)9��{��#Wr]뎸�kfօd�lv�r������
,��Pz<O�$h��~?�e�x�ǖ,��]�$�+�Zq;322�n7/��ʚ��b�2++kU4sČ1���חi�I<�PR*N�C���#@�*m��Е�s���
Ι��GO8A�aX�2�C���i�����k���B�#p8)!t�������I($��4ԁ:�Ͱ��gԺ��Zk@�9	\�T�%1���BT�U�x���/Q���M�b��1�t;��*�;���k���4�*��H(%q�F�c!�y�(�z���.Uk�8��b!��!����9�6]5�S+�ߊib��Qab��@H#y!d����N�](�~P9�C��\E/�����9���R<�ŕ�U�<y/D�Je�`gX���Ӏk�""�(8�D�@�5ƺ�-��O�d��H)>��Cag��+t���6N�B����> H��S���0,p�y+��p�aX�Bon�^��Ul�J�АD�LQUTyB�֏�KAh������uU�J�[� ���p��-)c�'	�\�t)N���	/ �،DB��`u�jl�ن�	����VV�|@G���)b�LR+�X�	\x4�=�1"�����D~�!{9seSl+�>l$�H�4]L��F��k�P\3�rR��f�\)��Bv������;��
E]4����������H���ĸP��j�o��I�y������)����*ԺF.7[�l�6�A���蕕���G��DD{�ܙ �k���8�Mҍ��⭉�E�:�Rh~�d�ü��u��ְ��M�^C(���IX:�
*�mB�2�&EY�PJ�i��MUT!b%W	#%�l���@Pj���ΧIh)�?D�p�r�R%�j-�Z2BN(�e'���b*e��$0Þ���������oKĔ>���TѣI�R>����5�J�;Uf�hHeB�m=�-G��F1N��a��K:3�X!���ژ{� 8O�)Dn��1dy�o�j��-���>�#�'.3y�wC�\l�>�d�1N�/Σ��"�,V@�ɡ��T��I���ZJMn�ҍC�6���4�&K�$v��j��pɪ Ӧ�v�)�98OD���2}��x�0�@U��f�.�0o�G��>��]��yB���)�( ��x)��A�ii��r>6�����c׺��uU�i���U�`��sΊbj��5q�Y��!�B��4�5�7�o�l��Z ��w!�t4�� 9VC��Ѥ��פ��R��f��3��/��y�s+�1���{�Su�^����kDYeFa
(:�B�*(�)Q ǜm-
�
;�I:�&)HA��[=�wt�H��x��B Ł���&4M�11@ӽB�@X^�@��e~�Ͽۼ���ݑ N�)*(%�u\�.�mrZ��k$�jTM��1���0`��4x#Yk�2�e(��(��҅����qd�ϛ%����P5���"ð�e��=������x���x?�a�@H�Zo=`DJ3P2Z�b�|I�k���e�(p]�nR��H��(8$b\�3s�OM~Ec�y��1�T��d� ���X��L�V)��96
!_��Xl���U���T
� ��0�J �]�~7�5o�ɤH��P��%1(�k+�SdY@ѻ}�;�^�(��R�6�?���S�;�7@@�Tu��/B���D|�$�&RH�ع?��S��T1.�x�5RάC����6��6%�fC@�'\�dqЕBUiTU!E���!]j*�v\�JאR��R�uWǦI���d��m�۸�@3�R:�j���Z�i�r�ZH�^ѫ�
�<�`�.�0?��_�Z�J���_|��x3[h)r�1�z� (o�h
��3!�J�s��;Fqdn��@�jkh��j�5��@���>lgjM��8�٨}��������Bб��K�7$����
��'�j���Υ�T�ˮ%A/�G�A��:�����Y���J�
�r,�s䱵bg��Q;�\ۇ�4"��Y�ɲ"OǢ�����������K�C. S�8������ l���>=U~A�Q��&��g"���	!�8�"��ݹ���@�QE�s�<�PJ���Z�&5����p�§X�xْ�B R	誊	J�͜Hc���1/��֧���)Tl$B���a��m�dS�VCh%*4�
U]���0�a��0�۲�����\T~a~b^ �8�y� G�. �����(Q)�u�l 圻�i��U��B�q�-:�$,6�,,�痎n6�	�l�U�K(Xga��G���*eJq!�Z�]��U4�J&�,�0J��I:g��E��1P�ڠ��ζb9�5��/L�p �����t�i|+y�IP��3��K���c�w!l_�n��n�Y(p�S:�M�	ڝ��H{��mbC��wM�t���/3��(~G.p���9���OC0��p� x�\���$�O�<���;m��:���l�JB��t)e�!�h�dS比*5X�(p�p�#��T�G���P�����ڟ���/�_)�a��0�;�>�������F>��j����L���-�I�I���[�!eHB���(,=v#�b�Z�(�ԃ����f��Ϲ�ٛh=fG�*e�T	Zkx������
AH�4%�yx@z���U�W�ԗ���X�B��*�OW�Gp�`�YxB��п�z��? 7}������$D�L\�D�����`:�ⵠ��Z����oS
�O���~��A�}�6��F�n�v�"$?nq_ �n����mR���+�����r.�al�ଁ3v�@�.���D9���h��n�t9cfc���Z)�Beq/öڿM͈k%$��'��[T����&�����5��|��aX�2�tO~����?�u�\hiD�>w���|�f��c���!C�����`JB`G �|X��Ԫ��-:C$��l�Y&Ql�]!W��FU���<��R�R����9V�����䷭�Z�,�B �Bx-EA���(�I��
BȜ�u���7L&˱X�B�FSD۴���,BĲH�?C�؊=Q��zH�^��i�jv_��kw�6�9������.�2V�_�\���g�I��z��v~7yC�b�nL/���/8x���
��w�:�ӈ����J*4u����_�a�	�4��n�!��		6�e<|aAB Vu��:Z|`\�O9~O 8%5T��,�明+U��n8��aX�2�!X�=�p	 7_��o&���G�3�89��y�qX�N���������7Cʳݾ/;�`��1��(p�
ݦC��!0�&e����/��t\�S�V)=i(������t_���P*�s�A�!�[g_k���dS� ��U�m�j3\$�밭�R�D)X_���m�Z�~�uf��ĥ$1�*߾��&�NI��E�v��*�Є��CR��l�>i�m8n|-e,��/�����/s�,E(wQ��3� o�Kٔ��4�9�-����^���r�4c3lP�tU�2�bc����0`�^���ܠ���u>�z@�"G8e�J!BJq��!�z�eF�T����@'���?:B�\rsð�e�Cs��__�����8�Bv˟��7���qk'��`�6�@���X�[3c�&Lӄ �2U�ۆ Hcl�;����)��J��1Y���k�M���Q���Q�ʭ�VJ���Z8���1�L�ѫb7b���w��͕bg ��J��nCWL�ڕ�;C
? ����>�gSi�����>U?}(t(U�e�rg�pY�VD����	d�.Ġ�rOA�l�^@�ײ}%l廠���!�me=O*����{����E.[���Ƨ5-
UUaj&�M��a�����Jb�U�E�<��[�N'dj0�PUtU�5��.��I"A
�+��Z8�R6��CO�:�.%!�}����	���/����2�a��0������o�����_,��'�n1��0�%�� c,�pJ��Q�b-�
2h��X��Z7кI�KAH�H+m���>KC϶Y�A�J�n4M���Q7��_)U��h��
�<�-=�ĳ��*_��!�t��0�,Š���em;���mՖ*���K��T	�"^ǘ�
)�S[w���&a)�kٺ� �6i�b�q��4����2>-j�b�nA�M����ڭ�����~S>-��$�� k'�S=�����+��	���.6�y�4G�A�4�A�6��Ø6^�VU1X!�8���$d��+���BƟWU����k�Ҕ��n���i}BV��ആ�5�Fw|�nu�����ݓ���0,p������_|q��?������?��<�n7k�~{���#J���I%�Ӵ��U�5�Eӵq�T�ߺ�'�6���?歃OY�6�p>6��*Z��A�X�m;�u��*]C�(b�:NU��V!�*�����aR��(!f������e�V�8���q��x-� �H�I�������DP.�9|���m�o:�'��v��WWV\�=bv���d���<h����W��g5��;d6$Ǳ�R�cl���1[�i�!�M�[�f%8cc�u1��k�y�w�4b�'x��:h� �����*M��J�����GG��4oB��F ��j[��Mߡj[�� am��+UEyӡ]�Pm��+�nЮ��.�_��|���-ð�e�?��G]�|��/�����~�on�1�phj�J+c �IG�QDVM=�u��kQw��p.`�f�٠�{x�ଃt^Hx����Z��7�17�Ϙ�&�	}�@����M-�d%jԺEUש2+�wW'q+��������B�>% ��/����;�a�y���b�3�8?U*)�5	�M%�!Q(���D��;�Ҡ�bllQL~M��Wx�,;Mi"dA�vz��a��9U"l��H��*��{I�����	_��(:���
��`F��<�l1��3M��n����K��Y�p)tS��:�]�c��W5�� ��}��275ƪ��7�����]L1Ʀ���;P�M��j�~�B�������E�.�/��+t�D�!����n�_������-ð�e�?���Q��/��0f�����������n_BVU����SɄ��������Q�񈸮*X���]0!
�ب3IPQQ06I�!��I�I���� �j��D�k�M����w�]����-A(I5��%�Jɢ�J�3�#P�ņm��;�V�������A��҈Yʆݙ�g1�j�/[�[MJ�y�E���ҁ��Bl��2�
��{������؋y�?;]'�Tp����ɬp�l���RT�t�ϊ��	5����`�7k�\��4��[?ϸ�y�o���f���@����=��A۶�t��G������M����ZW�MJHPp��;�0ΰ>�����y�q7N��&�ӌ��b�:�������%�n�~y�f�*}�����}���%���0,p��_L}���������Uu^�5����®o�����ᒟ��Uՠ�z4}�D�+�´1�	FM0���1jL
+i)��*��Jtm%$�9E��3F�Ԩ�]�a�Za�uh�M]�j-���]�ljfӨ��"k�]-;�C��t;-l+��گ4/D�r��lӢ
j�I�Υʪȯswb�/��������� ���!Y�UWbWB! C�ǈ����י�yjI`��(�݊�w2(T��V! kb^l����n�0L��o�1��3�Rh����=��W8==�r�D�6��u+�R��F!��N����� �Bݴ��L�3Ͱ�C�����/О�a��1�����1�n���ͥ����ֿ>y���-ð�e�'V�G�����������ο��`��� �аp�ޣ�����X,W�M��m����f�yF�" J�ʭL9�������ZjT�`��F̐J��X.�p|r��r	��T'��P�PAA� cc�u�*��S(	��nD�K��T�?%�g���$U�� ��*��P�8�%LO�^�o��n���x,�;�vo��ص'�4�.�$r�Y���t�ȯ�5��(j������_��I�ݟ�>�RWq|-���qL*����8������9̛�<�YUh,�=��W8>>Q�
��J�^R�T!U�J)k!��FYU1�9���^
�*f�zc�tUC��j��}���~����K�������g���e����Hwz� �����B���[�Ͽ~uLѯXU��"&�9� P�ʬ��])����TA���� �HG�'��OB)�A%$U��mq���>�у�PZ��w����X��Y � ��8$R�5<�_'�y�l�ΜY�q7��B��	��^ۚ�(�ERC�������%ok�-����������+�>�����l9������1eCQkr[ώ�b�1��V��U/+Hx!q7���[c'�J�oZ�=>ã��]�ղ�b�@۴)�BFk�syܳP�c+h�$TUAH�"���QX�0[��<�X'$d�����gO���'8}��rurzѭ����.O�Z�0,p����я�������|~��7،#f��h��ԧ�q�X    IDAT�1������*v��&6�丮��Q�5� �T06��$0�����D�X�>֐:V�ONq��V��1_w3`{��l��X�&�m��H"G�A)rLW�J����l&^���RvoQ}}MR�]1�c�S���*}��6��$���5�z}Q���}a�Y�<�� !P���������F��5�u�Z3|�Y)r�:|��(���i��jx�09����C@�ھ�у8::B�dL�PU���V��Q�R�Jny��V�`���6����^��	z����|���������/*]�������4�0,p��s�;Z���?;���iXcs�
.8� !���n�r3 /�ѷ4�!
-�4��0� � ��V`�(!bޮs�������by|�~�B���M�,�9*���#SdW�Zn�<P�R*��e0�B�qm�LNaO��4�U6�.�w��j��B�����֬7>I�s���񶡲�������7�s�F�`��l�ss�W���$�C�y�=;�,��!�"�)�P�w�5'�x,c��nz,V+�q@WkTu��'e3�4$DJQKH����y�G�������K/߇ <d�ayr��g�/�������_,�G�=~��aX�2�g-pOt���߯<s�ׯ^�n��13��|{�<���5�̀�j]��*�u�����=  c,��Q)+�>	[��]��&y}Ӣy� g?�1��ե�B֕RB��-տ'pAqZ4�7}U<�VB�����?��yxy���s E��w��}��]�b��ds�)��o+��Ui.�[aG�z���zx��!W�}��ϥ�硨$���\��1*����{�~�Zk�-��<:�����
����͐��!�)�Y)��o=���)�� Q�&�뜋�lF�0��<a�'!qtt�jy�}��~�c?|�E�����[�a��0�A�X�z���-Ϟ�_}��wW����2��
�uP!`\�������k|���U�, x��u��Z���Op�駨���^,���y���sL�����7W��><��;�����<�,�gk]�5I� �4ڶC�k�y�����aϿ���0_�i����s�}�;;`�&��k��lOt��`���5Q�{�i�Fl�	u���}�O���p���R�Ϗ}��aX�2s(�G/��/��]����^B*����VK8�plfL���׸}�b�h�
����<Y�ӄ�̐Z���P��X!%dS���?����G��/�T?��S&����D���ů�}u��z���O�������0�k& �$`0�84d��<�4�ù8����Lӄys��L�����#<x�>yry����~�7��.�0��ҍ�u��_`u�OVx��'8=>�R�y�〛�k���k��5*�r��������!�1��!�������O�꯰:9��m��W����`  ��/���?|�����7?���K�^_c�Yc���<$,��!��� /U�k�Tl(����	���a�gX�0#�nqv|
yt���[�a��0̡
ܺVU۠�z<8{�gO���gX����b7��1{��&���45꺉Hww+�A)�y���z8�a�ű�X<~���g�]����-�ϳ����?|>��X�����k\�֠i[4��b��[B�)�.�􊘿� �����Ơ�f�q�q�1���[��%ڧA�>�::���3\�aU�V�B(�������1��a�Z�����op�����+�ܬ8�=�n��� �N`�S�����Y[�r��3�8Fs��[^<�����y#��?�����}q�������;�g�<����'8zx���)�����X���	J�,��b	)56À���dqp���F�/�ɧ��Y_ꮻ��0,p�9Ta������?],���]��G������_�z�/��^�z�/_`7�����kt�u�^��:`v@��e�z	�<���c4�\1c����G�l-����
J}�	���8}�m���f���0Äoo_¹��j���
�|��ip{s��@)]7�TM��>�ݢ�Տ��a��0�A��Jꦅc�T��0��f��Y�o^b�8:9B|�S�"8(UCU=���G�),K<���X,�/�n�3���a]_����Ï����0�������ӿ��������+\��b|����ǯ0�O�<�ٓ���P
N �m����)���q�7���o����|��.�0�.,t���1�#n��899F�v8:>���-n���<X��l��yL����	XP�
G�<zt�e��x��1W̘������_��?o�V������i��ӏp��	��
߾�#��w��ͫWp��իW��˯p�^CW5����b�gl�M���Mc��_|����+�0�ɗ�a�q���g�����<Zay�B��Q7-��F�+(�! �Ǵ�0n&8�����g)�.z,��h�US�)��ӿ��/��G����v	��f�?��O����������߼�������u]C�i�pww�i���7k-�����?����2��_���0�I�:o-��PR@J	)�))E���<�W+��n`��36�'Xx�P�]�]�<�[�-P��u�A�Fjr��b�[c�FL�=��ӓS�u�'����*��i�ཇ�J)8�`F)չ��q��9��n��a��Mc\� ������o�8gB�R
u]��:t])%�q�1&>�@�"��D�0�Κ�H��n��:,�]ע�+(%ѶVGK�VK� ���6[�9�y����Ͼ��Wq��\��oj"()�����>�Zk��g�s!@J	�5꺆�u]c�gL��5B��Z!��/2�6!�:k� pzz�g�>���5���  yt0<�w�����!	\�y� �D8��<Wq�.�0��oC�J�	Q�<c����,	�$X��۶E��h���&?�R
J)Xk/������zB@)�E��>�s��
��1I�ŋ���>D۶h�6�4H)�ȵ�b�&(�_e�a��0�=��T��vl6Xk `:�%�u��%�a��vG���x�����C�j ��������p�$���f���k�}!ڶ��۷0�K)a���α�e��
{p枉�$,0C����<gA��BUU��j�㨔���Tᥛ��� ���?��m��6JT��?CyFku�睍=�{ ٶPU��zg���\���"w���S Y�N�#�
�-�\Ta�Zc�����d�����R��Z��Oi���	C�{ww��(Uui���l�X����a�/���0�mW���HH�h�R�9��aR�,p阘�E)HJA�0o��Y��ߴ	��	����6C��{crE�l��]��u��aX�2s(��]סit]����d&��G��m�=� r���P�RR�˦i�}�@�+�Ƙ|!�i��Ni3&�D�4����"oȼ����a��0�=@k��-	]���U\�}������V:{&٢��Ϟ=���6Ft:@�ϔRh���*o�h���BK�[��2�=��K�0�zӯ�*G~i�Ѷ-��OӔEG�S3��6��3��h�7�e��/p���|z�&+�w}�a���\��\���X(�o��ι�*Um����߀����GVJ����8b�睓�rSE_g��v�c�.��3qKb�>&B)�
F�z�RY��cH���N�.��$p�i�7DB�^�����Ib�a��[�~	
O��R���l �����=�|���e���.I����R���.o����P�`��0�~Gb�{��_}^��s ��E�R���_t�Z�����b�yWq�	\:E�$����2����=?�0�Wp�Bx��:/���]��iv��覲q���+���Bk��k�u�7��"��y�Y�i-�i�A]�;2n2c�.��#�E)�X)%ڶE�u;[j�)��4Ռ����	�y+�q��u]�)ni��OO(�g� I�2�s���q{ಬ�$t�t�S�U˨���:%��1�2=?��`h�f��1&�{��� ��MU��r�;m��I��a�C���Ǘ ~Y
\	eUx��X�D-��K�������%_e�m��0�-M&���TY�-?g��z�ηi���C�4ϯ����J3\�a��������ϨZVg(w��I�j�)�F�G$F��%�[��l�0X����9�i�r�-�=�dA �fd�������<CJyBx�W�aX�2s�<wΝ��k��sDIT�� ��B�4�Y6��� ʡ�6|���g�Ξ��q�o��4��(��֟�2�&�?�Z�st�1�X���0,p�9`�Zc da�]�K$r�һ?팛y������s�ޖy��&�zK7k-�}=��l|d�8E�a�o
�/.�K�K"�{�cWx�s3�[�"��*S%�l2����p����k�a��2�=�*����mr�aÐ�#;��2����0?���
<���	���А}�[zoi�Ek�Ԅ���U]������SH0����	@�o�RJcpww����Jy ��0o�RJ�u����X�Vh����$��Ԡ�S�yn�������\��g��/u��5Ak��i�X,r�~)*�y�8�9i��!�&3�m�Z_ ���UU�Vu�ɱ����m�Ik����QSJ�m[8�.�����0,p�9tqKG�$n��L)����u]�s�8b����N�G�˼�?���^�}�����i��iU
\���Z$�K��d����ѣG���0�q͗�a�T��Zg�@
!�u���T:���q�1p)n�O�y[������J����HI	e.�i��G��M���d����K������h�J��_��K)w���؍c�˼+��hi�B�4M��Ck����v���F�R��sV�0\�a�	�q|��֢i��ϳ�e�#��E��a���noo1�s^�M��{��i��\J�����iv��0��a���~�ז��I�RdX�9�^ډ\���l\���د��pww��/_����4�V]��ޣ���K�Z�u]�m�,��a��0�=M�d��aԸS�Z���Hv���&�Ee!���z$%#l6���A믪*�}��/�(�=؎����R@3��a���)e��g����)fT���&�����v�*�3�51
!�ԼRĒ�AJ	)�Nl5��H��	RȼN�a��0������EG�49�����#�LG�t�A̻�I�B��%8)���ni�5�s��
�Z�V�|
�0���;G����_�K)��W	Z�����W)n�x쫕F]�ܭμ3WWW�m�>/-e�b��qa�m�m��j.�BLӄi�rTX/�����pمa�!��R�s:� %�NR���&�e�M*	�U���e�aM~��>��#��]���qrr������L�R�,zi�E�6�d��TJ�3���p�a��{GB��u6��E�y��K�\V��۽�H��i�.˱�$`W���%���i$b�;v�p��]ס�:4Mk���Ǐy�ð�e�P!�-u����3ZVmI��oQ(#ļ��RJ��1oţG�._�zuA�a�Z��m(k�f���9�s��so���j�B��e�3��1�=�-
s���c������/r_�aW0��+e̻B��	�?�T���j�ߘ�A���b�+���<ڗa��6��y��z�ƫW�p{{c��z��D�l�\��^�hU`%��e��>��p}}����V+����%� '/0��a�GJ�K �J��Rӎ1�0��o�ŋ/0�sn��V��Q5�>.�m�.�m���b��l�a�z�Χ	�9�u���!�0��d��C"x]2\�a�2K��r�y�6�%_#�Z�#?�1u]c�g �{r�=7`і����i�z��<q��	���?�9��f�DК�u�0,p�9p�s��)�:��:�"���$,(t�g�u����0��YJ��f��i�X,  G�Q���2�.��lg�a��ƙ/�>�ZG���WLA�9V����19{�b��ɇE.�m�L6�aȍbmۢ�:H)���/����K�.�0\�e��!p������w�e�� �DV̇��Zl6���@J	cڶ�4M�l6����z���lF�h$p�	}�>�.�0	Z���3�sqJǽ�%�QN?#(Ɖa>��-��@���}cnnn`��8����F�[[B9��#��a��0� �\ ��x%����x�t�.a�0bV����g�KM��4�XhM� Z�t�k�aX�2s�Xk=�ᓘX�׸���U3�$�D()%�yη}k����i���"{1�����5����<c�\�%MY�e��0,p�9`����_�z�|��d�s�8���҈�24����|Vf��eއ�m�I�R
m�b�X�{�o��6Ws�����)�����]��;���q��ið�e�@��?�R���BNF��8w���hK��u:
�4jV�*�!��!T�%�8�0Ơi<z�}�gQ\���^c��1}���d��8���QY�I'{}�Z6���-�Gix	�}�-�վ���1ٓK·i�|��:�ɶmѶ-��1�]�aX�2s�"��dRJ�u���жm������ԸC��>�8���*.�� �1�� @���ٱ�(^)$���@<����uLk����a��0́	�"P�>�n��H����'��Z��.�!צ��8�1���@�`�0do�GO?B�Թ�Ĕ�����Ϝa���2�=�<�ߕJU/R��lV7u�'AK��n�>���B�|r�Z��X,PU�q���noo��9��Al6���f�����_���0�L��W��⥵��3�Z�,8�E	{p�%p�$���*ۛ��,d)Ҏ��d�y��U���Ϟ=���	_\�a��0̡���ｇ�2^�e�>5��}��+hGGGX.��ļ3d���M٣�5M����IB�ؒ��O$J!����_\�a��0�!Cb�-� H)s��~�9�"����ȥ�n۶X.����.�^�NJ�Kq_��Z.�X.�9�v4M�c�ʦ2��,0\�a:ƥ7|���y:ń�Bc���}4ʷ@�Ufޅr*�,������&�,H���Z�`����i�֢�k����Ӊ}K�0,p�90�q�<Ϲ�LJ���3��neV.�z�7��*H)᜻B\�UfޅB�PTJe;���:N�sq�CUU;�Z��Z�}���c!0MWp�a��0�5�)� E�'��	`:�%�M+s��Ҫ��x^)%�y�8;;��̼-WWW�/^�x~ww��;���b�@WWW0��t�rb�M ������B��ݱ�e�.�:R�<�Wi�ؑ~s{��<�e��ct��Nj5ȼ!��J���>SN,��
�9��k���a�l��fI:Q�FH��G������>�s�!r7�R
�;��a=�IQ�ծ}q��uK�<��8Zw��<k-�hY�fGJM(3sK�H�R��0���2�ᣪ��
�$Z�Ʊ�\���?��.��]�%��B�֤�:��R�V@�Xh�q��\c̎��a��	Wp��	!�����P�>�S�H���wKK�m[�Aqa���uGB��a��l �@��X,ي�6m�*��^�quu�'����-
��a�f�Z�|Q��iʶ�2w��XN>�Z�m[4M�� ���]�����6U���a�TF�?������Z�����˗����1��3ð�e���1�3c�O�y��7V��y�UU�a$(�
F��|�$��}���/ϻ���\W����%o-�H�盦A۶;��,p�~�\�9p�yv$liꘔ��9�6��EM�*�5�(����&�}��}�m)p�cK��t����sz�n��6ð�e� !A�/)%�ޙHF��MU/$HS3ü��,lgW�u�����LT b�-M1s�eNٰ�0\�a�R��pY�}S�R�`V��D
!(e�U�NH)YhMj����Y����B�f��) 4��?!`��    IDAT��UUq�a���1|	�^����Z��a0Cu]��%�[�6��WU�����:�+̼Ú���_6M�O�p~��h�:�0�y�'����(���c�.�0
U^�D�}���l0�3 d�K����jT�B�{��UfޖǏ_N�t��ނ�Zaʁ���5H��\��0sa��ܧm ��6���R���}�myc����뵪��ΰ������@��m�X,��IS`枾��%`�����R�,,B��Uv��MdeD=�� \
!.�*3o����y�u�˘0�`yﳰ��)�.PŖ֢������0j�0\�aSD��i�Ϩr��0�%�wD0	�\��>�2y�/�>}z�W�y���s��y�����O
�S����1Nl��<���H3��8s�8 ��9T�/ H �Ǒ������M2�����U��*�ܟ�7M���B�x�ð�e��.���q�� b+,�Qg�Y9�l_��בy�ř<��ZL���4� ��r�45LR��}߳�e�����LJ�S����P�[*sH�h�&7𐐥��q$*�w�y[h�E^[Z���[���)��u�R0�`ǜ{K���+7cð�e����:�	-;�I<�UX�>��3���4ˡ�J"��d������7Y�q������j��\.�\.w��ð�e�0n���U\���κ,p�V;�{��v%U����e�3��R
u]�\�<�Xz�r��j�ʑb<�a�7�.�0LY�-����ZA*��y��ݜ���B�@��0���#��uV�r���$!�v:Y��z�aX�2s�"UU��k!`����R��S�%$2���P�yǵy1M�%U`i�m�H��?�6V�G�2���aX�2s��g��s��P�]���Gw_�rU������]���]�u���wFI��!��5J�	��r���!g����%`�Å��sB�,p�"�lLU QVx��H��i�Y���ü�L�:-�cZ��Fi�	X�d��X1�ð�e��)	��"潇>��}�¾��|�$�/��<��yoJ�AQG뵴(��,���Ƙ���a��0�R6���/���}���ֆ  v2s������3�˼�����a��*+��-}��6�@J��͆a��T�*qr�R@���S�;�ۀ<�O�~��ހRSY]�y��s�8�A9�����"��ҋB@UU\�e��*e�5�ёn�#Z6��� �E.WĘM]�pΡ�{�]�5�i�<��l6��fH��ږRBI����'��0\�a�ar�y�4Y�5�-Uê��b7G/�, �y���T��BI	䡥Ӆ�^Zj���BH%���+2�yG�0�>bd�f�^c�gH)�u����f>�d�:���Ąuv�S�~�}�5�^�q}s��*m�H��[g��$���zL]�Ͽ���s����a���ر TU<�y�9�}S�:Y�lR��|(h��z��0��昰�/^�sp�4��g��9���2ð�e怸���i����h-�a!��n)rw����-��C�a�^�����h3F����Kkt��[�<$��c���\�9pʪWو|��=/mF���s��1��P����<�S��.����� r%���2s�w(�9P���~3M�/��^$p��6��v��X< \�QZ�T�LN('����4R���-��������%`��e_����:��k���z�y꺆��h���f��a PU꺆1&7�9�vH��i^�s��(WWW�M�<���7�g��7M0#�B W�X<0��u]�i�<�a��`�\�%/.yǩrK▢�����>����a��s)�9��� �OUU�\ ;�Q�I��Q1�C ��b��vZ{��|||��a@]ׯm�h��Yôqc�.�0���*�~E�|�etX)Zw�ъ���t�0��Ϫ��4�ֹ�������ɪ�z'W!���p�5�0,p�9@H$TU%�@%�b�#J����$p�Fi
%,��e�Y������i�0��4��F����QB�<�0,p�90���i�X�R�;�~��rp鶟��G�C�o�i�v�k[f�ZkѶ-��V���i��2[h�t�aX�2s �h-�	e�DG�������,p�	�PZ��:7�y�s�>�͜��tB �o:q`�.�0*pK1B v2B�iډ]"�Q����7%.0̻ �ȧR�X��kÐ��s��=�3�q��u]�uN�w$�˩}ð�e�xS������}:楊X���	ü����53�&����8�y� �s��y�0,p�9p�[6��wߦ �ȁ��k!��x��>�<�C 9%����1��4eqL���U|��.�0�%�S$Б.yo�ex~�z�Vr٢�|�����W�^=��M�`�X�H�u�g��4 �f���:u��M%*�.��|��.�0&p�&��L\�)Rz�� �8���2̻ �����s�%��V9������Zkt]�7f;�{{�4����쒯4��O��a�7yp��(�y�U[)v������_�QJ�2�pIQ_uUǬ�oW���7JL �{K�f�>~c��ι1�#\ e�vo�٥���w�����Z�K�M�@*� v���)D�#�9���\�a��0������d]x���*;���i�x��1�2�����s)�g4"ZH��ic彇1���0d�m�ΗNJH��u����ꜯ4ð�e�![zl�o�C9���~���y_�8��7�T��l6�q'���$Xks��k)�y�9_f�a��0́���m�_��e����o�jv�۾��N�*/-����0���S�m) �`��V�c��B}ך�RBk�o�T= ٚP{PJ�Z��/��1���+�sO�4M�l6��9k-���^��T��\�ߗ��0o���9wI͋�RJ����&I�R��(iM�c��a��0�a��,���1�6�i�p}}��z���IP�ӥ�x0�;üϞ=���܄�*-�M���fI S��33�E�a�_��ֳ8MS�9�H �J~[�!h��}t\�\�C����ƫi��iz���f��i�����
}��Z�k�a�s��[� ����xK�K�/��1���֩���P���=�֘�y��M�a��UJ�{�a��l���{���#c�\�f�t�G��a�C�<�%aJ�9$�x���d���16{����P*�1&�hf���}�CcL��M9���>�tIS������0�=�߱�@)��ȿH>G�}��]סi�� }j�1�d�Qz$�C��r#��UX)%ڶ͛�7�c�x��b�{l6�_����0���p�aU�_�-���2K#N�?i�)5�����v�/�|�P���KJ	c�N�-%$�M�OHضm��sQWU�����򳫫�K���a����w�㸲w��˹ש�wR�D�R�j7>� ưA������a��?�2�|Ӳ�d��$��DR�۹���C�
Ȍ̓%���B���\�DF����k��x����lv �O#��6LA�|q��哢��l�h*� ��r) .	)gj�P@D��$�Ƴ�1Ґ*`���6lX�kÆ�����n�պ��-MSѠv>�m�?.
��o\����F��'N��@��D���O�N��0��_�q���N$�a�\6l��H�y	&�� �Q����h��fJ�D�����`�ƪ1��3�qDU!�lAJi�2Y��B>��$I��}Qq�޹6l�xu��06l���1b�-)7f�ch�M2C���e��*����;���w�^z/����}_TĚ�#aq�*�k�l�gA��nX׆�3
pѝ�A��i�X,h�\
[0�+�0�f56X�w����X�����R�r�����$�nmذa\6�`���9y��j�C�� �#Se�`�[�.Ӕf���s�t9Ē)z��M�D ]0�X���g0$�nX׆�38�E&��-�q� ��X� \���cذ��:��f4��^V�eR�:.9�s���č�����X�x-ȵa�\6l���cx����v:r��(_ _���>	�`�\MO��$��bqB���Z�<!I���� �$ID��m��aÆ=�l�8��5�\[��!@�ȿ8��cq�k��� .�*\; -��-��,ȱ�`pQ�� h2�a�ƫV�k����lFQ	�-�(��u]����F�N'jU�	 �  ��ڰ�*��Map�@�%֘K��Z��K���ڰaÆ�6l���<@�<���4�n�K�� p9P�A@.Xaː�X5 Ryb�%
 �i�����랰��Z\���a��[g�a�F�����]�i�����u^2``�Е΁,J� � "6l����H�P9� [�]^��2��ڰa�6�Jt:J�D�i��b�e��ryd��'` ����Pmبpr�G��«��wP�����OI��s�]{�m�x5�Jl�8��P��}��(�� (�&2������P���%:rFÐ��6�a( ���Fl2����>u�]�v����X�X����l�����={�mذ ׆g$��)�q|�ǖ�}y�t�`� .�\�u]1Bպ(�h
���OaR����u]JӔ��)��s`�[���%���$�|�a�{Jٰqo�c ��.�k��E� � ��%"�3Q�b�ӥ >�A��qm4r��)qGT�!MӜ'�*��aÆ�6l�8c� p���W x�� 7�ca+�e��K� �^������6V�-��A[��u��Ґ��{h<���6l� �6�d��/@+�- �܂�� `X���r�F����Eѽ�%bt�06�Ni:��	z��	y� �KD��k[�ǵaÆ�6l�86�`��BL$�KD$�F9#FD9��&��,˲�W��*q�ʕ{�����Z�^�����v�-|�1"�c���h��aÆ�6l�8Cl:��l6��|N��B�B�Ec����^J l[��a(�3��Z#\+�����lll�+ )T�4k�O�˲LHmt�,��a�����a�l������^�uB�F4r�e��RMD�ew� ������#Ib���%�a'�ٰa��2�6l��x��ٝ ��7�L�d�
��ea>]���ʃ lبpS���.���G������6lذ���g8��}���Y{�aHq�:Չ�\'_���eh*C��c��ڄ�Xu��|���kSNи^�W%T`ن�ڰa�D����8�8 �[�	 q<�W���
I���4M﹮kG��X)�c_�X�|t�l&��F��Y��6,��a��\��m�q�b��D����fr9��C��|����;�F#��Z�E���)��k�W#lذ��Msm�8c�����]���{b/�P�  9rW�����ѣGw앶��u�@�Z-��z����=��c c�r�6,��a����uR'�X,��3��8��F��_����=���<�����j��d���[8{`�S���@p�k\6^�6�Xo[���K��usF��3Ȯ  ���0����Q�6VY���$G	�p����Ɩ'q���aÆpm�8� 7;q�;��{�Q�������>�i�����X5�t�I�PE�8�AxTi8֋�i�k��hr3�6,��a����O����we�+w��(?�cj�Z9&�x����1cf�M6��J�X,��}1�2�剡�,y�3���ڰa�\6�X�iz��rӡ�����l��������m4q�|>��l��DDA��8�19�#�-�2.m��O۰a�\6l����l f1�I���w4I��r�ǱE6V �4Mi�X�|>�n�����D��Ѩ*�O��ֿeqm�x�Öm�8C!kU��*���`y��%iB�v�_�>}�3{�m�t���,�h�X�b�81�o4������>�a��z�a��+���a��$I�J���KZ
�#�m���t^N��d
r�Y�G,p���F"�c�����X���4Mi>�SE�\.s ��<���6,��a��t���u]�җt��n���`h����-�`+6���[o�g���U"�"��H�"���:$"Z,b�K�v[��,��Jlذa�g�ʃ8�%�\��O/�k��%d �c��J�l���A@�v[HP} "���X,rβkd`�kÆ�Wx��������
�\n�� t�ǺG����X&:ۭK��� .4� �<�� w>��.��$I(MR��!	��؆�nX׆�3rU �_���vq�c�$Bˈ� �J�6l�>ek� �(���<��	�L��I}pc�kچ�ڰa�d�fi&���z�qL����M����x���8̈́L�������-�8@r�9t����9M&�iÆ�W7�e����h哠 Xe�ޘ`@� ˌ��.������.�$�$.9b{g����fÆ�W7,�k��Y�\!Q ��$�(A@��Q���K!K�ߨ�6�
����*���� C���-�KJ�#��t:��phש�ڰa�� F�.�:��%���$Ih�X�ݖ�Z&�?Ec$V�`��$�q�v�tA�uT\�%��s Wn��:q6lX�k���G����1
U�����P�}頀& ��-���X ��qL���)�i*0���bA����n������C.��<O�1ذa�\6l�Ep+�,���)M'SJ҄�$!��	x�y��hI��6l�ht���8��s!K��-�K�0�q(Nb!i@#�KDv��6,��a�,��`羠I��l6��|&@/7��X1��nK�6��z�|>�8�)� x6�Q�$4�{_߼�̮�6lX�kÆ�3pq�s0�C��\4�aH�|��� W�'�a�ɵ�5[��a8I�$b��.��&I�s�� ׆�ڰq��7�𿣄��� h���?����m�h"ǡ (a�+��Ѿ�#$IB�"�$=�mƿ[pkÆ�-b���`��,#Z���6A@a���Bx�ʝ�2�k��l4v��� ���Q��c���bM��KaR�ף�pHa�)y��װ6,��a���g��-i)���0���(�Ds��_��fۡn����p�v���~���� ����p8�v�}��U��ذa��+Q�a�\�Qt\''C P �@��q�$h0Ð:���m{�m4r�0�n�K�n�� ��b�2��t�u]��ˋ�E�+�ڰa�6�HdY��Q�|pg�����O�n��$�Y,qp��Rx�n�+d6l4��a-r.�� �Y��|>'�#�|>�$IDe"C1�Ć�vX��g$�={v��n�0hy-�8�$9�M��:�Q�Mg*Pb�F ��l�����5�ig���ۄ�Z-�Z��=�lذ ׆g"�,��y�.Q@)�_ �ސe�K |����rm�h��Ma�߹!�"1�CK�{\��Z��ΆV�`���)���`��r��4;����K-����B����v�����E��-�:���� 	��}Z�5kÆ�6l�8+�AU��r�hn�~A����"���
|ذ�Ě�ZS}��8�O4A�")��(7͆�ڰa�, ���/"�:��y*�`4��ѵa�4�+ �z�$���A �F`غ(ذa�jpm�8c��zZ�0�Q��$"�Y�(�ۢn��Py0s��!# ��� ��h6!�aÆepm�8C 7�ca��ǜA@�NGX(-����\Sgoa�DD� ��8λ�j�h��kM$dq���y�5�?1��Jil�x��2�6l��H���(ޠr�:����+�E��8�s`��x�c����˗�٫mc���x��4��!# � �X�x��6l�x��2�6l�������M�@�A9�nr���a6)��h���R�sV`��6MS�Nϳ�;    IDAT׆�ڰa�88��A�8Ή�}_L��=~�hȃtm�X)��D(?�A��b�B���1M��\��6lX�kÆ�3�F��6r����8���}j���"lo�$4���	A 4��ٌ����6]�X�|��0p}-���m�,��b!t�Q	PlÆpmذq�u]�W�}_�X(EQD��L0��� ^�����(�h:��t:�ium�h"�,�8�s�w���Bg��;�������qn�p6lX�k���\���ǝ.�K
�@4�@���Z���Z]�ss}6V�"���y���(K3��f���ł�0�7ʲ���i��ڰa�\6�`��Ep� �;�L(MS!;�t3|q� �.���x�1�����v)ZD�<p���8� ���|�FJ��l��+6͵a�DY�4�$	M&�N�DD�n��8��tJ����9EQt��2��m�$RK��h$�4� f`Q9@e��=r[.�qL��\��%z9��k��Z+�4M�#���^e6^����?~�������x�"].����`qx�j���e]�N'%?7�X�xE�+�q�����1��Xꮁ�]�*�(Vѷ=���0y�{m��O���>��}ߧ ��jeY������qL���txxHY�Q�ۥn�K�VK4�G�"�޷��f����<x@�V˕G�6y�T�]��.[�&{Q�=A���cs�W�:T�{�k�{\��L�?��8�X,h>�W^��/Xv���f{{{?�N��)e���=x��%��(v����e���䦃���~���q��Z���E��ֹ_�Xsu����+[�u__��[���]����gr��|�M~~��hb��9�uXb�3��zн��{�u��yDD�|���www�������,;1��)pk�!��<w\�oe����d����9��U����	�=�(z�*�k�+ʵ�VP0��h�X�+p���]�!�"z��	��f���`?�]$ye@�΁T�����qe0w	P����Ӗ����Qp9��W�e���Oϟ?�~�/[�u�#�,�	�@X�!�]�2׌6�����_@s��� ��h��6ȭn��ek��4�7���9T��*�l�
M\�:2���������_�5ݿ��8�M0�> .�ȩś��& ҄>�C]n�0�NX �����I��`&7�.�1���M^�����C�n�0icc��]�F׮]?�E� �`x����9`�c~��%M&z��)}��'���i%yek���4YgU7~f
pO�@x�.�kW�G�%�Y�Q�ӡ7�|S \��9��}�?��IX�a��qL_~�%����|>2��r�#o�q��V;�MS���)��l�{��nr�rWyU*f���j���d��[o�k�������Ç�ѣG�?�A \�ī���N�V�]�����kʒ�]�eYI�ke�u7���-c�L��u.���o�[ L(>��u]�t��Uj��t��q�� 6�Q���O\�!�;& 0�iJ��<x@ϟ?��b���6����Uآ:�u��z����s�V���%�XC\�����,�v�M7nܠ�ׯ�d .	���&�	�f�ܙ�.��Q��8� �Q}/Mi�>��s���h2��d2�G�c�ϣ)i�Njc"�)c?�\@��ӄ���ֽ�*p�����a�-�&&�z�ul���MLׯ.�����z����MewwW,�0���O`Z�o"�����F���j
��`F���1�e�_�M7��ܚܰ&x��JU�����9.% ����F�咺�.�a(rx��~�p��.��X.����������[����n�E��*��jO1��ĦLV�4�8�g�f�Zu��H������>]�p!w]�q�b��,ˎ p��d:�%��i�
	"�c��f4�Lh<�d2�,�(C!MXE�P� ���rv��DMw� ��պ Z��M���$_L�W]�[9��j"UF��"�}U���ܪ ���U�o�k��O>X�OBƬe�M�-z�h��� ���d�i����n�&6�U���Y��7��|,Z��� (by� ���}��z|rg�f�H^��������G�}A.��n~E�T����W���g���I��K�T���k��|m� ���*���]nӭe>�����t:��b���=��,�����b�kn�Z��s��`y��N��TZS�@h:����J�v����4���IO� �.�-���k�ᴈ��ʘ�*���s��,��*�J<lH��a��tL;�N���m�u�i��e7�*%N�/+�&�=�i��֕j4����T�D͔�Ag_9X�=����@�m���c�.J���\�t\�[�	��n�AU-��%�&ZQ���Z�hN�o�V�_k�^�ebe�[�����e"�Ke��d�$Nh���j�t:���1���}h|��� �i�[�lɉ��xe͉eU����,a1"E����3Y�U��r�`U�N���\(���뫮M9��Ĉ�51�U�����vڴ"�
���r[�oO[dm��5N��W}u�L��7w]��MD�ߧ��*h]�iy���-��و�N�1k�� �B~�n���}_��C
�P� Yw�j�(��Z�2f�D#������~�l㭒 �:~MJ��� ��`3M�*����W��{O� �N�#4�?Hh�(��{�i���X�A���hI�{��j�h4�p8�Y�&W!9�Lh���zUN�ޛ
��$`��]�(:"h��L>�U�Y�L(����)�gR�� ܪ�����NEnYE���X�}�:�Lu<&4��EH�]�E�	vWu�T�C�r��|�m���nfij�֔~X���҄I(:m�iȞ�:�h�y�>�H$��b3�,ˎ��J��u�y>���`�L�#�2����J�_���U�X��VMp�2�U�w]&J�L��2�Aǰ󽈟9���z�qLqrTE$����&1<&$D$�����m����p���h��2PuI�U��*��c��* � ���U��L*3E֪�I _G���ϣ�-������W�u�U:��!<��"��覮��,[�EeMܦY骙VQ����s��z�2߫^����ܤ�T���4�ES�Q2��6a�@���9B���eN� VP�1WmD����F/KT����*��Z��D��s�
J�Xk��V%.��ʯ��	s]�Z^������m��`	b&I�\���_EKYWco��O�گB�T�ɀI�^�L�D�ޙU��5�}a	@T�$���j�w�B�{lLT'�:l�NWU�}<M	D�M����r���@�"�)��\5A:�c�\���4�T�l���e��O�N�E��/ \ ��(���M����q�e[��Kզʦ�W�����|~���j�Y��,ZeIk�w]�<ϣ(����W)��6a�}>�8m�=��V����"�F«��5��U	���ⴚȚ ��^G&I~�U��R�4�w����āZ�֥�20ɲ��0ɶM6��å�Q����JV�T��acҁjZ",kJ)��'@;b�X�d2��0�v�}�1�K���S���2���̛X�"�\;�����[U�SV23=��J|�J29�jH)�MuY��ԩ��id�q�%D�����
�\y�iHM��wy�T�e���#�H_vF�ֿ�9�*I�*ݗ%eա*I�I#��kT9W�&�!��$F���UaO�ؖ�V��Mo��檺�I�{.jb:MfC׀��E�D]��= �u��I��u�e�>���	��{�~q/Q4�T���&#�U��p\�I�{a�V�
_us7}^Y�\��*Ðm�q���H���_.q@���z��i�kd*#kb���X��z�U�6SW�*����G&>�&I����>�ڦ�+��+t��*$A���ҡ{-��јh.P&��>�:R���S��6(5��n²2�*�.;�M�U&��
�J��JXE�tZ륨�_�-���� �-S���_Z�(���n)f
L�]e�W�cȏ��ir��7M��U=L���Z&ć)HB3�ο���ҨJp͸��j+�XK���4���&��
�馩���e�Y��K�Z���ҪMnE����_��mݳ˄̩��te�A������SC�]����Fob���T���\�&غXp�²��&M@U��*V�L�Єα��YU�X4�8Vw����@n�����rH��rF�S�x�״;��L�l3�R�h���p�j�k�j0��UM�e Ȕ,�$֝U>�2/s��܋���ky�r[9�8 �,�)�O4U!�R�6��nSV)����~^�(�j�TIO��-E]�E��g(Kd�Hɪ���i	���Ȩ�>�wQ�(��Tu�d�Zg��I�\�2P�
3\VZ��/�d�A�$V�~���e���IF�1���}n&�*�e�r��T���ZE:�Kg�e�<�|ߧ4M�ky���9i���yb�����%���DF�&��UN)��+��@`���vh�0eEI,�s9���DSG���`6M�t@�*�@�����	�<�z��C�F��	�GZ�ȍ(I
�P�q��!����]�Y��X6E���m�TV�e�{]���W%Rrc�
ȖM,;t�?_���`=��{U�h���q�j��<*"��Tb�`4�d��,�֩�x���K�U7�U�i�2[[�R�B��Y)UY<e7������_�������2�R���5�����������'���s����Ư^�W��X�9p g
�������m�M4���"���u����ݦ��elOQ�]fz_d��l:��|ߧn�K�~���>�f3�/�B3E����u�㘢(�y9�@���OG���˔��?/\ݟM�U>����*K@�6��+���<��-˪�'�ViL_�LNa��M�+zn�5yS2��(�)[���LMK��zE����fj�b�׹�W�!��us&�8�t����_�V�P21�l���s�Tm�&`Ŵ*Pv}Ok���~�5�t0cb���]Ձ���C��jZL6�"-�\��5��W��4�tɛ�N�z_�|V�Y�=�{�t��Z�n�%�'X�X��^�5a�	�3�u�,���*�AOH����٢�N~,� Ҕ�ׁO�<:�ՙVEB���}\��Z'E�"R�.��v��~����*{����TRU���^�'���L��4�~V�p4y�f���U�F��㛠nnu�HԲ��1���+۸ʮ�*e⿗ϼ)f��~�� e�$Ir�<	u�в	?E���)z��|�:Ǿ
�[�����^GS�G�Ϣh5)�W�̘^;��2?d�1�}�K:p�d��$A�ê��TǍ��
�U�})Z�E,\��gQ6իl�Oje6�K��.Y���R�{������(����M��Ӳ�2%ʚLn�8��^r��;^j%�ŪlDՋh�wS����daJe�̭��`2��
 Ru֖�M]2!y,Z#����{�>n��n�V��c�44ᐟ�f�X,h�\R��!�u��n��j�T����qG�/[oEX�����.��-j�*vE�k݄\�e���[X���t�E�sQ�]u4e`�֫jl����k�r��%-O�q�(C �4��FFW����DU�U�N�i3O.U�n��˥ #?�*yT9���B��� ln�3����s�1Q�ĦsY*���r���,Q1�eR��,|�ا���}�1�e,Z�l�ʴ�2�VS�: ��ME��|��s�J���'2P�%<}��e��3㙳|0�ޛ�{�����M���>An��w���׮�jQ����,�h>�����l�@	��i���W�܋�gYNCX�Z�������Mz8d�0^�g��.v��Kȭ�,Y�Y��DKy�s7砠��`� ��� ߓ��5��⯲Ϛ�ݺ�K�̋��Uu�*���������$�/��IH��!W��3rO
>�G����H</�$Ir�S��Y�������ӳ\�Tn���m�?��e����^�[�w��,�+9VIיt�D9r�Ei�IQ1WM�f�Nw}yv��0s��k7ݗ�������zQ4C�f3�]���n����n�j�4+���&�0<���� "����g8�㓚�S1)�ҵ�y�u��(��p���&�rQ'|]�jpLӔ��`�q`w:��zJ&V�2QT(���&�_n-�_u:z��3MH L��� bc�Ab'�'eM?U�W]�������V���;��2��삤�VZ$���+��m��"���R�0�{RQR���y��b���k���<y���QI�L�Z��U��u��T����YY�i���x��	��I�2�U���uȞF��k�.�6yZ���][�&Z���m
�P�&|!#�}�:�����#��� l@�ł:��`�M�S��Wѩy�6壺J�cfM^W �|2��0i�X�x=��ˎ4�99p�	��E���X@xIY5Fv���k�ˆ�����_�\/��tr� aR�$4�Lh6��/L�3�<��~����Yl����	��q-em%L��㟁ʩbՉ��}�I�v�y!?�Ι�'LE̹�y�ׇ������u�]�t:9� _r�R�,��y�3gtr�󹰋�:`Z$��5�6=e�t�F����ׁD�ըIBV��,"'L�Ĳ{�+���0��Җ�T���^>XT^�&�U�U[�i�I&br�������z�I��g�kkk4���N�nzyÔ��8��a �Y�QEbt,��d"���E�;��?��u��*II�lҰU4���lI���׏����@Y��(Nb��g�z��J���yW�P�U�W����W>�X��e<���x��e-��X�/^�k׮хh4����lFO�<������.u�>"7���/��WreWE���A,�80ʛ��mR��_k�#���Ο�Ie6P^?�%^Y�����z��?ρx�Ƽ�t:sيO�r����{��<� с�_H�}�W�[r��e=�9�U��F\�{xxHG�s�V���V���-�}�N�X6�CuO�ؙ:�4�U��:9dQ��J�\v�e5^Q��ʤ(U�^�y��s�s���!nl˺�03E1Hr�
^�� �^�G�nWh��~S��Ef����CNf�!�ͧ�뉿�f3��ߧ�x,�����U�m�1U����ʲ%F�k��l!J�`�a��?G\K~� x�1����}�irI\��:�-s�e���}Yw��?$f�����ݼy�n޼Iׯ_��/���q�L&���S��%�������s�Ip/�eIHY)�(�.҂�M�R%X�Ĝ��*o\R1��sG�E� �L�+cpW-��YE�l�3ZN��m�w SL@;�8�aH�nW�'|p��A ^/$$r�7��3���u����?.�r�n�i>��|6�E��(��VW�.�$e�Lz���**R�D/^E���u	�)�-�9:y��z�$�9�.�b~,3fE6T:f@gQV*�-����rV�j9�L�S�"I�|���u]
�@lX��@�\^2�>d@��@���Z��5�����n�+ʻq�|>ϕ�T��*���"6���6y\0�e�nrM"o�(bUOCndR��2-��:u9�8R]I����`<'ʠY�	���ߦ���t��-��ަ�p��IO�SZ__���5�����v��O?���]�:� 0�UP��J��YW�fT%s&RY���j��5�;���|>/�J%w��W�~y��ԾP�7����Nr^6�]�pЈ3ՠ�`@�V+�'o��4h0 ̭
U=���;�\�@4�^Az��ΥY�TEQ$���De0�p8�%�qrD&I���IW�7p�|L�"u{U�ݲ��UMM�m��������Y��2���G��.�6Y9�)j��.B>`Tk�FV�el�N	������`0�N�#����$�cUpyAp����
`�FC�{�N�� �N�#tV���4�s�i��kյX��3��촎&4�:�6��$Ir��U�UL��봒�"��.��51��pU[�)g�g��5�L���PL��|�2��;�L��'���y��|�2����=�qh0].�,��/�M����)s.7Ш��MK�u'�ߓ��=�xp��FQD�v�� Su    IDAT�Y��֖I�D�\Wݟul�|U��T��1U����6����h4�N�CY��t6g,���ϔ[��� ��N�C�N��0�D$�� ���B|�,���"@���H�$h���m2�������j�	�����:ƹ.ƪ�U�ݤ�l"�3a�� w�~^�����NFZd�_e4l�U�96)���h"KXu��s�Xn�1s��!�z=��ؠ��5!I�� vVUr�_Q
��.�J~]�Ća��#���q��6�N�Ckkk4�i?�����F��:M��EU�Y�yv]N<� χ�M\j�-�V���$@������L�jD�$E���A�I�~�~TW��1-ʲ����hcc��~�mz�w�������+�`�x���ΎH&Q6���Ee���p$1)�I�iBVVa����@�.v��ـ�ւ�n<I��$%t��*���ܛ&��3m�ibORiW!5���gB����W����
T{6ֲ|N�	�d�p8��jܕ��{��Z-���'dX"��
��@y0�x<�7�|�`U�Yt��U��2鏎X3]2iT<~���̱�j��S�,�N�)zA:=�*t��5m�o
DL@�n����g����� ��t:������Q�ץ��5�ʁ-��e���y9�;h���;��?���*��҈8�s `�
�u�F�Ħ�M?�"��J�d��r�	���Xج�r��,�([fZK0�k2~P�F�<u���^�oS5`�I`YCaY�'؞4Mimm��^�J[[[t��9��H7_�I�A��өh؃F �E�ӡ��-����G����^�aew���[&��U�*.���u\��$=�\�,����%7�V��>�$�lz�i>�ΚOnPm�۴��N��@$�h��{��p!�����T������bA�~_H�&���Z���/*�GdYF�v[�y�v����>���w���i2����.����ѭ2|��}V��]�W��~��-#U>�u�I�0Ѻ}J�˪/g��J�U)q��*�ΐYnZiB���4��\�	neL���z��hD���Ma;,(��x�Y��gQ2 �f�ؘМ���q^�� �� �8�f�����z��rIA���%IB���h:�9'4����El��$.�R�Ɠ]��C�T�Ie��9䃪J�`:�{�$X�U�D������h}}��_�N���]�t��������t��91U��ޫJ�Q������Ao��� l���>��3Qr�6bU�L��uS���3"t�Q����fv����ɟ��)����ȵ��ױ�W~����s#��2`nn���ך��؛1.��|/AB2��i<���ǌs wIK�y�u��:4��JN��4�Niww�&�I�B��%��� r�P}�~0���YSR�_��f\���>u���.r|��C7�P�U����̈���ͼ������aU9�M�j�d��
l*�.\���r]�s2~��ʈ�d;/~�p��e��`D,����� Q�)��P�0(M��c�L&�2Q��,sǢ���Y]�)�R}N�J�	cY'��sg�t�"��-_�Cξs0Q�XvU:�乎��rMըF���/$Nkkk���-�ɮ_�.4����l6�uh��a�5�HB777�֭[��>�����8��g�	���ĸʾl2���p��q��c-�h��\]�HR�Vy� tw������ܟ�������1E��*�N�p�������p8�կhQ��b�z=j����P����:,��ߧ�b!@,���Ð��R~ �K���Hz�\;\��캮hJ���D���geJ�U�#2iQv�U!nT���!#�Xx���P�+U����5�o Z=Yg��y\w���-NIˋ@��dT�U�juV�5���MJ�evb*&��$v.kkk���I��@4`I�D �4���x���/<��_�<P� ���ʬ��ق���j �;�Q���� �F����|h�JX�٫hʓl�V��1�c�a(�P��N��,����I�;j�X,��/(I_JSd ³~�TAf��VM�#Pv����u�m��8�)���t��U�}�6���[t��ʲL�m=�A�:�\fp�iJ��4飏>�gϞ�]�BQ�d*1Y��Z�̂ϥ��Q���'͔�K�~Ð����&~�a-�����U��ʮ���Gw0��ʆrT�l8���F��������t:�c���v����s�y�s�:Z$�؟��pr0���4T2 �ɲ��0χ���c�[���}^�����AǓ hww����sf�3�WM�YL�Q����1&�؋@k��h:��`�*:c]s�
�����j�U������e�B݆[��3�����V�o���L�gmmM&��R��x�7p�26lZa�L
 1�`lx� �o2�4���ӊ ��O�%�n�K��P�0 �ta��t:B�+wt��f]v�h*���d��mL���u���Ѓ�3�$`2�oc.C��g9�*�[�����QU���Um>5�uY�.��5,{w�]:w�]�r�._�L�����>��s��TnzRu�s�8���+Wr���lFbm���VU/�J���}!�9p&���H�s脏)�+�hty�oN]�x1M �λ��]Vɩ2��L�����0�h{{�z���}������i���'���>`F���],�j�D�o���p �{�㘦ө �����@o�u�3C^� k���aONVu��j}��~M���(���Φ&�t��ݲ*jQ���ڝ�(��o�4..b5���EP����U��Z
�2"���u�$r��-���I�&�q)!%���t:�	�9���;�kX����|���>6-y�.���e0 ]�gd�A��������z�1��2h\E��.p�� ���v��	�E���%[�����V��&�ߪ�+7�G� �G�t��M��ަ�7o����i8�뺢�L���V���#t��������7�Չ��������u��3-Y��˫ZW��fe�r���	�E-{����%
uH�"�N�&�������CQ�#"� ���4��q���,,6�=�}�*��Cz�e��EB��W8�xR�#�c:88n�LZ.�4��F���,��,7���� �e��=(&�*�����!qt��2y�	k��	��ȿ��չ�l��a_侠�VQ�-ʇ�i��D6P���<_�g��P��ؠ�`�묏���4� �|���,�W�s�,Zl
܆,�� �Ȩe�}����&��ę�������<�żd̟_.�5u�����uC����cb��4�I�ex�����ۨ�!x63���*��<4��f3��ڢ˗/ӕ+Whgg��\�B7n��<5N�Xi��=��o�qbL6�
�y�	E��[�Ф���t]�r�&���T�-Yf�J���K���������ҝ�a:�V^�����\XC��ę �zU8#�����xL�~��J.I�3q�a/�~��;����\b��2y�~�\�;�)�d�HtqO�x�B�g	��ʘ٦��lS�{��ɕ;���W�Md����&�*�,�r_�ᬳQ�D�Ez�&3���ě��׳h1�JȞ����mnn
Cth��H0{����˭]�$Q6����v.|� ��IaC�:;>������y�bc���p`֍����@`��-6n�8�(��1د��M�:oΓopyc��n�����BQ"�]�䦢��M��ڄ�6ɲ{��K��)����h4�7�|��y��p�p%�t:�D��:�R�t)��dk+Tapw�]���iww���qn���O�DO��h�W}&2y�\��4����R�@�ܺ��h�S�BQŴ��^~\~.��K�~�666hccCL���j��pBZ6���;�̈́&Z���3���9���Z<���7���d�πm��4��#<	=88�"�S�2:��D��퉪�\�T����Pnf-#�T�aU`\�W�E͋�{����	�����B+Q�E��E�Ƨe��C����:=K�aeL��F^V�+�F/ӽp�b�^�G�ш�ݮ��WC�
 ���4ĜnhTUL-�T � P����a�̗��^  zZn��MJ>��I����r)XZ0�X�=�z=�q���"3���U9�z ��M����q�������&$'��i��)�UyR��D�\���n�M���k��$I���t��5�y�&ݾ}�Ο?�����G�j�.I��Q>� �����_��`���'�o|��d���Τ��@W5�Gg����
��G6��Ȏuט)K�Ҙ���E�+*�Ve5(�	&������)�ں�K~��-��,��d"�S1��ȣ��9 �d��|�9� �����2q��q�����x �tƼ�ů��g�����7��U���#Uӱ�e����a#@�U�u���Hh.��.s��/^�5����faU�*6�$kY�gO�:�M.p�L{�?�A@���F���q単�(�ߐ�C�}S�bs_��Uy���yV����`i�	&�cs��`%.�oL h�.�KMn�R���F�6�>Tk�����;�N�MOU׸*��ʬ���%�%-o[ �i��p8�+W����A?�я�ڵk���Ekkk9��?�ܠ�:48x����������AaRE���Gi����>��c�t��]	��|o��g��_uL�����?z�&��Xryz���RehI��Y>���U�L|6�v���an��h�J��@d�����\�,#�~�mĢ(	�&) .����$2~�q�
'f��H�b�パ �O~^z�'\Q�\�F#���Wuk�˓�X��A4U�M��/�7�%���:�`S)�Ir]j�3*.coUTv������B:�r��)jn0�Be�})Zp�줮��>rWN
P�������;��Aζ�	��LP�k�N�H������Ol>2#�.kL��ƌ�l�U��?oٞ���Ti~���ȇ�i^>��o޲��<����ou��\mi��A՘��1���c-���ѥK����_�[�n�͛7����N<�n9�V�Ht�j�焉Kׯ_����z��dȚu]��㭓_Ui�2�w^�V��c�{��_��{T�C5Ȧ*�_�uX�{Ǆ]/��ru ��kkk��>-����!G4�	G�eG��lNQ�XM����
<7dox<�v9y���s	U<�pʧ�q@������F�p�d'p1�����@���P�!`��d?E��*I4�=��6�iuA��L7���y"\�ZD���j��	�6rÍ���Ab���Ȧ���
��D�4 ��ݸT��`��<$ ����+�c��b�@j��73b�q�tb�K�+��m@#*d� �r��4��e�.7��ch�a��l<�]�ކ�*a녍��"���lJ�_$M�]�|=��^Ȑ��v\����\&,>��]�4�e*�fM'o��v���ȿ�^�ݦk׮�O~�z���ʕ+B׎��;�9���u�(�r0���<qp�n��ƍ�����H����_���G��T�̋Ư��6'+[ �A5g�TI������u���Ƈ� Ie�Z?e~�e�Y�SD��}�c ��Q�>�F����a��{�_�|���A%h��W-�����x�F�ib�Bun2���	Mn��PH� ������R�
 �+T�~��$"1�4&s�����Mʲ�vww���#ዀ\��U[��=5�P�(��23-3�:2��x���k� d�(��kl��Ed�fτZWm@�~�E �x�dͦ?W4�B~=e@����A���ō�8�h&❩�+�K�Ƞ����F�M�Q���׊��o Y �|�@���)C���@ ����k�͙�a毇��a�u���xS6Fޥ-�u����JB�-�`��C���*k9ތ�K��y"��0/c�����2P���x������ܹs��k���o�M?��hssS��?T���8��={���>}*�Fw�]�t������Wvx���Z�mmm�p8<�ڄm������?ӓ'O��R'�*+��I�t25�͒Gr.OßH� *L׊�ITZp^��C����"�h�	����Iץ�
���DK�5L��։&=�I��2;v�iy9b%`sA>`����5�[[[H�-��w��=~���jݍ��t����h4���u1�Vp>�^��5n�(��8k��}0���p�����bd}}���e�#פ�[D�1��G=����U�\SBG'o��rtR�"��d���{*:�����u���U?�2f���<~���
���Lx���1;�{�r�(�$w���l
�=������!:88���Ca��& #��!�"������pxx(���p��_����ܝ�g }pqxx��r��.�}���f*��^�鷊��[�pSu޽��@f�� g.x9���+�ԘjqM�1S	E]�����t��-�q�]�z����s�<ML~/81x�ŋ���#z��=~���(���-z���ڵk��IH#��ŋ�^W����ۣ�l&�Y�*m����P�%�LL�� C�����-�P>�<��1�8ZE�c���u�����:�`����9블yQ�;�@~�Ġ�E�&/+C����[\w� H� ����3�X�~/�_]�t�}��?~��|>�����/����t�kfCU��G8"�}�,��	�e��5op㍸<��0�s��5�^O����v����$,Z�<q�U��0�|�֕��||˘`}�n�_��+{��.�W��M�����U7�:&�U3���n�0�& ��NT^8���/i�)6<��_�U�f��Q��666��ŋt��9
������믿��d�c���#k�l�@�:�}��K����?.2uc�������JMU�_ݪg[U �6
�qI7L��n�C���p�L��b7��[��_�Kɞ�����I�^��^�Jo��6ݸq���������"���E�7�|C��ߧ���Ӄ�ѣG�8mnn�Ç�7���h�s#)����(����X�I��_��W��$K*�m�=�ʁ\�E�c۱�L�S%[,\�Ċu]�W��D븨;��r`)_��~����m�r��4K�!�ܶ��$y����Zq�p�	'U� S4<}���n��.]�t���x���M���J����a�����r��́Z�����XC��!�=���gYv�^Mm�2��>�X�<ѹj��Qu�����eM&���bek�L¥epW=�MX��vYX�V��^e�R7/Mxrk.ܰ�h��r�����^�"���l�_��3��I�nTr(��6\���M�B�����>�0!f�X���d�`\���˅��ǈ��hD�v�iwwW�� ���x<�8���iy���ǯ�X4��l��ς7@�)�E������C
Rd%��=��FY�ђ��J�Ł-���Mz�7��͛���x�`gxb�f`��-�Kz��}��G��҃�D��n�t:��O�ҋ/�T���۴��)��ƥ8����:W�\��v�M��h<���IEYy\75�ȫ��VQ.��\N�7,��	}�6�n�f**�:`��*�)��	���x���J�$r\�D�����H|n��e��$	F��vooo�����V��w1y�u���nll����>�m�۽�{ �%$������s���ޱ?rm,�g��'�.�n��HX��,��V5ˡ�Y�TU�����4��H���*�*Hm����Mf�����=�ݦ�*���U��Uh���D);?9���G�r�&62��������[�Bϴ��&�+��O�~_l*�w�4<��`��4�n�K���M&Q
�� ��FJ�<�f��@��E%q���"���
en!e qVT�Xr��!�0��b6���An�.{��U�so隙t�~=�D�,����ddYF���t��U���'����z���U
���=��y�>��i<���=z��߿O�1}��W9_f|F8h��D�ۑ��    IDAT�]C^�e�����ӥK��A�e=|�����k�6q]vU����f�Ǯ���8���� �cs7���.�3�ƭ��"u�J��Z�ER8y��j�|��M�mFe�U��"?��%W9&V�����'_�s�l�77�g���J�,���q]�?��wt<�����>I��s>�Ǿ��m�Zwx��t:���!{�v��}-�c�L&�=Z[he�l5ʐq�醸6���Ƈcr�c9��\��n�l�
{ib�Z�G���sQY�q��6X�df� &��TS��*��lVeeΦE�M��:��K  S�-3j������ h��-�)��$p�_t�������S����OZ.��z�M<88���=q��;�_��8��\���!�}��aT��°�;?�����Z�<$��e쬩~��R�hL��e��d2��l���-�4�5bep�,�Ȱ��ҦhO�A@Q)�(PZ�v���?���z�n߾M[[['h蚨�F���W_��Ǐ��Ç�����/hwwW�N�u�=����/���>�H�4�?^��x2���i$q�N�._�,����)Iz��v^{]�ܔ��N�s�{0O�9(ᠡ��i�T,iٹ���Ua�����<,��U|p�sOY��{�G���a�彔r�y��M���~1*������RL��~�>��pH�V�뺿�<�w/^���r��{D��ӧO�[.�w�,K��z����7M�;x<���}���a�g_�ݦ�l����Z��I�1p��n�`0ȹ4�-7'1��E�ͪ�/W��u);����*��&��U��R�߼�Z%#0��R9%����,�t�[]0j��"��yS�>�7&�S//`�h��?nZ<�?�z���N�c����i�������s � �8�����܂39(�sSr~���{�C��j���:�Z-H���k	�!\?Ά�ZrS���d�hPu��	F�m:��d2�Mؑ��0�آuX��RQ�^����*�q�ݦs��э7�֭[t���Bc��)UY�O�;88�/���>��C����ѣG�����ޞ��� �+dC_�5}��'������O���A'���0�+W�����ݥ/^�t:=���&��sA�@�$���)�{r��֢��u{��勆mཨ8�,�A����Q���`�l�[7xqS��L�[^Kyc������6Y\26��{a���{p[�V��s���+����?�3�~��{I��M�4�}?��n�w`�ȭ��u��X7��h����x�\������$�W}�Vh Op�9�F�`���@iQI��ɓE~U�d9e�n��i���)EU�����.+	������HT�/eF���B��/�p�;Yl*��;��t�Op��!�Y*n�^�'�$.e�f���_ӷ�~+JE|��ښ8�x�/�����ŋtxxH�N������amm��H0��\	���R����Ǖ���Y��x<���|>`X7����p��ˑШ�:q�2��Gx�`I��xS >[�FNN�l�Lt�e�E������I��I(unllЛo�I�o��ۍ��:��S��b��d2�O>����?�����?ы/r.%�܋�Պ$I��ӧ�����^�xAO�>��_�.]�D���"!��!aSi��4�N�C.\�۷o��O?�T�����j]��s�Q������Zቻ<
�����뀬icXQ[vޙ7Q5�q�P��|?�gH��%�����DG.i�J	O��p_�f3�N�����ܹst��E�t:4�i<���Dto:���u�����?���x���s������iz7I�x�X�<����f3Br��B�N��vH�~�m�[r;^�䖙x���=�I´�\gfj�j*q,��+��"�ćW7�S�tWm��ݟ�
p�Z�fȄ٬�E]�U�L-pT��ASc��U&qB��������%g�WY��`� n�0�0�q�����vigg�F���sz��	}��7b888���]ᵸ��G�{i����t܂Q�Yw�4����qȧi*�`80\�tILis���)
� o��'���m�����F,2J�8 re#r�
]٦�&��[k\��2�x< �;N�Vb\o&�7rSs��+�F�'!UoL2՞�;�M'fɺY蹷���֭[���H���q�T�	����!=z�>��3�������9�w��I|r�,�[�n�O~���O*4�|��\z6ikk��_�N/^����b���Vv�e��U�:ܟi�
p�'�$	��e�#�l�-���HbF7�W��A��ٕ+�"�'�X_�����7��b�a�
 6x���[��{����͛���)��W���z�ߎF�����ܣS�0��Or�0����4hkk����`kq�R�W���@c'�Y�9����� U4��*8�hLv�=����U�S`�}�M{�y����Uo���R�XR��_d4\5sVe�NĤ�,�MXݢ��d���*K)I�/W�GVE�`Iy�h��(Y$���ODD;;;t��E����7�П��g���(MS��y��5�8ν4M��������7n�(��>|�^Ew[�V���q�����ߧ/������K�L&���t��%��ݥ��]aC?\�ǳiX����:c��.�H�d�U͹�+Ah���n�5�+~����<�Ek�
kQ�L'�\���Z��١.�����:��|���b�� +��?��>��1�����u�4�p�����i}}�._�L�ϟ�~�/���&!�~����йs��ҥK���C���osvI�!���X"��wX�׍Wg��)Y��ug��{q�	��U�]u^A�ם�eMRr[G���늟c����}b��t:��١۷o�իWE�r���/��\.u�����{�����{��?���/� ��*�HT�����<����s-x u��>y�(��\`?1m�*C^�I�L�Ϻ�����.��Ij��Bu}L���4�u7@մ�n��N�M��?ȸFQW��M��c;��7�y��>U��Z-���too��(ʹ!��Ƅ������6�F#�|�2mll�t:�/���>�����h0����i4��F�nmm��Ѩ���ޭ��_�rEd��~��{qߝL&�|>����hD������髯�""��W�
����!�����ᡐJ��>��l��M�n�+P������8[^�Z�6�C*�B�	�q|2��~� 2o �X.;�1G�R�<?�$t�� ��V�z�mnl����� Ȓ����)M�S��>}��G����W_}Eϟ?N\3�_����[�8��` ����6u:���4�':.-��ަ˗/��˗�ɓ'�:�D���`R��K����?�ޤõ�܆P�|V��{,|Q���ΰ"�T�=n(�3�/�q�Ke pq�P��+rEg0�˭[�������.f�7�~�ﶶ��pKDt������gϞ��$ɯ�8�){��fY&*���bD;�-�(��ʌ9wh ��\���e֋��ʤqRU5��VӄJ75��/�m��sP�]t.�dh��X�)��9͐���x�4��S)�~�R	���v��vH����8�d2hcc����i>�S��'g;���L�3M�/_���uZ[[�'O���L�~�)eYF?��i4��}����ۿ�я~�X�issS��gϞ�E�]�q��r�M�ӻ{{{w�<y"$7nܠ+W���+Wi�=~�!��8����R��P���$�J�<#����CeE�H��ztQs� ���{�_�Ty�Hn�YL(�P��l�L@D�������G\��sp�;ԃ  �q�p|Ĵ޿�����<x �'��e3�͙���*I�L&��g�	�{������5��-�9[����������{۴
a���F%ˠ���$	%irro����| �BPZ@��Y��A�0B�q���t@��K*��մ\q�M0�,�<��/oP�6Y���nݺE7o�$�����4M�_.���x���l����~��ӧ�"���/f�ٝ��d2�|���f�={��DS6*�q�AJ��@2��T�C�\�ϳ\Q-ccUթUH�l� ����ER!]���\l��mꦮrѾ/�\��L��e}��Qu�CW�����4!�t��y�p�mnn�p8:��l&J*<����->�3��%���/i}}�n߾M�����.\��������!��ݻ�۝��_������C��/h>�ӛo�IW�^��`@��[����,~�r�Vg�^O�D$0�'�qmV�Z� ���L5��Y[�R� RG't����oe҇�{��T����~ T���`�q=��FiV�X�����O<��?��<x@O�<!"���iU�jg���1����o����>}J�����[oх�����2�V��n^�%�&�������TI(|q�ʥ���yns��T���~�֑E�GV�7��5GԤG�)BQ�C�� �ЄE���������p8���-�v��g�q��� ��o��wnpax��������A�����ɺ��Q����c_����CAq'8/��2	Cvxҍ�D�P��e�:2�2��=�������U�LΈZnS�)E^k�6�}���-����[�?���޶8�$���OW�\rLC��>�f3^1�H.e����}�L&���3��/h�\�?��?�h4�����ۍ��ߝ6�Uŝ;w����/7�7~����ӯ��J�ʭVK����uD9��B�5Af���ܭ��j	�-�e�?Ee��Ъ�������6M�E塲�T(��3d�
ͤ�>��q��_��e�df���o�>������Ǣ�����+���#����7�⻻�tpp@��F�mooS��?��u�$+ .�˝TN{�,�����KJ(�_�8�����濪�D�z�+Mi);#M�'�^��)[fb�$
|�%�-��Q�2&>�wmm�666 <w��/�|�Ϳ;p�ckk��O?�����ۿ^.�?}��)��c���I/�h�#Γ)8�$�;�b�����J`�M�rO�J�Z`���2��"���>(�TQ��,cM��yǛk�*)�L�u����,;M�ѧ��,\�b[��]�(��#yQF][[�^�n�䑆r�=�$��Y,gnnoܸ�~����믿��n\�/_~���ǿ
������u�;>��rI�/_�~�/��i>�Q>`������(t�]�W�ijd��)��OۓUK�D�ϒWub��A:���HW%j��b�z�5�YD���.>K.ݑAx=������C���飏>�'O����8�mf8�ýma?�}+�oEI�Ο�f4��������t�Y�.q�� �}���Cɯ�|ϯ�d��1MI�L�7��P�B�
��b�\x��=M�_��kx���-�txxHQQ�׻���~u��Ϳkp�x���߿��/�8��l6��d2��xLB����'�\`cQù �0�`�!�t��`q�M����Cv�P��z�z����T	�N>S�����U�"ݮ�Q}�����ۻ�����w������(:Q�,�5��(�əf���n]�锱������|��Y̦�t~�<]8�������$ed�Q�w&2xh���)���җ_~IA�h4zo{{���Ν��s��.6.X���������/������W_�쫯��~�/\�΢̄��׬�%�u������˭N�#t�����F�� ��8��%7�W�] �U0l�wN5�ș�i�X�������Xʚt��]�6z��L�J��9���{����F����O?�Ǐ�l6�uTs �%|���(�rc?��A6�1���P�ߧ7n����iccCT���7�#�'�	�x�B{(��r�ָ�r�Zn����\��*똱���,��V�2MlS:U⦒g�����e	H�9y��<�~�p��,�뺴��E;;;�����������[�͛7����~������|~�ٳg�n������Ɔ�� ���{ȃ�8Rt�]A���F_��2U��(��`N�ZН#|��4��tI>,�,	�	�"�Ŵry��M���s���ߎ/�UE�&��e \Du7-c(zmE���[U6Z�`�pp� n�۴��A/^�������/��'tr���/�Q�<yB>� �wޡ.����o���ӏ��{Dt�������/������S��ܤ�/��s�ژ���8s�3� hq������e<ͪ��@��*߈�[��<^O�&5�W�FW�p�b�t�+Ӳ�nS���xI��ɛ�8K��>H�xi"��h$*,��(�@�*���s��_x��Z�z��(�r�R^Η�o4�{堻i�����:���8��	㯏�ޑt���io\ו����<�,��<����	� P�5�����ŀH����V��H�8�ٲd��8Vk����\G��to�[*��,�U�����k��6wQ�QY;�wM��&�ܪ�iL��5�j�X,�3g�y��͸b2���M�P����iss��X,�)� ������E�����U�U*�J��issS$L�Ag�d2֒�~��1UĨ��d,ȓx<�4>]��.S�lc�MxE^?~FX���&Z�����ʕ?��HG����_�A���].亃�:��ɴ��U��~�:x��o2��|>Oō�� �t:��	�+0�(�� �B�"��j5���T(hcc���k��������=@moo��<��x<�����:;;���PHmH&��l6s��.l���k6��r�h4�;
	]���cCmf׺�uAK�<�[.u��ȩ  ��b���P5e�>��ު�)�Ћ���+�
��c���T*Eׯ_�~�/l���U\ O^I���4|L�:����d2��Zu�d0���d2I�b�vvv�V�Q��RZ�%2lq]�N������	�lǁ;�+���������\qY�6�W����1S5�񳆿Q&�6z����������}�z
�O#��?�f�����F��dD��w��(�xpmd��tr��M�&�@73��yᢙ�M�t�����Dv�8W�V��t�wO�ò��i����Ϻl���?ݎ�R�(9.�����z���6��rg&��x<.��rI�D�Z��Z-*�T,?�����O��X�������?�N���������b�)��a�E*��z�.�r�ө��FDB����x,� B8+��cCs	�	�z?:<S �Bެd�Z���[5�t��ecrM���gd��`����@5�Jћo�)tz��H \YÈ5�zx�Q,)�͊k� x��bn���X��n�T�B�@�JE���L��3T��-�\p�dW�D>M�3�\������l�b�9�U��&�&��.�A�-��e���y��!�["��ׯ�?==����|R���0%��_Y3W��b�ߐ���b1�'�4��2d"������2�'.UuUl��xr/7��w��9��H{D	j)�J��]�s_&�Օ�\o���|v�|1���BG
ۖ��-�z�n����k�X,F�d�(u�e��q�F����J�B�Z.
�wvv~��_���677??88���?��'�pxr���-z��hww�F��`ua�-x��z��r9�=����Ҫr�S�d[C�5R�����ۀq� �@�?mY��dv�D�t�@�̐ˣ�1��B���3�_I�*������%ʕ\�(O1�vVX�O�j�l��<���(/ۛn���my>��t:�t%X��iZ+N��]i����h$�Ur��sq��R�-����M�"1��O� B���:v�q���PV�F4�L�[M>����nD����o?J�����r��}��-����:��'�*d3�&	A0q��\A�ߊ���m�2�^WY�q���x\�k���<ϻ[�V?�<����~fm�~f�N��;Kk2�ו�t�5�;�x�Y
��ܿ�;&D�����cW&�D"a/�n�i���9��g?����{?�����7�������n�����_���o�V��p8�Y"�z�.�繝F� H!��&�*i�J�.{����k2E    IDAT_4�}�֐<�k�d��hW;��i��i!�d��d��g G��`���F"
��K?+�+�+O�N�ُ\.!��E��8k��ɽKU�:�3 ��&��s�{����F(t�:������@�4s7���C<���_�'W���jQ"fo����6V �&֝'GH�J������\�Sz����/?��o~s��ʕJe�j�뀘�'��~$	�C��Դ��=�[��^u�'.Z_S|Q�����U�ν�
����/�r7����m��j�#@����������V͸d��t�X�k�-�� /r����7p�ٌ:�u�]�q����7o��A�����>|x��?�qy4Q�ݦ��c���� �TJ$d��b��@�^�X�^O?���ʗ6��ʆ��O����o��#>'g*xy\�qQ�G�2�~�f�d��z�5���_�S��^��0��(�i�a"3�$�3���_W�����Q�i2v�㫩K�Mz��N�>��>�<$����ݮ �<�s�w~GM�5���-[�|�J��]��� �ޡⰵ�E�D���0�W�Q*��`n1Η'������x��]Q�l�'ɪF���d&7!�#��]:�'Ⱥ^�x�7&짔�
�L�t��q]W�-71R6�����U�<F-������Tri~x< '�p[�F��*
:S82�J%z���)�L޻���~���O���?���{_~�%��֖8��"��3�� ��i����h��2�%x��"L�J��щ��4�Yn3��]U�뉃4��<�� ��..�&|n~��F&>�3�.B\�+3��nH���}*�5���a�������8��3�ȯŏf�T�R�N$!�h����	�!`'�d����>�Z�:m�X7�"fp�V�; ђ�',����qdss�R����t��bo�H$w���~�/@`��Y��8�n5�$ϫjp瑫@*`���Mհ?��rL�]t�7�P%)a�|�&�Kb<�����3�A��ӧʌ�&
�O��#�pw�F�XWA&�	��p(,Y1�2���	�.	J��\h��E�����g[[[��r��z�����'O�|�����[���j������z�H$��1h @��	:?$
x.|��ݮ ˰����>��8�@�%��� ���t(��90V�}6��^S��]�ߵn|,b��y�N�)�Ɉ�3�E)�N�8`\C.吽[U�E�]55-�#i��6I�F%{<s	�x<�N�#&5�1�V��v���J��֓_�)%a0��P�"�ſCv 2���nS���d2I���
��^lg��M��9~G��ה����y�m9F��U
.m�Bb`I2��������h4p��ѯ�/���~\�v�~�R���>���f�I�BAHBL��:��ˠIb
�\m���k��8�ʜ�֥��ˣ�u6��3������ǃnJ�eC	�C�3(�cw\�+��󜳇�d�b���b�Xb#d-%4��v��ͦx4VA�����ׯ����������JA�w������nݺU>??�o���Z�mnn
7��|���3��l
� 9�N/ c�E����
+Ɓ����`'O��2�����sme\f���!�r�* ���8Ȋ���'{�TVJ2˭��������f���	>�������v�-F���P';�Y��փ*ֺxZr /{#9���F!!�t:b����
��~��ѝ_.��.	\����H��Qq��&>���1H K�{ 1/�͒�yT��i�XP�ӹ�O��O�$��c{{��������J�ʈ��� 10I����1� k�K]⟎��K@�O���ٺj�KM�6M~����.�����L`��]l\�-0�"Wc���y�Cr�-h�x���0MgW<�����x�8 Z�P�b�}EKM������|�|xx(>?:ȡc[��i:���g�N�i0��f4�ЂF��Kk�O��\ZD@��/  4U�A�/��U�$ {%�)��|�$�:f�_7����<w<��d4.ɣ�U�D����2��t'��|���謶x���R%.�f`���*��jJ��5����g���DD��l�l��:2گE��f����|�g�j�<@� @���z�gt`	g	*A ���,|���<�����锪��1�Y[�̀WOdOr���*4(6� ۶�]�5*�*ΫH]ѭk�����.���Z���g�x����=I���m7f�+��EI�B� ��k,z^1q	,$~�G�H��ݮ �������R���b�z�w�?z�����n��ӧ4���l.y�"`A��� F�x,�z����+e��V�w��ȣe�\0��	O_�@'5���9@q��j޹k󀍹re��Tfd�A5���� ��f����U[?�Y���uz2�Tͫ��Qy�P_tkX>�L,�)�J��hOٕ�7�ɃFx��t:��l*�2���Tٯ�̲�9g�����`��J�4�M� �\�k�K���{��f�CJ�Ӕ�f)��Q>��� wcc#B������RR�+�Ĕ���!���nׁJ���s��6��T��-'U<r%�fwiK�Mxҥk	��aү�t�*��N�º^/HӐ���V\,	G��M&���4_�h�Tꊧ!�z%��P(P4���o�U�T&��4�L޾y�f�g��(/���{���T��<_̗������0tmX4�8[��Z;�ƟH|`i�+q���drE[*��؀]?`]��Ě���9D����0a�w]�8���剁�T�|x�%M�c��dF���o ���N�`Z��Q��&9���v�!�^�9C�.�QFeb�X��R]UΤ�1�.�!�sU�Lպv=kL�R:�#'�`7�Ni8���AvW��尜��L�.��D"q7�J}���ˏ=�x<���u��@
L&�%+;���l��
?���y��l�Rmp�c"\��~����L�m�u2�~.�M3�2��n�2*����L&#&����H&�g ��lF�LF��L����T*����]�v���㽷�~�<��n�h4�F�!���ٌ��4�r9�THd\�YT������!)2�������kR��܁��	@O�9tS�l�y~�}������L,0/!N&�v��3�>�M��0���f�2%W�i|�eL����D���**F��]�,�b�T�nM�,gyd-��9[6�Lh1�H8yR�N�)��J�γ�ow�y�ʄ��c�u���l\S���J�faM f2A�\Nż���oߧ�౻�{�ѣGw��t�dh�q�J�I�+1n��w�*������_�T��c�&��n����V��Z(�y��mot�j�d_]3q�&�u]/y!��s
�.�i6��T*E��H�ns���sرɰ�I^���?��O^�`U*�>��z�s�\��j��Clѥvo2��t�H��0���j[��n\UI�3�\��}�",�
G���x���Z� H�aD�}���H�6pȫ������w������u�h��u��@0�^�Ľ�d��2�5�����*�|�X�U�_r_�j��9*M�|.�&���s���2|mM`A��\\�)� 0��!�@�?�?X.����r���M[[[���!��nܸA�D���27
'#�(���uC�_K�9�D��dgU£j,�+QA0��h`WFWrun<1�%�~�k�\�l�n��:��+�sL���j
�.���1=Gx���|�Y"�X�ܢ�!<0\��J�(�Ͽ�������߿7�ɔ�ᰘn4��D}<�X����B��q� ����PЯ�S�%���+�ԟ�p�T��dB��Ep�Ec4�ϖ ��`��MA�&�k����jMƯ!���<.X!)�M&HjP�t:��ǃ�1���7|���|l0�t�Ѩ�,�\���X�p��l�W�]�6�g�U�-Ѕ"��f3J�R�y�;ߓ���lF���{1�/���u�����$e�Y�,�5-�s�	�L&�X,���6�J%�f�T�V��dDE��x<~w<����p!B�?O�+��)�JOn:TUՄ0ۜ���OY�bdug�j���I9�=��5����*͐��ej\XG��3!�rg�Ҳ� �Ǯr�#�L�C2��d2cw��(���ZS��f�e�Y*
��f_�`���½^Oh���Ш��y@��������`���T���:�����:0�xm1�<Q���H��l&|����F|j��!��Ԧ�4�05P��O�� +�����v�Mgggt~~N�j����(Y"�n.��b�(��`t8��$�O$��&���#��r9��١��]��r�
���'�ﺀ>�~��C5�M��|J3$�,.�GD/$8�6XH\����&��*��6%:���`d�=��W�d,��yC�4o��>����R����(��Q8��h��y?ߥ�豽�}������f��r���'-��E��b�"�Py�s�@يPnui�j�j�Rh���uW�C�����8��:m��"�)/����
�ڂ�:$6�g]�_��A��������1�_���Z��dB�X��[y��b���k��M���\��٬`9p8"��l&�#�} 
	Pd�u5�6�#T K���L���rI 
��3 -g02 �P�@��]�>2\`�/��<��y�4���t����lF�n����[z��=}�����fv8
I�ܴ'K
do^���	܅B!�d2��[o�O�Sz�whggGX��F���#�L'J��ʂ�|i��x��wZ�iQЉN���, 
��(%	��!+���b��4�AרK��I�k��~>.�@�6$5�9���#�e2��ؠ���p_�iss����ݛ7oާ������fS뒀�G�L��� �<��&g]c���Y���_�`ۈm[�-�Xefҍhwݻ^�M-oh׃�� �n�w��Y��х�b�G.?�������Wa,����e'�hF��I�p���$s.%	:m�f�dZo���qk%>� ����%�U��:���l�_���88e��Z"02kTE��&U*:88�gϞ�`0��t�l6�؎�OvS��x��D"!�4�R)����.����{��*p8
֞�Xu��]G��?g+�ro[yZ� ��2�)|�#����7BD���5?��m�ɖ��&c�\�/|.��r�@�~���T��,e2��bb�<�#��k���M�`m����$D$d<�do��M�:��J�LN��~�#[���a@����0y�y3��n�f��~"�ki ���Qw��g��[���y��`#�x��ş�7npU�ݮ�ӖH����I]�-{�����MT�ߡ�{k��BA���.B �62��� ������� X�iL�+@!��{Û�P��t:�X,�X,R�V�a��E�d�s2�P�ߧv�M�NG4Z⽪��n��S�$����^��N��rrI�l6��0/W1$��j��i��Y���J.�����\����k�4�q$;\�+_���Y ��nx��0�}����RN��C��[[���I�<�*NA�~�Ժ�MoՋ���� /�ac'Lڭu5.���(5s=�p8�H$�T6�d�{��M~0�N�H$rw�X|�N���d�S4& ,�l]p=����3�S�J���<h�_��
��<P+3
�Q�+ \t�w]�&��z\�<�>ê��d���U$
H!q��זkx��q�>`���pH�^O������#~p �X������Cu�t4�a�Sb���<�� h��@�������a�S~*c��S������uꚜ��{���� ��UN�d��F8K�:>�~�.���)�@-\yz��bR���^C%U

0U��e��a��4��ʮ�&���=�`���.��O����A��p��8��B!a�k>��u�ׯ_������wc�Xɀ�yc�%�R���X<&@-�Jܽ^�
[���:s��������%Zh�㌍jt+���j�w���m^�0���*���.Ǖ��f�)�"�Q �tν�� ������x<.��̪�4�<vyQO�3p�8��3��&:�Yg�G�"���Eԋ*��ޑPp�sA� ݥ�<H���Y�RR��u/��%
)�︖qk	q�w<�>�P�5����"O	E��	 `nŇ�brRPU^m���)|~֔n⟊=^eX�K�Gw&������&ڷ��*��t�M��u���nB�r���X�C��`{�R:9ѐ���3�����0�84(ob*�ኦ�H$B�шZ�u:�l�nnU0h���<�%n�>�Z[$8�-��fj�Xu�6-���.�p����R�F�A�F��ݮ�p�MMx�b1p��R)a==#�q�u��d��c	�^Bb����?�x�H$B�d
�V� � �D��'��	����쑰؋��'r ����PY3��X��t���Ϲ �G�\��7��d|�W��Pb�#�㉠�Q��<���@
��J����c!}B�}�y磶��^��V7t+�ǬK�L��z�S2�yg\�!�Oҕ��ź��lS'��9��N�2����L����Lxe򑫂�`��|>�,���c�Zr!�� ���D؃��7�� �T�����Z���L��1��HF��PY�'�;�r=.sA��_-�)�p�˾uI��` p�h6�T�ש��.��� �k���3�S��k ��7W�>e�s���u�Ð�%������ >��䄟��vC#\��ërC�2_�m/F��/����z�j��R�1��6	W$UX���ƣ1��3����/ ��,�e�p�:��';�/���h�dÆ�P����4�ͯH�x��zj]l�����Q�f�uU��"�q�:@�<������k���d��Ķ��&�3��X�q��q�h��lve.;,���Q���.t���u4�p4z�-[�Fi6�	�"������:�Z-1��P(P2��Z������[�e�4]|��-&�����#�!5������ �i3�$��z��[&���2�|����	 �[م���˓h>� ���YL�G�?�3�.h]���~HWa��V�s�J�����t:�%M-�̅�:�H�6�m`���#W��5V��Q�Qx���P~m�"K7�	|<�F#�f�w���>���y���z���\����2�͊��� @w8R6�}1qpq�?-��}RUad��:T�ӵ��!~�� & ��98��q�3�J����׶jp���TX%3	:�ΕQQ������0���a����F�L�����>���9�%@+�C���c>��`8�f�I�F�:��8Hq .b��h�i6��M�շy��JC8&
��!r&͊�ph	�A/�W��w���rPR��=�Z`9�ʂ)��Bq]1!����d,��\skbmuX�ibܑ�`���BAL5���?''�\�J�<fԔd�&f� 2��Y�	f�PH�c!��R$p�������D⦫L�q?0%K:ͼ�F,�xV]����(`�%��ItB���
���}�`���<i�F��ˋ���6 �����?���W_}%|�1=�>�J�d 
	ɒ�A,�Ų�^��4���צ��j$���s�J��<�ѵ%�..W�u=�L6F�UY9(��s�eK-]v�WJ�2rTu�� ������A?l�>�+i^+AU�R)��������!�{Í�;�u�]��ā��� ��e�l�,p�S�A�:��a�w�\.�gԭ��K�I_V#�F�$;t�����'X�ڷ��:�i�<�2�d2I���b
�.[n����>@:��A<G�ѕc2> .l��j|?p9�:�m&�=���	ܪ�[�g�܈�np���'�a]!6��H��Ľ���w"�Hy0P"��l6+�5Hy�Ƨr�.�\Թ��6q��)pf�e$�.v��{~}�M�]���a�+�{�L n&F�1���yO*�D�U�	r��;�r�&�<�������9��:=���p8\Ã �Y;�1��B� @�c�,�.!4�qT�$    IDAT^:�LT��h�E�p��_\s�aA�R��_M]�G��'�R6��|>�$30%���+&p�n�h�T�3�ܲL>��q�����F�A�^O\��Rb�����E��pf�*ry�*4٧z���IL�T�d?k~����Sx<�6�b_*�ZJr��v��6��d�_+n�ݞ`�E<�l6+���p�0^{8.y
sͭ�"`���p��W�D�� ��J�_}�뙨�ݼ1\&vdP���燱1�u�*UeM��ѡ&;�ui�L,�*S�������v��|�,X>�]���c4� ���S��Es�<�@�;���������#;��
���aο�:Б�~6�]y������YL��~b�k,1�A�k���D��١QGeo>�M]�x�*�H�x����R�٤v�M�~_0����!����9�j5j�.~nUͳK)Qu(�%F����芞YN��4:��9�_�4>��I�V]-7:�?��1JĲ����������)��&mll�999��ڵk��L���\�V�t�]1�,��rƿs	b���׹-��\�r9W֑�� ��N߄�L�+g.��z�fa	tو��5��lsc�x�l ����p8M (�Ђy����X��~���(��!ID��J�ĵ�t:� �~�4���5�%�C�O��$c�;�����4���Z���2MG�ץW7=׵ӝ7?��.� |��3�M�S*�"Ȥ5ս���+�
��u��ݥ��M��9���a�h�ף�p >��rm^�&p�Y|�oCW0$�H�F�G���REtu�q�*�]���Z�L&�d3�}�x��3�xM$x�ł��'���)�Yy8�:��`p���;����D���#��gd�|�r�I�>�x�	N�7mɳ*�^_�9�$5[uS��do� ���Օ�֑�.�M@m:��4��f��[�6�e>8X�T�ߧ�pD��T|�&QNB�K��v��Z��������B B�Q��&"�x,N�d��ɤ ��`�늒?4T��~A]	ʔ�q�����m��3��N��TI�id���:��K��}�3z��yل�Uh]A��3��Ľ�B����C�7��.{�uX�:r����U/���U�sܟ�� *��%����^�cb�d��=��M��Bkȕ	{�	|�Ѡj�J�h�������Y�R�N�#��
 ]��\:���X�y�ɇ�eŏ����[�yބ��T;\�\\���np���L5EK5�Ӥ4���.���\�����Lu#l6�L¥��;�e�~�sS��řZp�wlN�&�wj��g[[[�EG,k���� �2�qd�T�"��40 !��B!�&���O7��
����Z1���hD�A_c-�2Ɍ-X	�ٻ�K�:A@���A��b�*"�^O�~T��T�Ώ��*k@���:/��々NI
�6�L���<e2J�R4���U*�zUͰWFT Q��b�Mgʵ�b��.p�K�L�k����]��l,/�c� Ԣ8��)��P&�gɂD�x�Z�J�B���H�ј��O$�-;�@�Ǡ�\�kV��r.\�/
�i�`SdZ�M�j�I~�g��Q�Q��/�<�!p+OV�M>ҕ~t�DMۺm�TS��f�a�rɼU�%x鉈�l�0����P��
zB�K�ru(��`@��"X���V�5�&�LU��Cj4T�ը�j����;��e�Oggg�l6���
�l��6fF���J>�A	��\
&�-
�(	1���7������s�6[Cލ�-�Z����%?\/�Q,[�6s�0L��\9��6y�ր��T�"`m���X<�"�hJ��T,i{{�666D��i ��s�H�LkC������uf��W���C��_�^
�0�rN���R��~er�s����F�������X��8��1᥾X,��l��yw���˯�y��g���z�;�FCT���ǂ0���'8� v�oc�\b�r�O's����OL>�*�(��K�v]�b��o��*�+�M]�(O@ѡr۸O�uaEVaI\��lZ_�hPW|�5�����˃�3����s1��C��6�F#a����l6)��o�A�l��(5���?~|���	k04��f0�N&�B��N������P�d���9�z=����n�Ž���l`ƴ�]�wu��>��<
��ʲ��1E7E�L�ʥaE0U�L?�>>��xL�NG���~��<ZLK.���M��-�	�`$�G�-I {�/hnʹ��$
h��g{�6ѥ	�d�fKL�(�k�3���N��nK@�$m~˽���?���𤗻���hX�`vy��2�ͨZ����|vv�!��:��������ǝNg�R�!�9����{�U��hT����1�E焈	d����!�ث�!��e���\Y�$A�~���K�<]IǄ�m��L��) ��t��ߡ����	�.az���ᓑL�>|�,I&�K~�բJ�B�H�(5���ߙN�ed��~)�G"�f����(��Ƌ�p(*  d�wbP�x\�kW�����,�-�b�E��`���+O�����u=�ue+k�oQ%?��vq��3�:��<�k��W��	�M rb��慩cVm�A�j�k�`P��V^T9��]/�S��%K�t����_u��VU	
jmI���1��w�VvH���`�~���8�J%�V����O�����~��O�_�r �V�}��t�*�
qF@�I����+߇%��|�44����+�r�~q����y��yW�Wu>��᫃T M����<��z�T>����=1S�3uѺ4���a���Ἤ���fɋx4�k�Z-���w�������WZ���ɓ	�F(����S,���M���"���n��p�nW�`��h4D�1 ��t��~6����LTMa q�x��^���(Ib��^3
���t��䶎� ��TTA � S\�@#	Mr�������Uq�/@ԕ��T�AW�������ui��5F���D  ��dp]EB��Y_�ؾ����Ϝ�C+�s�M�Q� q��i*��L���r4�����|9�;r,�g����={F���Bc�.@.����!'`���E�p�n=���i�Z%A�U2T��b3�統ȞˇS	SI(H��,C�`�f6�^�t��̐��Sm����1��v�fJf9�t�,�	E�\���<�b1�N��L&�s&�I��鼲�&"��������7wŵ��2�NS<������>\����sj��bD/�$C쇵3e߶�&���d�94B�X����orѓ�b����e [���B)7�JQ�P�\.'|.9�%�?�����*������KɣVU�F�����*V���u��x>���O��b&�% �^u��X']�Ϻ�=�ȌF#qM����'3"yŽ@i���|N�BAh�)�N���o{�����+3���}8�����k���[���Z��0����A�����ԏT����E�*��U,�\ާ|>z�UeE�MPILlTF�ԑ�Z�ӍL�1�~�At���>yJ.��@�3�D"! 0���]�ۏ?��G?��+rONN��v���b�7�)�NP�@?C���N�&�	e2q���z=a�˘ L�j��@����� |-ֆ�?���Ж��诀)r�l�s!Q}.S����l��*�>4��tZ��l��W���[9��,m\c>!����{�`q�U��N�}\���/ p��D�~\'A��yȁn��:?����~q["ə�T*�t��ȧZr�����%�p���t:M�|�NNN��h�www?y���G������ثV����΄��$�c��g3Fg��%���2X�����n�9]����G��a?=S�LC�S���3u��6M��okfxY��*s�]2tμ�O���4\�`_�K�Ќ��h0�4��x\�t:��qw����V���j5�=,��x8����n���ТaD�ӡ�lF[[[t��-�f�4�L��nS�Rݳh�	�\4T*������\���q�@ם��[�s�����#��@Sc��p��
�6?�e�Jy�*�P؃�pU=�9��5ڭ���3���$f��GG�Q�"Q�Ře�_ 8��W%��L�u�I��c~Z���2|�8���͇_6*X�� ���!�`(����P(��r�ONNN~�C�n��ɓr�V����l������h���2H|���{�G%�r&N:��8:[>"�p�Tk�Y�5��T�L8~V�$t� W.Q����r�|@Ws9�����g"��Ⱦ�{��ș��bA�~��ө`(c�� l��8Z��^6HM^5p[����������\4PD�Q��ܤ|>/��&���R�ݦT*E;;;���!,w��0����_��vww��h�Ç���������A�2�o�(^j��h&��� I2�`�׺R���Ӻʼ�&*���בH<q���Lʕ<O5�Wu=]|�M�����*����O�LW����FMs��
؍��@2���s��% \���r �X�  הL��F��n� {I>�	vwМ�q>��k���R<�t:M�������������?h�[�����l�=}���ժ`b!����� ��vX�8c1����5?���j��R�נl��6eÔ��Z��g$�K�pi0���ܧ:0\<u��(����U%*?����Q�B��`9��G��<��ͦh ���D>�����|���]��٫ p�����n�|vv&�O�ӡX,&|p�q��i��ڢk׮����(+�z=�u��J%�v���i���N����V�:@gg��*�������gne9�N+���~l{��yl�i\X1c�u�8�F#�v���7
�|"��R�7M��~����\-�v�6�P~��&�k�χ� z01
I:���lY3,7U	7/J���
��;x� U�g�Vۆ��J�A���F#j�ZK25��qi��y"ч$a8R>����h���!�Z-���i��ަ~�O�|��F������}���pR��>�l�ٳg������h,Ux�,ax�UL|����.��ف��_�:q[��%>���3��蚡]�ZT.9���:{��$3[C�_q�i<�ɴ]G������6vۼu?�k'�|q0��@��e\K�cI��R��������+����_�wzzz�ٳg�܆d ��w��b1�v��R)��rT,��ݥ�`@�l������q�v��`��
~�6���\0�ϩ��.�62ki�Zp�ץ��M�T��\#T��#���J�"�&(�^Ȗ_\߉k/{��2��%��m<q�� �T�x�ʘ�>��c�?@�d2Y�X¿��Ƴ��'�KR���-�S��V��2H�)�:r�6�Ǐ�����F�A�ł2�e�Y�����5ǄGX���7��S"�6{`���8mllP(�Ǐ�d2)���۟�����G�������ӟ�>y������!y�G�Ba)F���v�D�2���s����҈oU#$g�e+<[�e��6��B0p�C/\��\i]2痽55��(�f�A�EP�_]�\�����=�o����q�8 �P*��<���f�I���DD��<yr��w���6����rvv�wzz*�ء�b!X
��l6K�bQ���ᰰ�I&����8�z�Nϟ?���s�|� E~�m�R�}����:J$�҆��(_r�jP�Df)M�����
���
�����f�XP�բf�)�>���eI�PD�Q��Şr�^�:�UeǛ]��9C���eN���]��1���剸Jc�R怘�%'��ݸi�+ ଷ�����dw�.�U%Qa@���o8R����n2�P,�~�O��x)~��B!1�����L&����'�����\.�ϐJ��A�V�����퓓��G�Q,�B� �TYgi�����
�䨂���y����@6�\���um��E�c���Qɯ��)���N����
�ubAf4���M-������v�]�����%� �< c���j5J���d2�ɳg�~��o���TGGG{�f���㽇�|>�l6+ ���С�J%J������^�]m,�hp�-t�ۥ��3:>>�z�~e�| �������% .������f�t8���M��U�F�q��T�a�T�s�Fy�>g���ؙ����-D��l4�f�:\,����y�� Q�Kd¤I����z���\���/����Mӹ�&y�޿�h:?\���,W���d2K�ceg���*�f3���ԟ���<*�4�(	/J�u�s���6u�]:>>��t�w���O���?~�w�w�[�[��U�������tttD�\N�������L4���nWT�dG0�|�4���	���:�x���wq��ItU�Hk+��
 u��ݰdӈ^��6(˫���:����F�n�K�DB���f� t��DF��t��������d2�M?���Z��w~~������W_}E�^���$M�SD��j�Z"�Ƶ���B4�^�S$�B�@���φ����zT��^�0Ȁ֦-r��N�|�?�8�A��EA��$yM'j+�����nM���kw${���f�\���d7�q
bMqS勌��q���1������Ye6�x,.F��2��l�e�{V���\�$@�Á�������n["*?wU�N�(�d��1��^�S,�b�(p}�N9�R$��b.&8B�����k�ye2
�BtrrB�f�B��}����{;;;�nnn~oΒG��+�����������Y��Ɔ�#C��=�Ѽ�feH�&�� �`ve�:޸���g
�w�
�����2�.�\UT=��xM�1�]�L�/{�:��~�Nw�jR�?g'3������E@��A���j4����͛�z��鿦��{����{�{||��n�?�T*{>n�HDh��h<��-��R)�P�B���f)��PԋR�ߧf�I'''T�T��{Q�S9��a�\J<\&�A ]���=�(^�O.U ��c���{eKU�i�u����?��9���,a��D(��hi��-gz1Hc0��ˈ� ���r�
;��m9oL��i4Q�ѠJ�B�N��X"#V�A��$���A9�ЃӍ��ׇ{��vN��S�p[�NPp������ ��������b�r��������,�DD�s,�Pb
"�%o�B,I��4�ٳg�����p�<������G?�����l�_|�wvv������7�|C�N���,��iAA����d4pc
b2��L&��x�s�S�1�?t��V�Б�~��-��,�<?J�b�lf!�w�������\�y݁-��E�*`sBc} f��Ց��s:����1E��666> �;�J���g�{||��j�>�V�{���4{�Q�>��	��p8��L�L�|6�t:M�l��٬H����>���ѣG������h4�eHW��WTo;�Q2��1I���rrp"�Q�����V�p�r�-���N[c�h���h<�h,*X.μp}v�ӡV�E�z�:��������=D8;���R����)�r9�� �4'�d2�z�N'''tzzJ���4�@����e-�Z��w�Đ?6��l:[b� ������e�n�r���r�aZ.NE�ʁ�YTF�5�M������h{{�2��r9�v��#k?�>� 0� �|��h4J���4�N�^������uz�w����?���~w/�N����;=K���ʣ��N�Z����ݩT*{_�5�Z-J�Ӕ����<!� #;S2�{��R�$ r�ӡJ�"K�������<����z6�ړ�j1�������6�6MASi��}sV�����ʈ���� 0���b1J$��v/��ˉU�LF,��"�D`���p�z�=|����)�����}o�
'''{�^����.i�u�g"g󙘱l>��|6�[�n�����yJ&�4�L�V����1}�����W_���xm�M� 
�^��H����|ҙ\��5���W���_۠�7W�    IDAT\��v�- �h4Z*��\g蜻�.5�����f���A�`U#/`G�=}����"e�YJ�R��f�C�t:�p$,�L{�5����n��ŝ��b$u̡���4����h��DP�Y^�b����Y���*V�/ɢ��F�#a_��l6�V�E�j���<��if�.�������.��H�@�L&A �j6����_S��(���r.����_������ƍ/�Ly���^������|���NOO�Z���y���H4�!��C��)�J�3%�P���ʅB����E��d"�����F
B��������]0�k��� �ɡ'��_Sk�C�5��� ��Va�U?�uV.vc.@X��T cW�(����ek���B܎���+������?��_www����~o��Ç�*��'�Fc�ɓ'�l6E0����
�K�^�ȩV�Dt�C�!�J���lR�V�o���<x@ϟ?�~�/��G�\���v�\np��4s��r��y�8�0>��ue?0���;
���{5h�Q]G���y�=y�n޼I�\��z�+M9`{�ѳgϨR�P��`B���2��s��d�ᐞ<y"<8��0���{�d<Sԋ�����m:;;�j�J�fS����֮)ʬ���_ �H��f)U�i>�ӂ.��x^m�{h���lv_��� �ka��W�t������X,F�RIT�d�x�~� `��H$D�����i{{��:>>���cz��w˱X��o?z��^,�t��̇����px��lN����t�ݽ�����>}J�x\ئ��i�$��s˵��9M���!
�I��v�Z���j	Om���9��M�D�^\'��`�xgld��-n!^�U�}��y]c��i]�L�LC���y�h ��L�;��x	>�L��<o:������n�Q�������i<��>��f~�������[[[5�[������ó������{GGG���X�E�:� ���!��h4���3�4�F�j�Jtpp@�jUH�Q7gtV�.@��B!�Q$�4����Ć�Y�YA�W�TK~�0ҦϋCf��|�7��F#z��Т�f3z뭷(��S6��a�Ѡ����/�/��gϞ���t\�kL�L%���pH��@��rT(��A@�Z�����ѣGtttD�~_4�֚�]u��RHRiXQE�k��G� 1�c4-1�<a3EU2b*y��.��&Y��
�#�x��5� l��di�C�T�L&#��0??�� ���d�J�LFH�@�q�/��J�r�P({�w������B���;ＳҙR����z�����۽^��h4�QoP�٠��sai�F��&�J�9�@� ����
V����l>2�-�H(���x.�����.-�)��j��@W�m�돎t�Vy��oWݡ_�����O�J����Au'��ZM'���`0X:��hA >� �,L&��c*
�7n����??x�ࣟ��'�y���_�W�V?{GGGtxx(��Ac� �J���>���F��F#:??�'O��p8�X,F�F�����,�p�x�D���!��0G¢�7���'[�r��>��B��x�xOn��b�UzW�m�����V��
�B��M$�V��~�m��ަ�dB'''txxH�?������m�ޮz �(p��v�- ��Ύ�D�f3!�x��9=|��NOOi0X��m���6�F%�RP�uǟÙD�g��ԹN�;�an��t�ӟ�$b0��sccC�5${ �:���=:��ZT
��,%	*�J������^�S4�����7ʝN���{��z���4�%yB
&��K�t����;�Ѩ���Sz��)�Z-�s��6��V�	��."ܯq�5�W�����a*�<��}j���l6�^�&�!W�\c�KC���~W��c��h�E���L�\�஛�^�E	���_'Cl*Q�f�1�6#8����E9�����~>[�O��{�@���t:T*��r������e�ٕ3o����I��nX�Tn7��=x���iJ$�v:�Y�A�L>�����j	M������0#7 W�O��C[yI6���% �^�`�d�ˁO|8h� ���X�p�� ��/� Uy�4X�y��������7ޠ�xL�~�-=}�����[:>>(:����npk
��74A&�I��b�n��X,��yܞ����ᡘr%�o�ˊ�J�A��gd�X"�/ L�����$Q�%�c:�mZn]���;x�(����.�r9a��}<�����ϵ��b
b.�#h�*�JK���'O(��c�X~�h����L8���v��k6���$!�H�����\�����A��j(	�M>
��rNj�ZB������%cȵ�U��5��{dy�*�u�ky/�û�Yב�Asl�G�1]S�i1�L�m:h����:Q(����D.���"��B� �A�� #c-
��x\�v����⋻�l6�L&#������Y�V���px�^�O������������������V���ɥН-J�RK%7.d���E"�nc޸�:�Ĵm�Z��H��9��D"��u�=\���;���p�~ cY�˟�b�t����B�}�5L���(<pc?�rqxxH׮]��dBhR��t:-:�m��ˬu�ѱv�DB0Ph�|��9�r9J&��j�����"���t�t��I~�c`]?��}��.{�"����  C�]7%�&�?�ɏ�\��҄�"*;?�&�yH��#H .�����񄳭 ����H>��B�@�l�&����T���%
����`}#� �AV�D��p�i�D$�n p������Jp~B{��)����W�'S����!���L��d���鮗�E��Ig:�_F��.Bf���R��YȘ ��ߘ`����8�0��D)��	�,�7� �`����bA�Z�z��r�r.�+�E�����>x���x<�����}�J�R�N�w&�ɤ^��i���J�"����#���c���K>o|@ ��f���@�/$���Ri6�Q�ۣ��O�~O� ������X5�V�_8��i��_� �D$X^0���<�e;Hx$3٪Nx?+K-�>v�T�q����Cz0����j5z��(����=�m�v~�z�`Κcosm��ё8|T�c"���Jn\��U�<*�?W4���2|	*,` ��'��A��_+#3e�Os�v��YV�[N1nR�|>/Q�CO^ۼD�؀u��OJ�g�b$���6�J%���.��C,�D"�
���)�d@Lb���x.�#����7iB��sc</�����^��w�d�����T*�v�"�b�(cb��!&~������nW�[}y�*�?�������A��\�7�ar�htu�T��vent��b�U����u:�#-�J���>h��,{y*�W���J�`0�+�����&�r�r&�)������߿�L&�ܶJ���f��t懇�w��yR��ϟ�r�|>��t:-F%6���H$���l��~�O��
�mllP*��P(D�fSؿp� �fA@u]֢�gd��Jʀ��A��8����7�q�w��d
6p��>��ua��h�e��5�8���v�<^�� t���3�)�挿�9�$2n���`��6�
6���iz�z0��h2��h	 ��枮&�:�^׹��9M E�\�H���7N����@ )Ryb��=�砱��1���f��h����S'q���P�3$H O�W��F"��g���3������X삅�d)�E�R������A��w�!.���B���3��Tz K(]_SEh�8)�dT6Y����[ۆ7}8�Ւ��B՘�
w1)_��W�U�<�|�5ʖ0b"�ew+��G��r�*^���]��p#��@9�N�3�L�4��	EUp��b�������ai����A��1�(s�f3�l�rs�V��dB�f�������Q$�\>�����f��a���Gvc;<]?��"/롼��G�J*�Q�{������?��{E9�W������'S�QW�o|�|��[��q��5U��C���s��@#(��s8���wadL/�&]�	��~�W�D\H�&c�o`oy?��� ֏UX�FgSS�n8�i��������R��p(H��� "�%����Ǩ�$��+�7�ϋ
[�ݦj�J�F��鴰x���?��r�W�3���c_ ��\wx_O�^��,�����f������!�����ٙ�>?�e�;?ɞK�˖ۘ�u�]��P#�՗I���d�].�92(�TV��
��3�E�ua0\�K�e�
WM�ᇾ�^����X*��T*Q�P�\6G�TRБH�R���%�C ��D�L����L�ٌNOO�˳zX���q0��N�C��Q>�_
t���nX~mnnR�Pe(��"���-�G"�N�Sj�ۂ�A��yȯ�	���I .�pޘ�
F���:p[1�O�b�\A�jOؚ+M��5I6iU`BN�<�4�J��q�б~���r��ʚN�Ӌ���ƪ"��L3X:��D"A�łr�� H�YA�ĵ�.HI�˹d#Q�{Q�i�*?�5��
<דW�z�U�U��r���%4hA��}��d����"6��
��[�CM�v�KL�����A�CcY����P(�����"F�QA�@��I�M�'�ZsssSr�����K[[[B�T|�'TɽK��GV��My-�Z���6y �/\c�(��&���]^��(���ǝ����h$ ��CޥiL�ErE�A�t9��=h�|f���耳|`@k��O�!Lg��+�R�\���6,ؔ|�`����` ��9�k����t�<y74ώ/�_q]�~y�,�\�ө��|��E��0�FND�⚶Z-1��~:�R�٤n�+��d�~tP��e� [4ȝ��h��KT��|$�m��ua��.Ur��oRlbmɩjX�qr7	�Y�$"]Õ6E~�8�u�����tX����e�����R��ޢ�n��"�J�8Ɓ .b��.�������:M�gk�sa�T��(�����>U�U����М�x�fJ^�B|A_�x<���"�H&�"6q�H ���<)��$ö"N@pq�\~ޱ*��>���b>X�1Q$�?��O�R�������dc~� �TT5.�'��e|�dǔD٤`~&Y���޷pQ�N�wJ�RY�O�l��*��������D��]��hbvU�3u0���(lv�l���"��
P�@��Csŭ^0���E�'/1r+/ _l`�\B;�K��%���pH�Rbz��q]�Дp+3wA%'~����*ݷ��"���_L�eJ���0�L�mO�)�����ⷒdJ�ul�M��R�4 A�?T�Y��u1J�t_�9�X���|	)4��؋! �����1F���dƖ_c�^��ҽ����o6����O��nܸA�BA�o^��A���,�F �x3&��t��%-���`��AV�l��Μ�r9o���t�����D"���!��|>Mχ�����:==#ґ �L��'ݺ-9�]:\s]��\��u�=~�Q������:� Me�b���ʒ�:��f�.�s�+"/VlT4u�]�T*��A��� L�����L�ȗ�I�0���p8>	�˵u��; �P��̒��R��f3���tZdޞ�Q.�[�ƃl�e/���g�2�_͸kӀ�}��v���ؘ���]~���Ac��q��	\b�𙘋 U/����*	��V�)�=���p�|UI�<ϣ�l.hL�J����D�Mp�q���Pꚅ�'�#�+7�)]����r-�jT)677����d2�4�rHC�΀��p+��  %�x]$3�8$�%���~p�xeq����@�#"!UH&�4��+�l6ECY�X�X,F��L�����t||L�J��� PB���B��舘�H�Ql,����>�6���u��p�T	]�O�yT�!��?�+a�\P����u�����V�i�C�+����Z�U�U~�moo�.p^�A��� �`��~��(�pJ���|���a�ȃ��	�;����U�Uj6�"#Ǹ]D^.����e�1�~����������/I�%]�h[̍�˦I��A��iԩn���M���U֋`kj35���.~P���\��� 2������=#J�|�׆��u�v�'��Tٴ��H�u�_ՙ�{��q	���-�k8�3����t* .hb���k ـތd2)dfܛ�g��4HB��-_��J?�{Jp�A+y�PnM��h1_P�ۥ��Sz��	�������|HT,�gl�_�K�:�Ϗ��oe�4e���v� �H��^� W�l؂���k�
rد��><\l��ex�9�Q,���C`�8D �M��,1�,�l/��'cA%k��,v@8�`{��2v����^�'\  �P�
W=tV5�6�,����O:B�тh>��t��'D!%ۤ���<�N�jc!���.AZ5}h;WFD�R�Ⱛ���V�C���~��O�n��� N`��>>Ek>��l:��492%D~֜��l�����U@��|ČJ���#���C��۰s�v�-�g �[x�L����#r� s���~}x�)�X,��� �h�C)�:p��u �ǅ�C$�8/D�z�NNN����D�4�H,9w�AI.#gm�)����"32)/�2���um�*�"���T�ٯ� vy�u��m��V)b�$�|��D��ή_�.\��(%	��B�
Cl^f@p�Lϖ f����8D~�9k�[B�U�"���׎�b�VZU\c|V0�|N8v��S��R�]%�r͚y�,�2�A�k�C�Bt��r�ٕF�W�e��ʄ\*)6�� ��� 3X�~�Ϋ4��L��
�� ��CR�'4i�m�;7 n�8��$�o6��d:�o^Ibb�\XlU2���gߘJ��$n�E8<<� ��	7�Z�F�N�F�� �D�$?C�J�8g���r+.�呹 �x?��D<���8L�� ���t���p`@2����-��3�L�rFT�V� $�]G�oж�U'��!
m.)~�>Y�N�iS"�㒪2���^�u�� z�<H��~�Mז�<�[��Q�TD��ƍT*�(�NS&�Y��D&�G�r�/[r���t�"�?>� ���닉88��}o�����9����v�j�5�MQfR� ���k͕�S1=�q�b�$p����d)3%�� ~5Z&;/�ɨߑ���c��vm(����Z����4�%f\>4tB�6?ȁ)� .<�*��!$�镡%6�æO�ug������ � �۵/��=��Y��h4J�l���$mllP:��J�"�P!{�Y��l&��0��� d��B6��q�~�/������ �xH( @A�b1��١P(D�j��ݮ��X�677)���h4���z����/��R����	`~q֨l��]�L צey�YW��
SE^v��}�Va~z����v�����X�e#�9�L�6��K�`�_'[bk������ʯ�YTn����
���"�������% .�O�F�܂�` %��rv�7�!Xd�9pZ@� ��GG*���%o@�>D����Toԩ^��F3�|�-���k����O%�80���A������6X ��cڕu0iQm]�6oYݵ3�O�a2���{}Wى���CU�����$���x]�<�i�u�@9��DR����FWhl9KëA�3�N�ٍ�`[�:kFU������i�G6��*�@���Sr4�9>>q���ߧB�@�|^�y�z�%��f�^��t:-`��^A2��dR1�'�H�v�-���$mmm����(��$Λb�H��ۂ���14�����c�V���W_џ��g�T*K$�p�������A��ت*��ΦD�%.��o\��utr�XU������+�Y~�"eb����L���Z�k�������X�|x.����ݣ(���}:<<�n�K�f���"��)JgҴ��I�tZx#��d<    IDAT�z�%oI@\���aB��f)�J�`Ǜ�p��F"ј���?+�̀@2���7FI	�%1H5��&�u1�����X�$E�:�FM�����Ⱦ�(�A�̯?�����.��`�6&\���.�@�0��#O�L�Y���Ֆ���!���,��67��]㝬�EeH�<�	+�x\T�P�F��l��+L��̶��d�%3�W��,R����=�z(�N>�gbq�ӡo��FV�u��b1����X���R�j�x<�|>O�B�2�̒����^�B�@�R��}�]��ަ�|N�v[�4�t:4�iww�677��wޥt&M�~�NNN����t~~N�DB��hr�$��hP�ZױR�P�Z�/���>|H�FC45�3���2{�7IW5����c�]�ZU�grq�<7�@�%Gug&'���
���A��w��?��*�!��]_��t�Kl@0z\0�q���9mll�͛7i{{�vvv(�S�Ѡ��3�v�"��<|�H
��6J8�cM`�����ہ�� ���l5>3�
C��d�`�9���~~7�	ܚ�?��n�[�ȇ��ՕG�")��R��!���S�{ޯe����:~�Vz��Tl�j����J�H&�|�`�`��\ʛ(��=��m��5M��[ž��� ��e��شղV��Yf6�����1
b���r��R�I  #�!W�t:������01lss��~�m�q���g?�[�nQ�ۥ��}����"�'	�(n�[o�E7nܠ�|N�N�髯��z�.�_�� ���y||L_~��`dONN�Z�^9@��l��\*�&l�G����f.����R��}>yB��sە�S%�Wܠ ��`�~�M���&⦒�KS�ld���� � ��h4J�b�vvvD�v0 �����U0��XG��U��s`3� �Y��b�l0 ,j����Iן�`U_U���T����:ȹ-ܜm��[>��
_\��Y� ��U���ت�F�������f�Z	0^������8mk�t�^9�)$��\g� .oT�/ّE7~�T����k���``]I��5��@��F��_!�d2�{��#�L��卮�[(�X,R8�F�A�Z�j��8�@����[��[o	�Z^���v[��� �x��R�$�|k{��`���*�z=�v��B��j�h2��5��\8��� �I�~ٺ�C[5K�Vu�+�*��y �~^)u!�\�}�=�zh�>w,�-�����د+��������= �m��[��3��	p��(��.y󑆳ٌ677ikkK8�nW4@���2t��r)L�a7����
�(�H,�/o4�h����pږ���UJ*��N��0��k�����.�pF� ]T� (��i����5e0亇]��X��Z�?�n������"T����J�Ja�=�4�/��������*���QӅ�2�\[�Ε�]���R)T�C�q`21�h���R��{�W�N���g( t<S�T��������R2���` d+�l6)�J-�pGE�%�x�r���yZ,tvvF����7ݎ�:�Fw�sa"� eR�HK���n����}��m���D��8"1O���?�8�
�13�z}��e�(Te�<Î;v4J�prr���c�� �|�)�H��#��R�K���O>�ȵ�ز�q	g��+�d�U�z~�������n5�T���X�+����a����l�����r�AZ���#�l�!��c��龜2KKK������&*����r�J��fS������h(сD�oޤ�\���A�`Z,�a����ڶ�mt�]�,��W[��V�>���������v\K���&ֆ�u�.:���P�F ��|5�!�|X���&�Iw���O{m�k����i��S��Բà��򟻴�>��6�Pm�)Ir_q9(�X5�o<�F�I{4�T�A��TtU��Q��Q�T���Ғ��P�01����������
������cܿ�^���x��F�VWWQ.�U�V�F#�ٳgh�ۨ�j�8;;Su#�v[���^O��%v6��) �I:k��5��z���T��J7�hd��`Qjy�X���ş� �(�@��E�!���>�٦�+I65
Pu�����M�y� ]Z���/��!��d2QU���{p�����S�T5@Yx�d&��@	����"�ĕ���R�M�!C)s W��������t�L&sM*�����%[��'կ��Br�n��IoM�4���>7JǮ(���m:�]l��ں�4[����= ��^����st�-���Id�x!�������}���y#ӽ�Ɔ�e��������
1���~�6�Of���BA`�n���^����^��Z����%��e���c2���� �V���8<<������y�N�w��f��>���x���3�C���);K�ƥ����KE|�R*����|�{!�*��Le�EU�(�wl�5�7����ݧM�-J]A�i����}@9_u�\6�杔�v(�7��K���ŀ�
!\2	n9{G��b�� �Gn�C�E�T 0�N1���v����:�P�r��v[���f�6�F��
���	���X`���!P�[�FD ���	LS�ś�@�H\e\L��gPZ��'f�4�\�K]�>����֮����|�l�Q��˂"��@� "���߇K3�C �X\8���|�����y�0�Zh�1���\��Ov��.1�>2�T>{�o�������gڟ���8Q�X��R����t�b��~����s���ϻ��R�l6��lzMFEM Z���\�r���h�f���Ӌ�"��F="Hv`��YeFe)Cj*:��#�L�mN-�ٌ��]�C��]������v6�E�m�6�
���Ɠ��7�c�!i/Wg�
k�wCo���%�*jyU,L�S\6.Ѹj(-г��r�v��v�XYYQ���rh�Zh�Z����p~0P��p8D��RQq��V,0�ԝ�Xڌ(ҧ���S~ȆF�>Ŏ>�&����=�8�KtQ3R�McCA��1�"\G|���>���)��2yȍW�1:xH�A?�A���ݖ]�U����W|������f���y��복/����t�&�T�z��`�*�epǿW�`�8��B�h%o:�]����iZc��._3rϡ���:�T�,;cf��2�a��ǫW��������R�4��F���d�v����S�ЁWNx�,�_#���&g:?���!����&v2�\�Y#r7��\�~\r"X�2b��N�k�g`�lu�=� \�"��d�mK+��[[�����L��6)}{��>SW�M�p���򻹟!J2�&�Lz�B��V����s\]]a}}�z]E�VKmx��*+�i㣖��^�)/ޕ��޹� y���&��ʥ��(m���q "u�<���g���LKr0���qm�|m�|ے��;h��n��C3#��C�"�l���i�%�!M�u޷��d����]���l�tsY�p�;��&=$i"�>�sF��W�^�S���>]��#o	]g!�y?��������(:7�܁�]pׅ��+�V�)���QV��3�����W�i�膤x�%��^����;�q��xd@�sk�����c8N�p�Y�5Q��
%LsZf�bܨmjy��o��f���P�hק���D�G�6J���l6��t�b"b�xZ�3���p}/]i�� m0��l"�N��SΆ��#f�>_�0��Z�4� ��i0�7��Fm�j�o!ޟQ[���3�(�6��`��
���"i���ǳ7�C�O�i����zH���Q<�I��E���ƅ�O�����o�{��7�B) ����r|
�l���w�۸e��B�<QfB���a!~�Q�CRr8_[2C�u�?��K;��}��qf�KP���Q.��,n6��o�<c<�,s0�m2}0�,��m��9I�����$c�כ�V�Y}�`�� ��\S� �e�d-��QJT7W��	Rl�m� Q"Ӥ�GT��:�|�(q^Ծ�w���(
sfۼI5t �Wn$v	P�EbQ)u�J�T�*]�o回��qF��*M)�&}��v[k�8�ԻY������1���r��鸥kB��e_]Vlq�#���;C���lR[J�W�d����3g���v�8�b �I�JW����vd��&;2��@���H��T*5�"5�Nc2�\.r���EY�>L^�n�I�W�N|���i��{!���� <@����v�Z�MF�:l�O~��BAy�f�Y%��u��9b�� Vf�m�w}���z�I���hj5Οw�ڭPk��M,(IM��������T�7$=�;y|{Ż��]�f���]o�K��t@p �e�^��tE���� �Z�ʍ�����2����\<.��9q1>�r[�Y��G\͍�������t/,3������&����6�5��Cd�Y�j5�J%%��ݮl)dY�����F�����l���:��� XYYQz�B�0W���4^@H'��>�}���Ҧ]�I|H���䋴���%�o�K��\�R�JE5��cjk��ۉ2*0u�aD9�d[⤨}���d� RC���v|2F�?�쩉��?Ԫ�T*�,$/(����.Y�+K7ȉ�\`�F9��Eq��|� ��=�gq�n57��w2�@�ml\ �ֶS��{�Q��x<V�\�JuQ�0�/i�H��A�m�:�ɂ�A�N�專�S�j;�v�����m�x0�A���Hw���H>.}q�|>�ZOߺukN�'��TmKcC��L&��x���K���D�~J{6ӳ���� ���t:���6���������i�y���p�n�;����:�NNNp~~>ז�Gj*�YK�~�m�(���:��^DI��<���W؂�$�ꚂDٷl�j�ْt�Q]іi_�1���ݐ�����{%�%�E P�����5�.]6"N�ۅ�|�i�b_�D�L8�<C+缫�wHgL߹�M*%�s,Х�tQ�2+�}��21��'��3�|��|S����R������m�7�IL,�N0�j�i�F�����tkIF�q*�ـD'�'�3o�3��(���[Ԩlk�R	����������#ܾ}�bQ��ZXJ��%��G������/���۷8<<D��T҇8cD,$��L&�z����޽{��j�V��Kgd)u�\�v*��Rv������U�J�E"���d�$> f6�������g6�U*�b���bQyf���v��Z']�cs����B�.IS�ֺ-2a�(ާQ�l��r9���];;���lA�"5SM�-���}�"�t�X��i��c-�-QXSiZ�\Wi[��-);��C�Jq��xvEZ>���s�G.�,�˾�\�v��P���+�b3w6-`����0o�e����qt�.Yz���Ng<���K��/`w��G�QR3�_�5���kloo ���6�c��a� �������!���)�����W��� �Z�bccw�����6�ݻ��I��=�M
^(���f���t;׊4I�|xx�$,������) �j>�Hs�r:���< ���j���H
��F>�[�=8Ipk�@�*K��@ȸ'M�*�m�Ƌ���C��z/��(�J*�j4j�$�9��>���j���B=lҒ�w�����皲2�웖�)3mQZ���.�1WK`_벤2ipML�+�[X�T�d2�K�
TkUd�X<bru]�l��h�pM^|W�mT܌�+ry]�>'ʵ��y����ҷ�ɍ�ɂ�\����u^�$��M�m�w9����g�p�T*x��!���K<x� �~�)<x���%e#d�W�x��c5�LP�TP��p��-<|����x��vww�l6�N��x�H�Oŝ�r������������Uv�VSR*�� �3�:��4.�R�̽�KW��\^^�/���w�����H�Z'�	r�ܵT�O��V�G�M�JE��~�_*=����Qlw�C��t��W*�L���q~R-�u�n&S7��l���:T�(�q���n.�ё��q������[���}U,�eB��HO|��-�e;�L��|	e�M�3e�]���#,�שּׂ�O���&]���6��8�.�x��O""s�b��M�%	�z=U���Q����t���^�%/�?�Ϳ�"�(�Ft�Y�
ߐ�D�I�1L�KL���/��R��@Bv��,�tA������.�7.����}�6���K����'�|�[�n��x�`Q�u�A �^�}u�Z�ݻw�����+���ȥ������n��L&���-|��W��/��g�����
�Q:��G'������t]�_[[C&����&vvv���[�x����8<<D�ߟ���
R|;����B��j��4�*��an��1怛���s(�#�����4tŞ��4I�-=sݜ�I�lY#�M�k}�@�"��t]��:����L�	��
���NJ�?�%��yls��l"mrW��m���	}���2�]k��8���)�r<Ԫ+J�sQ/W���^��cc�$�A���vIv��*���|B]uAH��;g6$��9��3�U"�^���Y���pM&�t�s8��B7�~V*<z�_}�=z���-���� &�kb�H�!�t�:'�	�ݻ���c�����k?�l$9lmm�ѣG�����?�����T�Ai�J]�ԩ��K6����W�P���VWW������m,--a:����Lu#45O���L�T�)�fH�q������u�>[�,.�uꮦ*6v5��%A���|����l.B6��d�\V( ���e�\]#9�Rv %��9)ͭ���F���Up�Z�Q�t6)�UM���X�5I����4	�0d��ƈ:����fQ�TP*�0,���,�cY����"��&�˙��1.V��y6���I�h��i�r��t:�`0P�q�b��Y�
ӫ�������u����������uTʕ�6�������{%����x�G����R����ĮӜX���/�����?���3�ݻ�L&3'1�A
?�)�1�q�1�%������:����N�qvv���C�PO[���4ϼ�zoʿ�Z�mt��6�>C��&�kkґ$�{?��"�un�*�jH|���y��KN	ԍ�,�(��9�<���Sq�s�X�I�����-[/���f:Cl�>2�9���A�i��L���tLMB&�.%�~�����.M/�!�@�B��Z��t&���+���L��˴1�>Z�$��븨�W]�%S�T�f�4��>�g��ҁd�D���I�n�3�T��v�|c��YL���昮��K�V��Ɔj�N�10�L�)������n4�2���
�V�~_�@tr�Y^�G��X,�Z��/�����O�vvvP�T��vUkR~ӵ�B s�==/�S�6~���y��elll������kww�����:��T���:�]��<��c}�ۛ@�<P%c�j0�S!��K���v\l�M�\Q�bpC�uC^��z*���"�=��6�VKa��$���`���re�ֵ��e�\������,ee���8 u�nhU�)���=na�Mo�������v��T�U�U��˫_�˅Ϧfc��ܨj��`t��>Q��(Dv��̜��0"悊rtQ5gcLL���ͧڷ5�L��J5�
h�l2f7��9s���95}h��s �fE�Y�R��;w��������|��7���A.�SR��)���p�$�]��`:��6� �?��S��e�j5�r94�M\\\(9S�A$�N�et/�M���|���{�[��x%�v�Ig|�	W`qӯнצ���{}�P`OY(��P�)�j�TD�W-:#�b[}�?$���1W��	��3�:�����s �7���4�X-*����B���*нGg���M�s�ϩ��^��7�ɠ�j����l�kq�ΝEl�q��z��5�S��p0*;�x�w�.�8�̽��L&�>��4�<8d�E�R�GM
�áj�+�M��F�`�Ƃ��	ҿ�
q�m-��akk_�5����/���۷�=?*��i�	���o]J�����P��t:UR�T*���    IDAT�۷ocee�j�Z�_��������2钥�-����%\�A
gSԸ-���˺=�t&D�"���X4;�jfdʼsKY���X�l貸�����,��-
��-�[]F��eY�j������&Ɋ�t�$	f8�E��u��E��$���s:�	�f2T�U,--ͱ=��E�*�s�V��t�Z@b��u�f�D�Q6}��!g:	�`�� RhR�ǜy��jB�B����B���6��677Q��Q,1��W�c���y �lNC����kn�FL�h4B�Z�'�|�o����߰��9�-�Ϣ������U*��UQ_���s�"�r9�5�R�(]���)��ϝ��Z�`�L$O�E�.���j����`p,�Z|��7����,���g����&@�t[��Ж����\�y�-�x�K��Y-��:���x%��~,m�.���+W����4�'���2�:a�ǌ2C��m�`�&�JW�<	]�>�0�k�����Ã;:\��L������H�~�Q��\���> .�f���ި:?k��UJ�}�(��ur~-|�r�}E�����s�a�T*a��6r������e��t�4^\J`����NG���H��t:���-|�������Ǐcuu�LFP�����
�2�*���N �?O��i�O�J�1�V�U����j)��/^(�m]*u@`6����Fb�e{i[��^f��6NNN���kַ�sL]�� �ɰ��F�4K,;���Y�Qz��3����|�3I�|��P��s�'�V�1��;��6�fsm�i_�����x�]�7���-#�P�H��	�8��n�ım��ɥ^*��0�Ǔ �%����MQ�8G�����<��B�X|�(��ޔ�|xI�H�M��"|:��1u(4�?�#��g��{����m4�{�.���P*�P�ױ��t�?���3����x�����>�?�_~��fs���ɋ�677��g��믿�_|���- P�W���;�G1��n�v{�%1�2&�-Y�Ei��l�
o�;e�(�ooo��Çh6��t:8<<D�՚��~�&��9F)�S�&$� ��9`�=�V��V��P(�_�¢3�>�Ox�\\\�kQ����)�"pr
Z��|���d�	HL���,iի�<EצϖR�?f���$N�� �Z�ʿg}���.�EE���]@'�&d�@c`���&�Q�M���֑�R��Z���n���nk$7������3��"q�g���d2��C
�
�dq�-pk,�*�]�l�d�T��$�/Ɋ�w�ޡ��bww���X^^��Ғ��������TRn�I2B�������T��x�v�����y����h6�s�ǥ$-������G|��Wx��1677瞋<4xȥRI5_9;;���.//�s$;/޾���\.�j����5���*�G ��$[σ�b����-|����.����fSi�}�\5^)�u�����P(�l�&7���hL��?��`GK�z���EZ��l�L���71U�j�vI�W^r_�ul�®��8}ǟ�>�U۾�;���R�P�y|F�!".Ƚ��7�u��ج\�T� F���K����d2QY:�F�R��Ғ� �Z���T�N�b����>���l�er�0U�/zNIy��LzN#FL�*���0�L�  P:O����rm:�������õ�h����BAu���������۷��g��O>��������#*T#�v8���{{{x��NOO���z������	������y!T�X������|������OQ��0U�l��K�F��Ҭ�Ύ�����S������\=���k�Y^^���>|�;w�X,�{&M�^�'Ks)�ϫ�m$��´��+��>������x����e8t��\�^�~_�v
�}�����M4!�Ώ!�%Xd3_�2�ni�RQ��)EJ�t�l�T�qs�
C��-����#-L�5ӵ�l��v94P���|�`v��榪���B
ޢhtB��}4��n�C���R���_O���L|7���݇X�����ѥOn��!�K�74֔�&����t:E:�F��WQ\�K`���u�.X��߶��MJ���a�IK�<{��������`�|>�z�����kzZ�t�������۷���o��?���D1:4>�m,���	�F#���bccw���ݻw�����l���?����@��;��"Z������_���ׯ�h4����t�{��dP�հ��=�<����z��|����Cruu�Z�l�fGGG8<<T�o��g[��T�El*��
H(УyK5�ٲ�D��t�i ��o���u�LF�\VAj��E�כ�7��d��>�L��؊�] N�2��Ǖ=�	�����,5M�w�,��â;��o���&A��@��*7�K���l61�L����Z��b��t��u"�+�Fl:JG4 J���>ߋ�7���r�G��k9��)r����9`�Q�dt]���0D��q�'Y q����qtt��������ݻx��b�H�G�#Yu��m��˗x��9��bZ�ި���FL&��y�E�E�J%u}�,H���v��o޼���~��������qrr����lr�P���!..����}<x� �JED
p����|>�j��^������|���|�����#q��6\��Z}��I�1!Ƣ3�� �C$��.+TL&��t�̞���.`��!�Ӏ�9���-S����&�9�m�Ԇ��O��R��k>l�M����&��h�v��ڄ��1Z���{�XD�P�K{�Â��u�p����"�$"X�Em�w���LQ�3���%��nhEMi�q�U�
}�|S�o[���áJ]s�.�x���h6����B�۝�ҧ�����\�cç�)������?+����縸���(᪢���F#ܻwkkks�����h4�k�Q(�uKs=G9F��*j�2'q������TJ]5�p9���r�DvӧB�c���h|�Q��I(��t��Űn�ؚ?� ^��c�]犫_�mpI>l*�k�}�u9!E���n��.b"�����=�[�5��&[�f!���֭[���m�כ���[]̊���k�|�ضBW��c���K6r�,�����E��XC��6-�猚dJ\�s��P�s�L4鐉ͥ�� ���f*����J�A@�\.�\.+K.�"�%Sz�,�x�tu 0��/�����<y��-����m�������π�?8i�E�6@~����]�á�N�/2`d�F F�q�U���}�4̭�	����v���ͺ�/ďy����1���"*��%pKk�������|� �F�7�n_4�w��5|�8ә�:]g��ͰO�J؅�C3�qɺ����ZB�T�ç��7l��"ہ/b[�������}�m�IN�Q&�����\1L.����*L�vE&�nbu������HC����>[��7q��C �ƛ .�׉�$拳��ЁyӦ$�t�����ӵ�Cݸ�|���w1�{��r
�):��ruuh���3�g�.�B��P(`yyYiW)� ���@���899����={��������>...�J�P,�s�co
Px����^�|��h��%�ܹ����J%U�E���F����J[�2���k�qR�a���?�|>�B��L:�����y�4��"����Z_Y��-�Y?!�V�S�l��
=3y�-� �I�s�Jʚ
�gvM@�+ـ0_�ZK=Þ��>84�2��������y�Ԛ�jpM�<��h�Fٿuё�m���g�l:�P�"���������*"�����D�4�%h�Ѵ�<:��v-&3�cmC���v7���tv0J:I#J�q�ߟ�K�-8pY|���(�T�KRn����l>5I�e��LY	�C�^G�\V�*��ӴQ���V*���`mm���
x��۶qK�~����|��w���o��?*6�X,^�|W�~������Pٖ?��O������D�T��6F͛��+\^^���{�A�i-��y��-�f��ܸp�ޕ�KmdQ��ۂ֤|�Yd�êE�F�]�L�����w8�%k;��Zn`����4&@��#����4^��ʹ�u#��M5M��n#-\��G�s^�>34���+Q�O1T�7����^�u��䦭b���cevϣ�J��~����E�K-� �$-�����ڂ���"�𼰌k5��${��[e�WWP+A��N-T_m�
6i<{���6��.��!��,F�:P�5�Ɣ�D��p����V����M���zI|qq���}�����T*��1NJ�*���ٳgsR��p�z�>w��f3�Z-�z=t:�{�{{{8<<D��S�p&�K�lsB�%I2���;f�sP I��;�ΐ7���j(>V'�(@ڇ�\�{<KpKsD��b�g
�u-�u��@^W�fcTe���wA�ma�	�����i��In"�\�O��Ȇ�dW5����?�w�,O}R�R��J��|�5S:�F��T�\@�E�I>c����lQk���
�r�b�L�;a���L�i�L���>��)�A�N�� �`8@6�5|\	���@��Jk���5���^�M;����Ņ��TR,��EJ랞���#�뵵5%G(���d28==���)�NNN���+���*�4�a��~}:��#W���\�_z?1�sU���MGAt��Bt|�Τ����&-<��n��,�M��d:���\�\���e=wh&-�鈯3IRD��Z8��)f��nm�}-�f�Dt�%�
�б'��t�n����R�(�Qb���M��b����}.�����.5�Zw�����,�������4jХ�M@�,�K'i�>~o��{�6Z<����V�>�1�Yt � ��<����n�1P�V���B}�)��m˞?��`���C,//+Vvyy�|���8>>F��@����Ņ�S�X�sޕB�n�����k�4�W�c:�p<T��;2��I����S���i��yf¤�I|�9��,�t���%���健,t�9�谄n0�|�}�V�f�Y)�H���]ka��|�F\�����n����i�����t> 7�$����D�*M�ST�UU�M���v����M�7´�ېM(�R���*j���}s�.ל�tǺ͙~���	���7� 7a{�s����<�ҩtA�'Ud��.s�c{�R��M�k%:ȩ�J�XT�*Lk$d��B� b4�����ӧx��-*����T*d24�M�Z-5?hL躸6�|�#oG���p�ӳ�F���w��LM2��rME:�?�a�u�E�]�ߗX��ej� �;�&��ʹ�)׹`���v�ҿ]6U��k[���\J$L�>5%Ir�晔6��KT������к�ߴ����n6�*M&�z��ͩP(�V��C��h��P&��9:�UW4�����3m�3���S�R˿�W�;��ه֩��T:9��J}Y�R�z8����ʒ`�M�GZw�jzP�P��rs�G@���4�mZn�}�Ԡ����̥�e�$��s���:�����'�����XS��84Ǩ�i��R�
N�%/1eT��;�0𲐒��Xt	(&�	f���?�Kկ�3}h�8��M�UJv"��o�:��,�ܒ��|�l(mdP���&A������f�L�VB-)y���8=�|� �d�1_�i��TA�MV�F�]4dK�$M��6}/4tX��H��Z����U�}��-��l(h�{���к.��8p�߰h|9�5�L0�l�ںMIm�o�ʤ�5~�}w܃^�\9�W��e_�A<�S{�n��lVS���z��$'^l&Ǐ����:vvvprr����9�1�g�/C�{�l�RII ��yKh.s1�V��w��q>2�0�N0�N��_���M�l�uRuIvs�KS�Y.QZT�H�ܺ�	����$l��bo}���&����_��]W��H�[�\���6��3��L<��}S*���6�P�՗PNj��IG�J�P)W�/䱴�����v{ή��8���6U��M�*��'�L�����R�TJ�Y���G�nc�U�>�5\z��M.� �aQ9�]ZZ���2�Ţ��N������ԤDw�\>2��n��n�����$&�Ɯ�Q�zq��m����E�pxx�N���y75���}om뉏���f���9�M��|f<�kIz�r�?w	1�\�s]���Q�(�}}��<`3���mkZ�G�>��
w!�� �$��!�s���bN},��,��Q�h��EG��f��n\�����6��Р0���bpM��$R/��v�~CTؘ���q&?O�����Mł�)"}#7��,��Q�[�oW�t@�
�l�}QMѹS����[�� 0��W 
��b�x3>.:6N��6Ϧ�6��lP��k���7�J��j��|>���N$W�l/s�v����r�P��	T$CŖ�Y���t�n�zo�}����:&�	����/]��|�S�5��1�5I��A�#��:`�+��y�J�K�J�	��䌰�]ܤ�m\��rm��q@._�.K�8�n��Y)���i��JY�.�%��6�0]��B�����O�s��6�5���۶W��8�Y��(��L������M3�!��DC�ę6X�e8n��$��v��=ڼ�d;N����샩=Uqs&��y��$@�dz�t������o��näC@�M
H���H VQ��(��m�u��n�����q-
(��qI��� lpy��u�{�rF�{��J�������q||�}	p�3��1��M{����$�~�������;'���|����셵ͯ%�F7��5��KR�.��)�����b��<����[���cշE��9�sR���>����`
rl�o�v�- ӹ���f�`0���]��⊀lzR�I�[��Z��0u�/T�JG�l��>��D��īͥWn�9l�~�\���2��~����M$�K@AV���me����6E�kC��]L�Nv����P��T*�Z��X,��jE����}�z=���N
���񥃜���uT*pK�޼y���S@y!��u��<�A�~_׌�}:[�V�Y��A�ߖe�ϝ7:�@״V�������5���7i�i�	���#�*X�]��u���L�Oq�KF��V�2Y�F�AI�L��mr�y(�����;(u�n�h �"r���b>&�:}zW�l��?������-���j(�˪x�*�e����v0��׺
�E=#��5sp�=pm$�)s�\�4���k��=#�iy��Q�e8�)�Ȣ��$v���@�Nj�n8??G��R�sj',3�����N^�Y*��������^H�.1�����ڨ�l����fS�F��2�}9@m�i-I�̃ L�:oҹ�K�&|\T�|q��P�dH���jY/���@��\����7Hp)>�d�=���-�*/�5U1ݏOѝi�l��n��wh�-I���\�D�u��I0��b��o���g�Z���}>���y�J����ϲ٬j�˵x:'���a�ԄF�q'W��Ǻ�XW�N�T�J�J�r�{ �
S�mHot��]?>�6: ��.X�&�ŗvC<unb�M)bit��t������]lmm!�J�^��P(���Ϥ�K�C����M��y����Mz��Ųl�"u�<8??���NNNppp���K��}����]/4�y������q�7���eҙk���io��=I�k##LMB�Fq\cLghȋgM(������k�zV�+:�a8�j5��9��>���Z�Fe�m��<��z7J�^� �&�6���� 8��h��\�.��~M�4��7����9U�Pf��ju����`� uޖ>Qb�"�P��wc	�ԉ����꺕�F���� ���|N]U�R��}C��ٴo�ŧլ͚����ݻw���Q�T�J��駟��d���������p��-��uU�F/��'��.�~:���h`cc�����j���������&f]p�r\�9��9���=r�9��i�}}�����F	r?v-I�|�    IDATpK��Q��h4Ҧ�C���Oݔ�-�sIF��7�z�퓡�͔�����8!�W6�@��ֵl4=\y@�D9��X�HG�4�I���u�eZ�Q�C��g��bָ�e�TRlg�de�i����A�K�Z0�kBa�G�ip�u���b��$�LM�8!~�L�l�.2��\c��dM��q�ﲚ��Zp������+��e���b}}�rY�bMzg�\�K�S��b���3	ݿ)=J�������&���P��P(���k))��l){ך�{�x��f���<Db�4�r~��O1���Iv�׳���9ר��
f��t�:�7��?�B�J�_�����(����B��L�wa�E'9~ٸ�0]4`[�4D�T��6�eﲗq�{}�������nH����P�BLn���l6C�\F.���Ғ�t2yd��ݔMб��Cħᄫ֕z�E���-<;�����^��/i4}�	�JQ��d����}V��+�N+�w�Z�����9�L����n��l6��������s9v��^\\`ww����T*�N�XYY�cT�- 9�t�CI��|����ϑc��Pxoݷ�����5T�UL�S��������Ĺ��i}H�S�����.V����P�?_�� Z�x&�Y�1`.p��E�xN�f�|��O��SkY]p��0
���e&$���4�9bޥ�ۆ!L�@�No.\e�)����fC��E6G�$�-���jpm�-Md�Dl�l��]����1jJ��	��m���J��0������p8D���h4���*����HGI�T2���죹���0�>]�B*jm�)׆K�]x=�]�V����5�Y>�����,��r��V��wj2�*��
�L��@���l6qyy�n�{�����]�PP^��_�V������9���Q(�y��R����q�ժY��y ��-�͢R�(c��`���K\^^����~_5
1�'�{ ��'��B8���n��B�����ڕ���3�'��r}��� n�,$�`����Ufjy���l���,!)�3���q�	͘&){s�ɶz	_����y�<�Z�"����%
60�èɛ���6��oJⷦ�a}���E�-��,uѾ�
�kr;��bs�y�n��-r]�M��AƷ3�+�F���p�K�@�m�O*�R��I� ��Q"dӖsN��V���d|s��luMDl�Av|��Ih�Zx��*��T�ݻw�s�f�J�J�]�@����N��;�������������N�lWWWsL�ND��dq cJ3=�ir�":���N�R
؎�c�j5�	�D�,�oܴ�E���s(�4�����+�<�{e��Ġ ���㦵]L�OF�ǖ�un&]�eo�ɨ�2�!$`�*���B\kf�>`�tv0��w��������*�k6[�p����.b�L&�ې��f>�K��<Z�:��Jû6�(����)Ի�n�<K�|�.��8r�+����ܵ���W.6D�}�8A$�\���^h5Q�>�P��7o�`0������~_�`K��n��m~�4�|�th��l��ћ��Q�V������E�y��VK������1*ȕE��t3��[:�_iy&�Ţ
�0�I��5ͣ߂�륫[�kDg%�k-8SOz[z.�'	�䎛�w�P�N�渮ʟgt�d� �g������n��"_>�e�N�(;�(B����8LAV�
�ڠ�:� �$&��5}���<�t)Wz�t��C\6. K�K(���/�� ��U���>ѷ�����0�D�R8�ǁ 5͠T�x<V�@zv4ּ���q1��A|Rx7�	�/J�SA�I�-�!nQڞ<i]Ev���C�TB*�B������D�/�@>�G�\F�XD*�Rt.���51dR�"���ƗkZ+�
j�>��d�YT�U,//�ŋ���E��S�R��v] ��d`B	�V�4������e�Ŋ�H����F�}SM�<�e����l6S:[�Z�NMtzݸ.>q���7�9#�4I�&��Mb��@j����ϊ�iɯ1w2$a�b�T�&R��'u�(k_�,4E����&&F��˕"v�CAY��Q�����%�? �L�j�miGSq��В�N��*����Pq�˫��С1���5N���̦�[D��� Wn~�I�R��$ׄ�m4V�����yM�@�x<F���������h`0(����M�j睜t�����%�(��r0(��J��b�'�	��"��:r�����Ou��������`��p�=������)�9-e��T�.�c�S�����^W�A��Ai��R��������Y�<��S�.�d�{��!g����Sa]��٧�9$s���e�� t�a[��l�ţ����$��#MՈ�`Ha��d0Ea��+W!N�h6*c#�8+��J��n!�͠\.���3Yd3Y��-�m�f�b�M�g�S�ɗ=6�"����s9P�6H�g�S��q�	�����@��]��w���N���9(��!�K �g�\1lkP�qJ�v�]�|�R��`�G�a}}�\NNq��+��/��RA!/L���K�Kl�`0Pz���e��y�C%:??���L��ۋO:�/��"PM�M��|I�̻�ـˢ,�|�����I�l�o[?��f4DPpח8g^����s6P�7�.�Mk����6��Π��1C�Q��]k����j������)�01+\%��B�XC�;q:��"���V�H�i�h������P��`�F���p���f��3�7������������Q6W���u�#U	�l�_�2$�ׇ��i-:�}��ܚ��Y��t�v���~�3:<����l[>L�l���o޼�l6C�����9>��S,--�֭[XZZ�{�\�Kl�+��8���zD`�t�@�u���&>��S���)W
h>�>��%�@�����܆���.�ݏ]����mŹ7�	���L7�#�� ڣ( �e1��ֲ�u�V��9�')��)���'� �I��$>2ٻ������]{Ȝ~߀=�&j=�EJ�Jh�$J�T��vu�޴h\����ڴ)��Iu���)H2m<rä�b����j1���n��Z͚*^���˾����w޶1E٤iS!�T*]Ks"b� ɍQ��ں���5/LŦqrY��#��a�ڐu�ajw,P�d2�F���C���������G�a{{[�]^d�En���\Niyi�H��J�M�b�	�\�d[[[x��1������t:
 GI�r�a����3�W��m�dQ�z���إ(`!43#�tk�7p�B:�ޛ�0Gh�q֖���b�e>��)��kFc��t��O��D�2@����Z�W�jwo���<����!Ğ���|&Y�h�@}��+�hKo�f�?����%�V3��
y�	�:ߘ�-�l�V�&V���?tȶ����X��T.�Z��C�t\�ؼr]���9M��6ދ`�谠�����|�����Ln:vϵY�����;NQ�I�Ol:�F�Z����Ţj� S�1&w��Wȁ�l�0�ppp���s�~������;w�m��5��y������VKy�V* @���l6C�^��Ɔ�w�R�~��'���t�R	w��U�n��w�ީ��(���ϔ��f�<��p���_ՙ ��zM
x��\�>�q'S�<CD����t��J��p3B6���[��
����p�x���l�<礍f1��v�d�t�Г ���ys�R���(�Oq�ou�M�c\���2u�
e�t�_�jk��t[�	j�l՟��E.�S�%�br%;�����vD>@�'���&H�<�Q���J�X;뫵���ӱ��>����]�L�O�/�p8T^QZ7��i?DVb�NGu�{���\�Z���j������f�t:��zH�R(�����3�VVVp��]ܾ}�ZMe �� i%��-��amm�T
�N�����z8==5�ٲa�q�	��<��� nPw_t�g�o�e��y�i.ᙀ�p�
�t�ԋ>�%;j;_㶷�鉣Xu�6t��l�	�)��s}Rklcq��ຮ�^Y�>�I-�$>'�>�!�pot��Y7�9���0�eU�h)��d2��/�:�����x���$��B@�]���C�������>i���M�sȼ
ej]��6/P� �XY��� �XC�`��C�];Rb���={�W�^i��l���elll�\.+/i�Р{XZZ�ݻw���#|��g��>
��r���j�h���n�XT��..//q~~������m����I�1�u
d��N�,H����f.J;��a���
o��P�u�$���jzS �$�p�M��#69)KQ+m����ԝ�%K3���m|�s\j~�E/����Qm�j�zMI5l��ob�Ml��K��M��m���2��*
���Jov��kN>숎���-�3~Q=��t�"�#�'�hR��-nL�E��wQ��|�D�]�d�H�Jz@����I�*;gq�E8�L}tx�ADvU�k!��\.��jI��^��w:4�M���������;��f������Kd2,//�\.�T,��i+�_(�In�H��;w�`ggggg��S����������H�y��{������S����W�B;����ξ^�6�}��Ao��5����|�Mx��v�� �����k�r�-�|�
ٛ�����
�n��^_!r[DiJ�0�vO�ժ�]�ɵU̚�ϧ�۵�����Xv�ռ����9��݃s���B�Ao��:ƚ��������(��T�E����=|d��_�5���r9�8L�S\]]�fފ����1����1��:��2ʥ2n��B�ZE�כ��&���^O���:��ױ������9m�dSmY�Ėsm&��Ȫu�o\w�˨�@�"��.� _��w�[. �SH�*X��Tl(u���y�k�I��c��&]'1$��{>�:S��y�ەi����L��F~It����-��o�>��M�5�e�e8��� �br���z?��<_} ��4ŷ��蟭�l.�p�K`�@.�s��o�:6W���e3L�����ϳ����#Ҳx�-]�~y�c��=��� (W�\��K�\7�ȍ@g����E:o�+ǃ�t�]����~@&��g���X[]C.�C��3fd�,�;ǿJ$kRH��ߊ�M��~�`����'[g*��a�}I�$H�(5����\.�)*$�6S��{!�����յ��m�t�9sCo���7nc��bK��-��M�wHi9)�M��(m}ƐEu�ݹ֤���#�+{���$eW�(~�>�yR���1��
6�͢�j�����%������jK��^��cFiy��n��
�r K �2\�J�[�jU3��Ccl��� ���d%u�/.=������z��D�����f���޷�����늱5e�8�Jş6��u`�9k�j���.�s_M��M��a11��w��7IQ`�+�0�C����/���D�>lbH� �<Wvj�Eqq�=\������o���i��dkS ���mmJM(>䁻&X����V���!.I�]��:B�]��Sxg�P�F�{�1J�VK��r9,--!�����
�nW����֪7D�lK5��9�R	�JE�Ɋ�y��r9�n�"yV���\�ivm�J�PI�ԴG��Yg��s��C������4'6�ƥP(`{{{�������*�,�>�[�M�S��P�TP��P�בN�����j�T�A�A��]����}���͛7���
,>|�p�WYZoqI�	pu��.%�L��A�\�V�|�e]r�L�.��!��:����qD�s����9Ng��{=�"8�|��w9�=ڧ�|\ɷх��*�t�q��˷���(Y���5�.�T��#��K( �a�B�����tdQ+��v�
eƣ���T��h(�J�@�O~��"Ȑl�m�ad|ں�>�X,�Z������������2����1�տ��4�~�Y׶ ����$������8�K�Y�|���
��j544�Mu� %f����"�l�J�J+++�}�6666P,�n����[�x�ggg*(!ɂ���1�t�(���s�u�e��?�P(�Ν;���R~���KT�����9���� �7�Đ�D���j�y1g�9 7�)Di���M�i.�5ʾ���q��.|$U!pK�'���Q<��˵�[��yH�h�'U�bd�|��2>�%��t��u��2�\4�������2�����|�nA�i��DJC.�(&t,�x����o:LG����c�RQL/V��&���j��;F���<���4f0�h��'W����ຊsl��r\��+w��k��Q�
t:�+�n7�ˡV�agg�l�����zh�����h�Z888������U#�8����!��?����X__���:VVVP,���������e���8<<T����/�11�N\�۵y�N]+��e�L���o�@�J�<��$�J�ͱl6�\6�6]�N[���"YBݵ�<��n5��b*y�H���#�	 �����t����g��6q�5�>�YE��ʰ��>Mz$f�JxE���Q?�\�"6��(�oc��� ������	�2�=����r�K�1f��uu��b�b�M>l��xp��X���u�<�+��3s��&j?�(�7�d��pk�J��
9��ۣr�dj�P*�����>������ϟ?�l6�������8��h���}��7x��nݺ�4��\��������JJ���o�!Ew�uD�r�[��3>�|X8_� emƥ
׊��ЌE g�5�6P���>)l9�|�vIt}�i3�-����2hߥy�?_>�k��4�l`Uj���e�c_��%�Ct�f�$`�rC��yr���еƖV��Z��R ����y���@7H6�P7iPgZ`Q�m~�:��1��~k@5�������P���FeK!F9tL����uٱ��	���4�i��)Ɠ�� �Φ��3ݘ�����S��۴F��dJ�!��� �� ��X��}T*\\\������J�@�M��eloo�����>VVV�{) �]��w����2,�~)j�X��ױ���j�z��8����r��4�,H��i]Gρ��f3L���#���f��沘a���śBqX=[������Շ׶?��f5�-.K�"N����d\mMuB�w�s�:�y��כl0R$g��$2����n��k�R(�҄K��a\W�"�YUD-�Jz��:n�:븴+.y��B0�]>F�$.+7�y_��W �X,zWU�^�C�4\ �U�Ł��&ɔ���N��h4�Zr�u7���� �K]���&��II��Z^^ƭ[�������#Ul%A_�^����ܹ�:���iȒ�@0�x�a{vv�t��H�d��)��w��V�x��>|���-T*�k��6Ƒ�����3�.��|>�rK0�]��I��$��}�Wfͥ���ZPq}� ��zu^�i+t����J�N���&&7�Mx�`�`�8 ���o�K���DٚS$=��3�Q.^Z������.�Nԉe����m��r��t	Kj����C���;�0����7;pݓ�)���'�t�?��!�N�/��\�#���81.QR��bP�N���bbUm�(���X� ��j����ulnn��`��P�.=�;w����sJ����m�����'�x��O?��۷jNKgY�e��]&����x��1>��3lmm�T*)�"5�.������ڃ���|�0�A��$�f�sB����y�yŞ*�}�t���lŝ2����F��u�MP]ƕ�H�3���`:�Mgv(�~.J7My��Z-�0�������<i���#1�:K!�c�zH��O�X[S��Sj��7_t&�����n�N\�@!�-�/lK�]��mL�Idz�>���[%�y#w[���>x�3beL���17��$��G���D���.`�%k8��/��� Y4FZ�Z����lmmauu�f�nW��	���a���j�K�6��$� 
�E���(�Kms�n����x����    IDAT�4.d�E�Az���u|��W��˯p��=,--!�N����C����S���|>p���"���4'�O�(]���D���9
@��w�v���}�h��m�C�e]�.+�S7�����*�@e�gq�L���Y��2��b�(&kW�5�$�I�y���.�
Ѧa��X|(q_'m!�7��W�v��*�lnۛ�MZ��φfZ����&�0�>�o��i��T���C�Ť�0�_����Gb
���b%(�(w5j���nl���IwL�Ciԋ�������(�jR������J%��u��u,--)f�~w<�\.�^�cmmMY���$	1���@���u��y�E��e<�Ϟ=S���h42�����>��>
��߿�o���?��Ǐ����*⥖��7][��G��A��F�۝k�K�d�_dc^0�]1������P�����k���g��w�ٹ8�P���%��3@!D��L�խ�H��3� �E9���������ˍ�%��YQ�Wȼu��z�H�L�o�l��H6F4l��V���4=x��c��EH���|��1C����v]wt4΢�ǐE�ӽK��6]Wꔳv�|�C}�AsFlgi��2�)�N���ŕ��R�46�� ggg���@���h4B�P�J��r�����t 	B�\~�0�c���#�^�byy<P��t:���h4Z_g#M��x��1���?��G�+ MVaRWKך���zuu���#����^OI
|4ܺ�<�M��[I�"��|,)�����}6����KE������:j^��%,:��G�aj�&6�Fr��MR�8�|ry��j[s_�l�5��h��@G�ߺy��sCrPC��\�H_>�D�1ηE�!÷-]h����vd��(�[\Rh���o>��K~�������EH��L�C�R�ʁ��y���Ӑ55ЉR�c;89sO� Q�O|���T���H��j��h40{L�p8���	�����`��n�����3��˸��z�X���>Z��bd��q�nll`ii	������/���C���+fZ�KbF��,��>��ϱ�����e�G��z�U�sɍNSΥ.�=�2f9@�m�}��P0jm��S��@�ƒJ�k
���6?T���,X�yF!���}�?����\�NT��[!��lf��q�nWf��w��n�:��9�B�(�">����?h6����tQ�>2[��7�k{^!ip�M7�V��Ԍn�����`��
m�"���&���!m @j�r�+�l�J�!�������+�8�@��R	�r�B�fS7�dQ��ū���6...pzz���3�)��F��!������;ܻwO5s(���h6�s)}~���a r�������[\^^��� �ϣT*��뗗�����;w��޽{�}�6��*&�	����C�z��yL�S\^^boo/^��/��2�=��ĵ12�"&�� &N�#5�:Pe+>��M��F�uG�}_�sǖ���@�����{�Oџ�~y��*V�9�]�x��u�� �k��D�7�|L��(	;���[�8D�d�*&I�耮���큻��Lz���u��|��\��s��*|�hM����0TۭKݸһ&�H�5���|�y�+�����3[��c����)J��3fK�W4���Fi��|�٬����h�& ���U��� �f����������\���h�����C4ܾ}{�� =ɤ���\ayy���C�����r���1H ����
VWWq��-UPF�ϛ^�|"����t�vx��vwwq||��l�R�t̄�K�'�{���@�"����]Bt2��:C��I1d.�����do�A�u^�W*Y׌�x�� ��1Q@s��Z\|`���,B�J�\��|t9>H�ꋜ�+e���w��[�br1k.P�Ƶ��Hη:0��mK��62�r�>ZӸ�����=7�@�蹢~�-��� �L&�T:�Rs �@*O�c*MEa&`¼�����#�yI�zy�0�L�<8���vqvv�ׯ_�ŋx��z��\�'�2e2�z=���boo�o�F�V�l6C�RQ��t���8P��T*�z��r����5�z=�z=��!ï?�ɠ^��Z��T*���v�s����[��l6���[���Ox��9NOO1��.׶G� \�o-��f�N��@yS�\�C?����bK�&If$qn�
X]�-�)��.Mg��ö��|�;���F,�C9*>0Y6��&<�#�t�-���R���e-���>g�Î�w곈\v���4��ˌ��.��-!^�I>�}�ϔbJ��Õ�I��#�'0@�^ �Τ��O&�kzD2$c����!�;�C-t?�I��̋����-@:%��0�+z����s|���x��)NNN�>�.b��)��&^�x���x<�'�|�r��ޣ+��d�r����� �:j��bQ��g��� �Z-��ӧx��	^�z������]Ť��ʘYy:h9��.>*_C~ߗ��_{�O���D�6~��	&��;��&�����Nd>�y�BV[�ɐ}���}���<�uq-<������� �5>RB"�{L��~e�z(Q@���8j�8]���P1�M�I��t��}7m٘x��OA��Ƿ�9q_�]6͵�;�Ԁ�
����0��J��D	BR��LN��@�CEZ�>JG��D�r4���/^���������x���ݮ
6d�L�����_�F��A:�F�VC�^W�ޝL����,�;u@��Gϛϳ|>��Ho2����/_�ē'O���S�}�VuB�f�J�`�>+u��g�/S�5�I�nT�e�}�u�`,���G��['��e�|2K���S�����x:
�c��]�.�����g�5A�]�2��#wr���[O|��]�_��²�p�Q$��S�e��z��·�K}'��>b�RI�P�/�)���R��
�ec���ݶ	���M��*��ߦ���-OWtf����Æ˃����@"�S�:�r�U]�R�+��B�(���5wD��uU��Ipu1���WWW���D��R���r� �G�����<{����_���ﰷ�����}�=��$Ă>y�D1���[[[s�	�<(���@��wt?�`r	g�9�õ����k��x��-~��g<}����J&Cn|.�Һ���kkա��w	���ԘD�C�`��Ѵ��du���E��+5n�G�9��g�M0y>�E_	0M��6V��d�����LA���|>?��b�9�u���Bcړ�3'}�sm��m��C�e}'�-�������I�msQ��L�RI�* ��t0U�O,EB�����u�����]:��~�R1�[�e�O|��kn�D�Ѿρ%�b�'.�'v�:�QŻ���x���8+@s7j�a����y���Z�����8==E��R�`ܕ��Q	h $أ�#<�������S���5Sa�b�n?���j<��׿��k��0��`O�w�r�$�&��f�Ϡߡ��v�h�Z����w�}�'�~�ׯ_+]�,�2�Pu���I�����-�� �I#�I_^��DǠh��4.ݑL���ڍG�U�]o{=Ӿo"�L~��=Ԕҗ ��o���u^Giծ#T\�5��׹��}����&D6�N��Xm��� �]n�A� ����`p���C)x6a�^X�y�U�Bvf�.�[���褊�L��xj�j�J�Ҝ6��l�@��"��G�=�i�ښK�0�鯐g��º���a��V�6�$�����l�o�s�keө�6Z�ZZ[q��,r?\S�0�F�������<�^�7�q�X,*�C�%�kB&��p8���1�>}����}�^�~��8T*��z�g�Y
���O?�����ϱ���
���`3���Ϟмx�_W��W�y�J�����������������H1���9����/���n��V��-�}*���(�,8g�}S�&��v7�~�Զ���&ϧ;��l���#ory�&����2L�������s�Q��\�+q���N��'�.�S=R��d)�s�>�v�XCِ���$���τ�9�dtI�~>�W)Cz`�������R��ᾍ� �N&�ߜM2�(�ä/ӥ�M����5��o�<�"��A�R��Y�)q]�nS$�0�8���V|'�D�V��1O� �[0��6����v�n������\�_��R	�lWWW8==ſ��o���ǋ/���kt�]�j5#�5ɗ��4
���):�޾}���+ ?~��?��Z�\��@�h��O�w$����`x托�J���l�F��/^���g��������t�i���4���lj.pQs�"�_{�ŕ��vкk�V	�C�CQ�>2	�.u�&pU3���=�|�.#� 34/)� ��tZfh4)��M��6ϊP����A�df�v�.]��
p��x>�>����ڢ�D��t����:0�\Y���Φ�Od�X9�"D�u��_�X�Q�c \�%�l3��[/rEq�H�e���i�l��}9:�)�澡�=-�c�p���s�����RPr���6��o�A	�|)Sjn:����+pKk�P((֖��b��b���`���#<y����?�����h�����T*�<�M�C{
��%P�VH��h�Z�L&���H���������4:M�n�ϕ�S���F���������'^�|�~��J�2'�ХYmsWī�7�b������8�{Lk���O[iY�'א�æ{�d��~n�db���n�L{\�rÏl9i%3�>͖������Y1H|��\��ݜ���/��m�Ƞ��i���|a8�V߼����´����8i�2� ��.�ڥ�E@�6)����O�nO��u;�'/�����h��5��:��� \�嶨_J$nz���\��-��)\�O2`�N�\J����i��-f��整�ůܺt⺂�ж׶��|	�v;�u��T�=�Og��U��/��/^����'���[�P(�\.�X,"��i�1�9B�I�A��=lww�� �R	�z�\���(�JJ2E�M,���-�ե8ep���qyy�_~�?��#~|�#^�|�V��e�^e*����3�2�Fb�p�0]Ai��6�'>�}�V��;΢� �d8}ص��Q����Q�w���ǲ�J�����-�$��T��.���r��5���x1�$.8�=c���9�#��7��h4B>��p8T�2ab�U��5}�K2Ř��]�{��R��A�À���2�S���:���3icq�l�����ë����(ū��d6�w��)n��g��m_�d\�B���MB�?�֗��>���Nf��\�][������d2�d<�����U�cr��	VC��;܎O����;�J%�C��9��`0@�����	^�|���?�����զOR&[�'���QW��b����}�������F������uՂ�Tu���w�!�?͙n����S�{��^���������99��2H�� �$������]�t2����H��K��L���Ҵ|�J��Z����k�윏�ϼ�ҙ��9����|��Wc��>L{T"�ߋ��׵������R'������$ڃ�'�����|~rْ�w�9�����,��ct2J]a�C�O��.>�

|��ЙR��R@��h��~�X,*H�z�^� ���u��d�,t:����v��+׊��봔�	�|M"�Mj��x\R����B#D�y����z��6v��Z��L���xn^�FH�@n&4�i,��������\�ui�_�r��p8������P�T�������z�>���vq||���]�|�o޼Q�hi,uA�+X�.R&U��������[%����q��T*���ayy�{��� }`yU�p0�h��Jmoo�^����޾}�N��
oi���L�N���3��M?d(Ȑ���懷m���$���{N����w<+���h�z�{I\ɟ����8�8�l�u�<+ľ-�	'����63�FuA��d�I$����ͤqM�ӨT*�T*XYYQ�r��`�a&_mZ�E��	�~��^�?�h;#�gͳҼH�kre�C]�R���|}�N6���ggg��x<��Ր�`�5�B#9��z�&�hzN��"��̥h�䀖ؔR��6,��Q{K	�i�e/;���j�Z���|?q~-h4ʺ���(�sig�u���اyA�ѿ�q9��(�tZ7�rZ�����ӽ�/n�y��#��$a6��ѡK��6��Y.���h��B�\����h�=��&9L�e+��iy�����8::­[�����J�2�==88���quu�^��B��Z��ݦ�+��e�Y�J%t:b8�������V��������5M��&H���>���5[�^��g��z㸲����S�<O�(ɳ�<vW�D6T��J�^@~l��?���R���6��.�ڲU�5�c2�9ϙ�!��v���$顪�%�LfF����k��V���}j�Z���OO�>�Z�Ɵ�QJ�-K
�u~�{
I�բ^�gs�����s���x����hT��$��$e%guZ{�?
Q<�p8̴��x�g>�d2Yp�C�G6�~N�%�Q��Z��R��u�?=h�:��3�ǰ��@�iϪ	��~9!�rK���`0�4(��@�)��eY<��C�Z�z�b��ˁ���s���GR���ˎ8���j����N�e��/Mp����?��?o!��,�2��y�Bnmp'����	�tFY���DC��Z�E�eQ,�
	���(�Q8���Hn���}���C�H�\�ۥt:�h�Mg̿k4�j���䄅�QQ!ApEŇE&tu�[�ܞ]ur�Y�V�b���H��*J��#�T�"�2)�mT9���.3�@P���k[�$�
��(
�OL��A�J1�B!�Jj�|>�\啝�Ox���Q[g�ٌj���u��Ȳ,����'�	�j5��j�j��C&%�tɽ��[��D��Z�ݻw�?~L�e�?�@�T�c��v�𱪀Z�4F�5ĩ~��_����f�D�2	1/�n��%ޯD�����u�t:g���\�/�a���ړ�A=�� �@��{<�t:��^�G�^Ϧ/���)q#�6��t�鄓��h�]>  :j��j[vWt��,��ppɃSGѫ��e[�_Fr�+��S��W�	�����@R�P�2���i.�-ˢD"�ؓ��|����T0��tJ�~ߖ8YT��$u0P"��*4X���l�D	,�Q�$/�	����S�q�j)+QL,���J�Y���B�1
Q$a�A2��!
,|=�sb�KeKP�`0���<E����";-������1�Z-j���n�mhH~dkwJ�ܒ��.�U�\nɧ�Bw�(,�A�ҾRy��}V]�ˆ>dU/�@�P�!9��^:����N�4�/�P(�m�J� \�2q� ���W�~W����e��)��}����"���(8�������ԭQY�������lR�^�Z���:,fK�Oe����@�0��%mȷD�/�pJ8u��{'�e�'QXy/��2&��2I@r�/�L2b��CQ�$�E�<�^ʁby8Qh��0E�Q��z=
&�0�{ &ՍJǁ\<��-�S���v��րS�Xf䰪6���I�][p
�Mg� �|�0�M�R���(�JQ2���;u Mv�U��m�K�M����������s1��v���p�ND��V;%@��Y�����kl2ݐ���V�M�]"O���ȿ�M�/$�$�W�H�L�ev��3��8�b���������l�H�CA�RX�E�iR�X�R�D�z����������������&M�FU�HK3
ɯS� �8K�<��k���*��2!v]{d���eo�px��*���hf2�� ��-ˊA��.�֍N���G0�E5�o$H�����z�ڍ˒%���BTU+��_}�Hml/��y��Il���H��-7N�U.I�D�%�/�rQ��i�z�*v*�������D�����j[G�    IDAT�y���q.X�E�L�R�E�Q���[(�3��:����-��R����b1J�ӌ����P�ղ�a��p8�='5��srXt����$׍;}Y1S�?V�#vKVW�۫�Sj�H���t �e˲(�NS.�c�=x��Т��7�g���B|S��Hn%��S匇\� �b1� �m�Z���t:��t8�� w�C�K"�C�n�֪ �J	�W�n�������Ps�)D� �m#���k�ߧ�pa���Xz�J�l� ԩb<�V�Ś��V�N.�/��x9< .�+y�"�b��Z�R�^�����ݥ�O�R���d��h9-/�w��V��\��e��k��kr
�Nd���e�t߃@�(��P0D�P�F9A��$�UN���#�g����q��g/�i%�����hD�N�"���4.XR�Y&jn��n�F�P ���k�3��-��q[k�b�D�����wf�����=H�����W�7�UZ ��u�s�3��Lr�ݳ�뉄-`�	p��|_P�T��q��|E��~�ϝH�0(��{\��cz�p8�u����������99:�2�%iSMc܆{W�yIZ���E(��/T<7�0H3�.��G�X�2���y�T*��d��͔72�Г�mo@�[�S��;ٍQD��J��"Q�o�ؗ�i�7x�#����yne�n�m{�I������	�E2d�6�E��B���Kq@�H���0o6��X,�T�` Hf�dB6xgH.P�Z-FRTn����F�t�����Z�%�4)�NS2��\.G�R���*=~���<y�|]p^$�\ '}�_�]�ĝ��qY�����:{LHE��.q��}$�@hKJ�|fw��IK����S�G$���t�^�pT�r�Fת\�v�4xfq+tt�G��+�>W�~��T�P0�@��@��F��m� [:p'���EZ�IqB�$He���S]��9!!E�B+���|N�h���$�Z`���^R�Xw��d	���L�iCa�=G��s'�Hp����̆a0~�:쨮�e(��$�I�@��_%�p3�q�~�ΣZ4��{u����=Xףшci,�ĶR�P�P`><kH���� I+rJU�l�6�Ϩ ��o��e�X���F����z����J�\,�J�� q���=����7� �c�7��"��ݨ����֢4'
������
hm("��w����DXL*�/����|>?3�����ق)`}pq��8
�f���fi��<y�� ��Nh��"ߗYE�% rmx���LZ�[�Ἧ'��;��H$B�`��0���	M��gZ㒳%[�Ʉ�#����kRNL���V�(���	"P*$$X@�6�W�h��pS��b<�����Wv�K<��H�|]�>��[u�W�%���ċ5�N6mY��A9I ����R<i$�ɄF��qc�5"�Ņn�2�k����p��Z��M�����	��� �b0�eY�n�����x<f*]2�d*[��<#%�Tdxy����+���2^����υX(U t� ����H�;���tzq��T.�)��r,E�T��`0`
 �H�C��K)�~T�Q�~e���R؛(�&}>e�Yη������Ė?J&�d�&��d�oYG�2h��e%6�}pj����X,F�T��}�w���3C#�D�ʕ2��H�=$�����Z���cj���P%�Zj�����;x�Xo����eY���)��P"��D"A�l�����������ﾣF��2 hq�~Ὢ�ë��~����e��{��9���*:�ջDb��h4J�T���dB��sN��l6�v�m㝣�5�5�rq���m\�؟�p ���Or����I�D�I��Zq[��e�<�k�-0;���R�C��,{�n2���6�*u�<{�뀡\�:
�,��d�U�����1��3�� I��8�b%J+-F%�!9�~�5uO�A
�VJ��4�i:[�t��#iA�gx�-����^�S$��lf�U�Jyߝ��Uy�a/��=��[V�y�aV?�d�"G�̜���6��3`%�;�#���%X�5�3_�ˢX�]J

!ۥn�<l�������\ǘoB�+�qvd���j����ؤ���	[%PzIlW�d�Zn�Na�0��F'ڢ��I��t�2�e�Y��^"1/
AM&�%����d���gY��Ln}>ќ��	���V���!��.O�Cu�d2��e2��>{��:��m�����8��P�#VI�W{v��_%�L¬	Ƀ��h4�-Ri�,+i��� $��^��Z8p��S+c�n�a$�*���/��A�="�SdpU�*,ˢ~��:�l:*�n����ƫ���X�sn�FnZ�n4�`�S�G�-���P�ڽ:dJ��^���'7kW�C�RJO7�.yߒ�JD�� ..���)/q�%5m0���Ȯ�l6��o�E�T��A�� ���|LU����Ϩ���^�T�ux�zMp��ewx�֖��ʋ��S��F��U� 2I3��G�d��]�F�N�mT�n��I���"���I�X�� ���%ו���&�񘇆��$"�v�����ဈ�%	�ۀ
���>����z0�t:M�D��3��-]�T�'���_��-�] `���'�	'�P0��ؠJ������n�����GU,]�p�ȃ������n�4�a���r�BC �I��̕���f���.5^,�h�*���K��~P��eQh$*�P��q�*��a����;����r�5sC��p����-~)��{ 8У��	$H5��%H�Q�I),h����� mJ���u�`.���m��!����R�̹q���C� ��3�n��VzT�v��v�=��oT]���g��kms�tH��9���5�ju*۪���`i�U�awR-`��P �#2�U[����ߥ��t��G�F|���q��t||L�����v��jq2�F�T*-Άh�����l� ����V�y=��4�/��p�����R@��y~A�<�mP�:�1� ]�z��]�F�R�U�����YX�� R� �t�X,�C_R�� �r��v�}��&�'��o-��{$�7���2�@4�O0�z���4~՜	�l���e�lL5�,w�a�	k����,�D�LӤB�@�\��\�B�R������a�A7Z���dK(�\.G~�����Ʉ��$��=���jNJ���-��X�:�r����!L(��'"nw��~�$�������S�#>�D��-�_M�2��UW�����rk�Dq��xBr+��P� �����|�1@��-j�Hm{�nA(�����"x�n�_-6� $x�8N�^���V�ףV�E�z}�	��!�uM��зJԉF�~�����U�ʲ�:%;����Lt���t�g�C�'����[(���:ȟ�:��0 gRzO}��_؟R�s�(� �k�f3"���Ș�I�|���������)������'O���*Pky6-��*��cˆ���.J�S,������3�/0l(��ǹ�v����؏5 *&bw0�h,�sF�����.�n��Ͻ�=:88�i�#�W�� e>:���h�4��D"�]�H$¼��N��g��j��-+�ϻ�̋��^��� �_�-x(��D"T,�R�P6��MND�n���j1�ӧһU	�Z�F �t#�q�g���B5��
uK1pi���L��B;��X�h.&���JZ�z�ग�JRz�A�ˢ<��@{�(v�luZ�*�ɭ|>j+NF�P�ʃR��^.+�^�t"���ˊ��+9�*��E���z=��y�lww�Z��#����`���T�쑋$����t7V�T��/*�
���g������1�N�o��z��������i�>�d�ɠ�a�]��2����:�*'��Wɉ���c$��X���*��s:::�z�N�v�|>�R)J�R��!������sϭ��渨�P�	��eJ<^^C��2f]�	*�P����f�K���mr�6ѱ�z�x��hY��)Jg�
�����i�>��	�:�(�g�D�f0�D�,A:	���1I.�8�á�{��� ȳ�B!^�����w4��q�Yx��m�Ln�[ݠ��)�d2I�J���*��y
G�l)<m	.�6�0`� i#<L8���	��	�:�2 %�/�\�1$��T:��6�8��_$�l��eY��F��rն�*�~��2����X?.k����ŕ	��� Z	Z7����P�]Q���Dle�I&��i���p��2���k�rJ:�� p��� ��e,[[���V�P��)t��P�eJN{�+��<���&��"ͫ�|�ࡤ��T��|f�U5F�y��c��l�2�0�iu��b��xViH@ڜ�	U�a�н?�#�R.��^��� ?'�	e2�,���2�f>~����A�SѸe(�zN_�^��}.x��s[����ſT����P&1/���S�6.$P���L�i&��\.�Bf���oe��@(ںv���E�����g�aܜN��X,v�4��~��Hk��g���t��xL�V��t-���T΀~��j��G�P���$M�S��V=���K��2���hA��,x�����"�Si
G����G�	��`�B$	<�1��^I���b��ʅ(V��U$Z&3�� =�4)�Jq����.����BA�ỵ�5��8ʲm�@�?�%\^�bN(�@���^��.�Է�E�r(AjjJ.�Ӂ�j �&0�>o�J�W��%Z��J.8�Wjr���B<�.-H��,��U=�p�wT�k�u
k��U�.:�+�ܔ!�Rl�I�yEt�4&�x�^�חY+{�X��\DD6�v����r�`͢ �
�"�:d:~��"�Q�BT�[�\�',��T�0�ge��g��\�Z��K�L�2���=zD�v��Ȓ�K�$���sAG��C�,wu�8���c`:��B�@�J�R��͠	�֦�H�5�M bz��n�R��X,�F�[/����e��R��MD�DD�Z��x|���C���d2��B
�X��p�?�vr��Á����(���d��̹.K��\�_u�8-:<\���*�0*����A�j����6C��BL���-�pS�;�A�Kj�ʊY��T�LP������RGW*>�H¤��:�7i<�P��Ɠ�%X$�C=����<<<�V ui=,՗�/]�>��Z�N�����y*Dr�X��Jz�D����n�F&��L9}~P$����P%"��:�I�<(�`��6�3?���K��H�Sw�.�Ӽ��	�S������i�z�Z��Š��
y��U�
nC�j"aK��Qʵ$U$}@x��5�=��T����l>�Q��>��Q�Qd2-��*����Y����hyK�R*��D��n��/x��R���4w?��9=x��&���C*ϓ���z�n��Nno���>T�5㌇n}*��B�@�B���$E�Q�>��wX��H&�L�6!u�L&i>�o�F���p�λﾻ�c���\��݇~6�Ln���|>�97ahm��J�P5�q�+�J4������/� P�u:�v��hzϻ8.���B!�҂�!��r�mllЕ+W(�ɰ�X�������������T�׹��v/l����LD���t+��dKX
j�;�f�P�a�X����Ф���|>O��B5b0P����k��4xc�:2��J��	���$J��]�)�	s/���(��P\/��W�t]��嵑�B�ɭD��A+ב�$D��s;T0�"\Pԁ0MrR7��[�ی@�;��`R����ؒ�U;��-'��7�L�{�_e�SM�ϓ0�PY��X7,���wz�n��3G�ڒ3�g*w6��t6���Ngl���``�lh�:��Z˂L'�%$9�%�|2ٜL'�����0�P����trrB�P�à��?b���q����mz������E��tJ^�S/_[���|^\������"��S�r��^�J�d�:���x�N5L0�:�)8��L&o[�u�a�ɯ�W�r����������`0x@�p8di:�(�n��7�{H�ΏF#:C��}�����YP0u�*��2\,T�h��r9*
��B-!P�T�k׮Q�Z�t:M�aP��cuٲJ$���NW�\�|>O�t���8�ݦZ�F�f�ۨ�\�B��6m��atC-��������s-����������p8=�%������t��h4��h���	ˁaڿ�b�r�u::<<���]֌����c�@����S�ۥ��}�U�
�-�e-�eډN�m|� t�v����N_ӽ7T�Hn��(O�JQx�o:QTz~Ed�P���"��H@��'��U���RuC&�h�IMF�B�yj�/*xt@��$t-P��N�^�47�;����y^E/�*ɰۡ�L��k2�K�$�U�P���`�<�pK!�%i`,o7��9�0�g�hn�)`��nV2��]�.��Tr�%=IRؐ�J�����.���ɽ(�m����l|�N��C>�T���2M�S:99�}?�i���t�D��r�fܐ8��n�ǋ��*�)%�Խ��#�NS�\�+W�P�P`Z���u��n�&�J%��v�]:::�P(D�r����v0�����\�~�gIluו+Wv���>6��d2������pڃy	
(�j���Il4�\6ǔ��b�G��3Θ�c�c�J��t���U����<��(S&��|>O�x�&�����P.��:�v�trr�~� h�A�d2��H���>��u2���2e2*�J��v����7�ܹ�E������ٳ�z�އ�X�l6�Y�����vww�^���Ǐ����oR�P��;����/�吐���b\,��u�t:ttt��K��ǈ�<�V���8�$]E�W�^��kp�� �X�0
�q�U
��w�K��Db �
ѝ �  �<�����B'�Qr��MU�6��A	3�3���e�L&l=*e���ܒB��"�4�k����'���ҧK�T�*�@���M������&*npX�*b�����S$�T��S"�)M�$��G�o�6���l�tX�
^v#P�ʢT�H!�<ɽ�bo>����eY���a�>�N��P�*!qB��.�,l1����R�����)R\ƹ���]En�%�5�ŨP(���:��yFc��:� ����"�&(x
���e���;�P���_�R�˺��2�3�=�u:�:������Y�a��.{$a�-	S.�#�0���Ȇ�b1~H���^Ur�5�<<�U����c�e�Yvꂋ�b��4U�U��r�Ռa0|`> Z�x���j�����^{�5�F��>�o+��,��*�J?ɢ�V��D����{g0��B�j�z�ڵk�����ӧt��}���T.�)��Q�P"��H$B���g���:���q��UF��t��MUE]��"�N?��2'�u(�[2$����$9�@B��!��$�Z?"y��2a}9��Cܫp�D�U�X�-@�!"��%�J";�`���$��eX���H����t(�>dr{�eCS�M��7����ڔ�U��J]� ���R{t��m`s������f�c��HHI0�G&��u�SPp��D|Yg[���=��:U��!���=���q<>>f�&�G ( ���x�g���v��:xO^h_^���(��@��tڔɭ�� ���c�F�T.��T*���`0�N�CD�y��-��d8���L<�r����fo'�;�j��ܪ�eY�#�)�J%��M��I�{T�K�iIq��3fI� '	�ġHĺu*��b��Ԋ��&�@� ��b���l��DȊ,y��)���S���v�|>�b�H�jr'�||�ʕ�m1U*�����ч~���J����w����>ݽ{���t:M�X�̀���V����HrG�'"�R�e���:/>�*$wU����E�H��f�D�
5$}�D+C ;��uAHB��h�j��R�C��?/�T�[�"�Uc
�D�.����~!�E[��nۼ�%b#Ql/Z��R��<��^ѝ�$�?%�+��*�B�����<f%ӯQ    IDATb����U��Hr�!�Z�C9��&�j��j�)M�χ糅��>T��:)�mu��r�T�b��~�����?/@�tI�*t�d�+ݪ����1�v/���Z-�N�< +��.�:i�J��W���cU�w'��e%ɛ��I��EZ__�b�H�h�F�5�M��\�� 1���0��(��R<߉D"�X�֥;�}����;�X�C"����m�j5�U<��R��"��P��4)bE(���P���טi^4(;UV*	���d�b��.��)��a�ڈ�b�ܢz��z4�ϹMK��`H�^���'�	
z��W)��o�b��|>H&�[�|���0�x���;�V��`0�Q�P���ۣ�w�R�^g�E2��1�N���S/z�;h��A�x����i:�ғ'Ohoo��YRJuW�J?��܋�h˸��-y��P��8��#�C�FmwI�8���:ɃU/^C�W�v x}v�wKp�>T�*a��m��s����{����3~��b�:�M�S��	=��ƪ��xx-~.���)֬��K�IM6�	�%!�����K�%�_9Hƿ�8�@˂((?j�*8)-��i�E�Ni�z����mT�3J���j�w�$BH�$MG���|l�D���N9�H���$+(Rc�*6�nH�*˗�O�8�N�Uv�t�CP�l�666h}}��b��Z��\�@`�q��T�B�m�P�����_Tr+�+W�l��_|����>���7h�(Je���Ui�$���ƣ1Վ�כJ��,j�Z܅V����6��,dME��� ����Q�ۥh4��-8�8`����-���V�j�>���	Y�Eׯ_�W_}�J��N,���W_�E/�SR���_~���f?�f�7<x@�~�-=x��666�7ޠjuap��Z����$�|��=zD�fӆ!pJ*~L��:YP%~t]�g��*�S�J%SdL[2�E�	�����x�P��s�mEu�L��(5������Iu�<1܆A��ph*��E*��lF3��p\�Z��h.ڣ���ӡ�Ja����l^��:�������Wu���/�N�p����M�fi�ٓ���LBU�Eg򠢷��ɨ����'y�*oX�<����ɰ��phQJ}Q����)�TH����N��l6ٴh0(k �����\]&�T ��LEr���.#�u���bϮ+n$  �hmm�*�
%	6_'W)P� er4Q2�$˲�����D"q秢F���{ｷs���[�H��D"q�O'''�D����T7(Ba���**P�T*�|p�u�uk�\� ���jCB�J3�ɰ�T� ��yZ__�l6ksʐ�5�ա�����z����\n�R���d2w����b�;Ｓ���Ï}>߇����X,����cz��1�6��*�R)�` ��f��,P���l��Hޭj=�z�s��.;�un<�mG�����d�J��J%�D"6�ԉ+������N�$���cQ&�yUZ�u� �(��� �p���6%�%�C|��d��	* "z���]��G�C*���T�y�=���&�^���)y�Nj8n.l�|^��n��~���5_Ng�����Tt�
/���<԰%���tJ$���3��򞙦I�#ج���S�������L'���ާ�f���zJ}�R�dӵF[]5�qKp���^$"�욝�U�U[��k���HnK����S:��X��P�f��WB����Q4�d2��N�?~뭷�*[y���;����B����G�^o��ӧ�/0�����1ǿe�Y���C��i��w�Au���|�HpW�@v
~�#Z��d�y�؄�ш��J%*��<P �2Z*h��EJ�R4������<yB�v�*�
����ھ����	t���V�\�4�N���o����uX*��X�B0M���&�bhm�%":99azC��bʈ�ɡ���Q/��-�׵�TN��p���sJ�C�%�	���<d�B���E�'y��;�&�þS�����FR#T&���z�t��L�%���� �%಄��\��`Ҷ��A��P?].'���e�E�m�#�1^�ܫ�[�A��z�}��-������s��t{W^6兹�E�Q7t���)�� ��'�0��i��j:�/~n�S1|>���ݪ蠤%�#6��[r��@8�d2ɪHn�����tC�q�&�}t�e:~��y7��-v��Kj�jT0�L(�Q�Z��W��\L�dA��-�X@n4�R)��ؠd2y���^��Knqa�h�^��N�ot�]�У#�3*(���H$���z���P��>�Nnɜ��Z^.����(�JQ>�g�B8uY�E�R���*%�I[*��B���*U*""z��=~���U�Uz���R���[�-��s\������������Z��O�n��'O�P<'�0Ŏ�����5$VR�&����~�$����
�䥭�j�j5�k�9X]�,�x�*�
�sy��F%@N0���Db%mA*-�j��b��ФJC�3���(�d2�R$}�Fjbx����H	"bZ�y9E>��Y�Yz�}�XGWpJJ��U:�P�W�����Z���]Pw�ִS�vDz�'_G�9U<_j��])τ�i����M�N����3�N��erc}9��H�\��g��gd�O�H0`OR�B�I=T�iP^��}�a�q8�{֙�H^0�t:�<w�B��b1*���l6i:�����o��Du�gPiON�mY�v�cs*<�Sn��)1�����<E�X��_~���*K|��I{�H$�Z�N���B����fo�b�����U*�v�޽{+
}bY��x<f�Z��`��@� ��f����v9& ρL�Z���K�0uU���U�.�JB?.ذ�E�HsZpO�� ���tl�6>x.��@ @�z���Xa��7������T*u�P(��TI�lv������������o��������!���+lE,�)x��1�6��(`�X��jQ�ٴ%8���Z˞ׯ�2%��daܒ74ω���؁@&�0J�DV��#q��"�p�u����,�����Oǳ�S�H�{��n��ꁂ��A�/HO�n�u����??�g���B�*�=�n�X,F�|�Q����5�e�u��:��2�rU����{E���n:��ڰ����C������'�uDԤZ�j�=;5���5�W���u��j��ji�3J�w�~��'��|O�v?c�1��u�K]���2�#Ԇ�U�S=�ɶ�`c�K�����u7��	Myt����
計�"ԍӫ[���*�K`,�3��:fV�ߩ��B�?���lj�����0��z�d2��dvR���/���_-r�DY�ӟ�t{:�n"�C������nRFl2���f��⢸�ك� �[~b�s���@��Y�MiYO�[u��h,�RB�V������y6����=|���T*��o�M;�d�*��W>��m��M"����ҽ{�h2��;�C�t��l.���&u:��^p,Jy�S���Dȳ��m\�^�j���@�1.�������N�'e�xxj:#��q�a��,�d@-$�{z��Ȳ,����~�T�nB�?����A�C�C�����h2&����z��b0Itչt��T�Ȗ��A�Cs��e���֦R���6 ��8g��.�%��:�G�ϭ@]�9�Z���T4�?�8HSb�Ū��RZ�:r?J>�D���]K�d&��J����-���u6�8�Q3��G��־DD�V�:Q8��q���S��W��e�nox�8b畝s�R�W��,���"�ѝ8'��Yh��f3�t:�G��B���;S�-�x<~g6��v6��@��H$(�УǏl ���Ca*���C�R���K;�Sp�K罜N���,�eQ.��L&cs[j6��j�h0���H$­ړ���ݥ�O�R"���6��*���\.o����"�O���������O�R�\懎�Di͊?�eq�^����A���~^ܐ��q/#��!T^��ː_�7���4�,
��"��m=��!�x<��D:�I�#�B'Y�o�).A�A���6�S6�eQn���~�������p�	D	<���6ί�_�rHx�d��N~�	��@8����25�qZ3?�`�.y�I�etF��'/	�2��U�6$�,�-A����D�P������.9p$	e[1 �!��n�p8��#2F��k�$�	�w�d�Ր���|�$�I��rtrrB�N�M
t�RR���ۙ��s�K.��zN�IJQ*����5*
�Dx�V�����,�|�ªw6�a>�����7��-f����?������)��I��|%g���N�y"ǁz��j�x�K��"�I�Hp�u~�x<�d2I�|��CؐC� �b$��hD�Z��={F�p�~��_����N&����f��R�\�y��魵��O���gϞ�w�}G�ٌeՐ���=�f��~�,���(����,�J%:::�v���>TP�Z���y��ԭ�_��N��G<�9� ���H��
����}���ΦTJ��_��Ɯ�(�v���!NF�6����j&�!��G��v���6�>�Si?(�HR0d�r�?D�~�}���l6��ns"�jR��y�k��{~l[��Z�^$¼R�Y�`�ۙ�&A�k]K�.i�=��Ǚ7�����`0�%����3�&ޒ��11� �\2	���5�ј��E�}vp�q����,��A�Q�����0� ߂"$���@�c>����b8f}j��<I�WtuY��D7�?ܤ��Bߋ���&	>�� �:�,�� :��a���F�Tj'�Hܡ����W_����oow��MH��|>�d2L��C����:��b,w0	G��ۺԞ@*��/���c��b1F1I2|>���LNu���/�R�٤��]�L&��_��*��N"���Hnq�����������>�N�7�>}J�a���#�hO�v�;,��)�A�ek��L�f�v!�$��ژ���_������څ /HZ�BU �� ��CД����n9HLqx�C_����~�ɲ�����R���l6y
{4�JG6�]8�̟�����>��>��1�X�.P��l��.H 0���D"A�zݖp�H�&:��"�?%��t��:q'�#�����*�0:�5��|[��P(D�H����k`�4u�͋�����0:99���#F���@��ݳH$b����.�:Pf��F�3J(vSM�lh��9�^�	�s��dx^ �{�{���$["�n��Ub�����尯��]�âV�� z��t:͝ctBF�ߋ���jQ�X$˲�c���ׯ_��Eo�J���������f��gm[��G{{{�l6��B�Cǖe�'"�-ht�WY���sB6�d`8�ne�j��r
�ʲ,�����y`%����J��`0�WMKp�^z饝?�񏷲��'�nw�	Y9�AD��D ųI��t��j��T�ը�n�td�vT�"t�emO'�07�����J�x@2��l3�N��Z�(Hn,ֶ�	m�����֣�*	>|>ͦ3������b�WE�p�J�	n�V��xlK�{��E��rT,����6 �_R2B����~�Fm@�!�!�4����uV��mb�`yi��)�����ܐI�!�e���5�]��H~�a�U�O&��n=�H��Z���t��Z�ITv8�d���&��u���Ϡ�!HY��&�4�d�eP�'?'[��0���e��*MJ�k"�F�A�������l6K�N�VX�`����[W��prJx�����e����g��u2��2`$5��ځ8�j����eYT*�(����K��W�T�����o����ǏS���n(���J�eq�VtF�o+!��*q'�;��G�����<�!�dVN�J�|4�|~!��h4h<S�P�B���Fo�5k�-��}�ݝ�w����>�v�M�\�v?A=�:��hM!qI����t���ےZ9����WMp���]��^5���dT�Dχ��ý�RD�2�|;�_p��c���y�ݦ��c�����4�NXJEN����,9� �K�l6�1���<@u�~?�cq桁���-�0���F���������(�N���8��1�Ny=M[5�s�xIr�$o^$���"�}�2$W�YT��e�����%�n*�$�T�49I-R���\P%פJ����u(�.u��= Yda�j�l{�+@������nN��D"lRT((��s<AA��=Oh<y^4Jί���7�J�4��Ǧ�:l�J�(��P�ףgϞ�Q�Wz���F/�Q�5Վ�2Y�3K��l��x&��p8�E�+b@��Z���d�o���^�d��t:�m:��q||L��������\�za�� K^�3��%�f�;�";�|>oCu�q4���S�ݦF��v�v ��������������������~���>��jl�� �P���C�	Z����tpp@�v�����w[��{]6��*��<��-�l6K�D�6�-�\aRۯ*⤢��왦I��Bk��n���R��a)�t:�()
G�H��2���Ku�H�x���#�X,Ƈ�eY4��';҂� � �Gc�/v�`(F�߇D"�ɼ�Y�0�I�x��Z6��jWbY����	�NV�[��%ʾl�8�=�!w�"�^CUM[YJ�丫�����#)���%���\.3ET	�R��&P]8X�z=j4T�ո�h4X��=�Ni2�Pp���:Z�.y�X��J.>��ă��U Њ�d2p�n�h5���TN��������4��MR^����3u2�r���D�C�'��|�666(���~�׶_���+��o߿�V2��d6�m�9�:P����=�\	��,Kr�	����$���Ŋ��T,�\.S8f�|H�]�DXw0еkר\.o����/�"*�˟�g��o�6#����X�|�@0��&� Y� Ξ>}J�F��+�ܐ���?/��ݒ�U�?iш�m<���	�1����S�r�Z�!$�vX�ߧ��#:<<d��E�R)
�E�	dy4�� PU$�*R%#Xh#_�~���(�j5��ߧN�C�|����Q>�gS��������C\5)��� ID$ad-Z8���q��z䰙�"J')������uJ
�;'A{/�ߩ��V�J=g���ZGܖË:3	]r|^��b!��T�U�v�jA;!��3b�R������L��|���Z�R�T�\.���`0؊D">$�N��S��l4���������z��!5V6 ��f!9��Ll
�d��ω*;��r��TҊ�[ޫ��3N��&%��&��[�EA�>D,�N�L�qI?>bC����Q:�~�޺\ׯ_����n���	�T
�$�͉���ME�Aj��S��J�Y�<I���'�� hx��<�收l��HnAk(
�K���	4z��1������+@�d"�F)�����h��^־\%p����{Չ�;]hE�"P�hp�&�Yp0��%�pU�s���Վk�h4h6�ѕ+W�Z����~��o�bq�I�Xb� .���y�~?8g�%�ɭl6������'O��ÇtrrB�ш�.r2\�"�3�N��7�s��ɕ�A�0�>��U�T���cˬ�u��[��$:�����2V�a��/�����K�UJ�|ϒ���~��+U�V�o���� ��l���SKί��z�ns;�T*���NW�^%˲����V:����q8�:5�Y����o?7C��8�J�|��W6www��nӳg�h<S�X�.����H���j�e�X(�����E�lY��:��lY������)�9��Qw�\�TuQs�e���E�����3X0�N)��Q�R!˲n��վ��P(tg6��v4�h�Z�]@�O�n� 3`Rh��I�`0��l���-�u�w��q��y�n:���������7�R�P<�	��[/���J�R[�a|�l6o|���(���`�#2T>��A�)�H�D��*�<-nU�y\��Z�^ߗ��P۵H���J��,�~@LdB�(lZI�CT���&�j5��j4��`�].��O(�ׄ    IDAT��n�?@����ns`@�(�LΑЪ�D��ɝ������{����V��a$�(��o޽{��>}ʟ��CʜD�V�X_DD�N�bȆ!Vక��3�V��\�tVĺ��)�]v �,M�Ix�ɂS���o%� I�|o��)�e�U��Z�n��eCFN��M�X��
�d���_F;�3�� �����e�666�C��n'��;��������D��d�����b��������_M��ݣ��C�V����l]8y���K����=�C��Q�X�
���a�E���]S<#��nM����)^��*�Qtf9��l6cJ\��%c�x<�V���n�T(�J��b����ʕ+�>�>	��8Ge�ý���h4b�־쒪`�c���ĻLt��6����v��h4���)��l�Ր�����_�T(�n�B��s��z�rU����������b
ذ�=k�۶CRȪ��y[D�y]���L"��-���J&Q0�F7O�9$�|>�Z-z��S,��_~�*��N,�����v����l6���hP���  �yP $Z�|��p�u~B�|��m"�~����h4��t:�(�Ln>y�������S>��XZ1ʖ�L��_I�S��B�ݦ��9���h���R�AT��r��$B&�x�hK�-'q{�UE(uS�Xrz @�!k$'�e�%�'YI�������k:�X���B��k�\
{��C{_M४ ڙ�锚�&�$������;��緓���\.w�X,�h(����~�T*}��dn|���tpp�1L�(�,P��Z�ڄ|:$�'$	�
&��'����e��vB\݊�e ǲ� ��[�u�ly#D�(��!� ����r���ǕJ�En��z�������`0�	U �q��H�8@�,�ઠ�c��j�.VyX�o�Jm!$R�e1��D���hȺ���퍍�ȅ������v�Z�D5�f�lH	*"�11��Ť#�_D.̋S�����\��5�k��8LTI�3���_G!~z�ף��#�������ޣ+W��D"�[�����CD̟�����T߻� 
��$WO:���ڵk�D��_��_[�T��P(t㫯��z�·%�|9E.[ǈPSA���M0�882���́�8}``J���&^Nv�҄�+�dw	G��r��3�t����ό��%�j{v>�S:���B"b���D"��d����t�v��6��>p�~��-߫��K,p�CZ*���˜X�lI��E��9�E�B��ce�x<No������R�t�P(�Y__����/�������ǡP��H$������{���ӧt||�S��H�c�j�z�
D�gs�$$� �\�pVD"
�O�K� �4�u$�@�U���H*�
J��G�dE,�gH�dK�3 �T��~��+���"7Y���C.�ܷ�A܍F�숉x!c���tk�鄺u(	�*��)�t�Af�Crǳ@ @�B����N6�}�/�N	��z��F�A�D�R���e�/�D�% ����ҭ�e:�n��+���P`R�%�G%"� )y�H$�'��(���L�S���tttD���T*���7�dw>���j�ͽ���@d�� ��>�mKI�0M���:d�N������w���[D�������cj��4�(�H�dA�:Sۮ��n�"��{F0j��:���(�&�\�	U�W�గ&r}���7 n�@�z���Q5���WX7jҖH$(���{P 	@p����j���5N�67�7���ŝ���0֪	���+Zg�����@���FTD݂v��1�T*ѯ�k�r��N*����x����ץRi����>}����?M&�7��8=x�����P(�֢�V=�XuGv���a��n�ޗ&5˞�y��^��e���s��z9ĤZ"�~x(h�{�@1�������E���������z������"�9��"�1�	�8�ີ~�x�R+��:A�yHXa"}8R����ѺŇ;�2l�����V��y���������z�{{{d�E*�JtrrB�F��$�pRϜ\]��}����uJ���]�V���tV�hIQ%�d�^m�ۑH���)ѓ'O�ٳgT*��7��mll�B!���t:�ߦin��.v�󉀠�8=C��v��~��?�񏷢���h��_|A���|OP,ɤ�����=�'cvj��}L�@�+�e���A+�-_y���ؠL&C�P�s��ʖ�Lp�\�4U���O8�p(L�A���H�'H��`�h��^��������x�5�X�ȥR) J�l6Y?��/\ ���u><<���Cz��=|��)Y����8��(Ȥ)��M�y!���œɄ������o~C׮]ۉ����eY������b�g��X[[�����������?J�R�_}����aT*�l�S�"��l{�F��XW��gs^R�B��:j�Ehb^P]/q�ˠ��Z��E��]��&:�z�� ��_d�]�pxk0|�F7э�9����(	�J7@���nL��r��Q���[%�^u_�������Y�a������ɭw7�6\�^g/�|>Ϻq�L�8���CJ&��F�~���1����(*8�^����{7DAz`�߃V �'���{k^�4a��hеk�h}}��r����v���O��������t���"E�Qv&�4��m�Z��@�{F��Fm�rn׻ﾻ����[~����|~㫯����c���X��ts��
�M*R 9�{,D�k#���Ce2z�7�׿�5��e�T��eGJ����H)�x<f�QX }��������f"�uҼc6��իWm���b��9O>cy� I��4���ݿ���NNN��&�4�Ӿ�M��8�E����m0��*�{<�@ @�~���
�eY��[oQ>���\*�.��ޮT*�yppp�����6m߻wo+~jƍ�w���ޞ�X�<���|fWP��Rs�����7x���,j�Z��;^:s��ˬ|/b
�v��I��n�^�������(?Uj�Z���)��S8�6M����9���{���`��L&C�ш�M&V<Q]�9�G���֭鴸�	��M���AU7��� ��#P$�D"A�L�����F�|��p8�9X�h6�<P���L&lG[���ų�!^�r�.Jnp�k�T'TX��0�/[U8h�խ��B2$��L��>?�<}��NNN(�J�������/����^{�_t�P(l�����x<�,
�L&9l6���v(��\T��ј#�g}������E0��e�v��Γ'On�|�Og�ٍ?��tttD����{���~8,��o�2<�^�֥R)��j����O2��W*�b	��ׯS�P���Q�=���j���<�B"��l�v�h�K�9���;p��=�%9�r���C��G>[u�H��>�L�|��l����M"OMp��ʃF"N��l��9��{.	$A�"�F���i�~�:����y���������]�����ݻwoѧDt��/����.
aƂdU�� 2��in;�� 5f��t5HB�Z��utC����E���9%6���"O~�ByH��x�������	��yJ�R�D��^��B�W0���=���<?�|A�J@G����2S��,Cud��4��0Z�ീ����D�����������L&��v(8��U�# �`�>�j�P/��Y��霨��׺�a4�![�@m嚖z��4�D�TK�o�h<���#��j���׿�5�ŝD"q��=JQT��Mg4�{i,�@���+<{�<a������o���V�Z��������/����t:��
�g�ĽF��&<R	B�9�;yP�vd>���ׯӫ����U�����R�����h$R�	�٦�(d�d�I"�N{GW��u����?�����1��R�P�Ra�rY�:�n��{�N�l6�ќ�6��<ؓ��ʂ���D�6�ɛo����_�*�����k���ߧ��=^�Ј8�N����8�.���dq����ŉˌ�����W��^7(�WI$��x9�(�_b8� w�K����iI</<�/���e4)����ʃS�(�,��t:,_$[0x�Ӂ��`0��_�J�Rw���G��h��l��a�
T<I$�������պ�"݆�&�nT��V�2�V��O)+B>��*?��k��ӽ�=�L&t��u�r��N,�U.�i8��Ǜ����{��q����k$ �.o��石�&��
|�7v���[ׯ_�t2���������]� ���#[Ij�]\ƒ/�������>�^e$�k׮�[o�E/���E
��*!g�b��0�(�䇩��T)P�j��bH�c�&Sb�3�`��BA&t�����=>�DL�|8�l6K�j������lR�ݶY�.k{qnS���(����B�G5��T��K��y睝���v4�l�������jDD��f�sϦ3^g�'*ʅg:�.�a�g0-I��r`�
�˴a�hr����X��a1J&���ɘ��T�@l�� ��	�_
��F��j�:�1R�8 r �s����j����+�P���$�r9~3R�	�$�[kkk/�����~{�?��?�F�����.'(>�D�K$�,�M����d�h.P%U*F�娇�O��^F�+�+�Ⓣ����D��4k���������!����T.����ǯ���Β�M˲6���A<���Q|�eY\���(�ܣ��ҭ��{ｷ�?��V�����jm~��wT��(��P8&�g��,!&H�-�]*X�C:�+9��V����������t��5�d2�
'QQ9\�r�e�|e��	?�ϮC(�v��>�m6]�,��/��۲� �luK3����H*uH>�:0��t{_'�f{:US8M�Ai���XO�~���i�lՊ_J2�ʕN����_�F�ѠV���C�Ba���R��V��7m{Z�&��{�����k�)���HyQ�/���Xf0�8��` H���5��)U@̡7MD�~�� w����o�|���FD�����P���|#���]4���I�m�����BPyWr��%�RL��~����ͣ��x<N�D�-�9�D"�C�$n�6hk�S��")&��E�j[��/]�$�|��%��*���(U��``�V�I�R�Do��U��ۿ�կv<�)UU�:gL��B!��n�ʃ��N����[o����MD�GGGtpp@���<�&m����r��$�|��VU'�^H��(��i��rL�@C5�PE�U�95���3���-5y�!�x�5*?'~'��Y�cY��*ib������ea7y��S2�t�,D�&A�:���P�����n��^�3�GE��W.�ۮ�����>}��o|���h4���
�t:����~�v;ZY\�7dwDʆIz�:pyF��#=eY�q�N�A]�:ICi %�8&���*
Q<��t�u:��:���{��V$�l6����m���dB�v۶.�ʌ:���e:-R�+����R�r�UV����)�h;����y���j4�mIy��rN�Y����Nh��`��p�*�-;%L�æ{YЩ2y�L�r"���^{����v:����r~���$��\V��		���a��!��f����߾���7P��z�� /�¥��ݟ�*|a�t�H ���.�Ш��-�Nj;_�ȪR�\�HR��U97U����ſ�X g��9�B�?�,T@a������R��dYG��'Z���4��I�,>U�>����GB�j�l{�/��d2;�=�U�T>�t:�?����6���g�f��3:�3��K#U�[-��˟��&�*#�K��L��Q��g��&������q�{���{�+
����LpA�Qe��������IkȿKN� �v�z���U��* �����\?;eu�_Ċ𳁞�.��	�:�48�
��%(^��^�"��WB&�2�����4��4�I����R�xZ�Ht�l�|�H�HJQZ�\L�(]�Z__�����o���OJ�����	�z=���������$��G�$ڲ�"bڍ2!C����a>$�������@Q`Jy��tJ�ɔ̀iSA�ɬD#A%�������}Ok+�JQ6��h4�kAv����j��S��@>/���ϴJ�۫NRQ�����^�5/���c�׭�߿�kccc����m�T�v�d2Y�4'���\WZA+Ek�V 贝u_w2S������U(UNÕ2���z�V؆�L��tik��x���8Y�H��yز\��uZL*r%ex @�u-e��H�G�W�D"�zQ]�
[���H$���vi2��i���l6����
Z�h�:�&|:3���u܂����$׋L^�4M�,�'9Q9����e���u,�=8���c�d2���F�Px�4M��|R�Yx��~��_T��H$bS� ʅ����h4z������[׮]����y:[J��dD�o�8��GC[�-+'���ʃ��p�C2)�1�t�ъ��z�ȥ�ǳ�s�!(��$UZ:� �dB�јF���[��h���LӤL&C�t���,�b�3��A�H���4������,�$u$�JQ�X���5j��ttt������Y��+f�}[�ť��L���*��eq��\|~�W<������K/ݸw�u�]N�L�I����p8|&NN�S��sCX��`Em�ʃwBМ���q���[������ ��F̔R�莘������n�/��]�`pk2�|`��x4&��ɵ��P����� 9&�N�9��zڣ�'�$�W"�҆T�H��V�r�����la
���`ІHIe ��=��A����S�^�Ѫ<�e(���upx������v3-�Y�#������rt���沷���������Y I���tT?+)�t��lG��Q�*�J`>����������`�=?�7l&B���-Y����B�g>�S�ۥv��4I��U�ݦ��������j�!ٕI�n��N�a0O��BA�Ў�@�]x�2���Fa $._b��Q]��?��6�����������y2�
�gY
�v�k��A�N�6��TQZ ��u1 ��2���!��^2� p�%N���`���/�*���������'�ht���dѕ�D(
�x2�Q��w��ݓɄ�4�Q�d'O��^Qy?�2�:ڊ�p�~�u'g��"�=�	�ݛP0į� ��.v�������2cs:�J��?m�un_�jG���7u������V���śU�5���L^\��|�w���sG����Rq�\ۍ��ո^V�;9���:Y)�}���aDH�^��&y�-����4��(��eY��d��*�Q'�#/��@���ޏD,�ء�	����������(A�px+|��f7��������8���G����=�O�b�Ϗd�K��h�C�=�J���� A����N�vww��ޭ��+���)Q�.V��IU�P�N�C����/��Ώi��z>�p�K���0*]@�ҕ ��ز�)�����r��4��7�)ѩ8�v�"�^k�9�s����իW�d2*��ԅyh�dBjǨBG�u�X>]�n8�0�����ZE�j�Z
ɍ��o�ƃ�������Ɔr5����~_ɉ�b�l@u}�딝?]K�L�D��qБIܻ���k{{��_|��o����&%���x�^�$^J\���]��,�4�y�C��s��e%������z�z�z�X]]���JnY�2f��#%WǳϮ1��e���T���p
��}Ƀ����َYផ��B�$�]�
եix��27lz<����n�p��n���p8D(R��,Nt% &	VA�,�٩����ŎZff����֩⠷�8YH!yY �	�ԞՇt�b����H$��x<�P"i6��'�2a�3�>�����"�����?����tss3yxx�f����h㫛����ϵ�O{�!QD�����|��X__G<G$�҆�[�h8    IDAT���f�H�RS� �	Lߒ�'?t�9�{��+������w��@&�|?Dai�l���XN�4(�?�P)sP����a�\.���L�`R�J{yV̐s�A.��0������.'���tX�^�D�DI[�����S�m4&�* �k�T�>D�����u�e=ɵ;�q�ˎӥ,������gw��n+�V�-��Ԁ�Md�.�<E�DrIG9�cJ�F~���}�E��͐?&�l%�C&rC�����v��mf#�r�کv��"˪-,)˔������Uo��)5�J��֯Y������Қ���-������J�����r��@K.���z�a�� �x�mv��U��V�����t:�B(��0C%�DNtɲ�d2�<�v�T��!ҡ-
!����`gg?��Oq��}��q�K�QE�L��~�BwH��R�V���xb�⩮��7K�L��C�D�h�{e��~^J�I����ass�pX=?�{�a�#rr�N��\6��Y򂺪�+4�lG��l1�̐�W���Ȼ|}��ǟ��gOWVV���p^��fП60��t>�OR�N�UY%�VE�U���=�"y��>fq�u�~v�y�er~H�9�pw-��^g��ݙ��2FJ���s��p�,��ҩr�I��?�uB&KL�����_:�'��3�
yҺ�Y�%�n�n�0u�.O�N⠿O���uY��X��e2"T�����rئ�j��v#����=]___��v9Qx]vJ&�2�%Ř0�z=�1�F����+?u8����$���n�U����� y�D��dBh���\Uv!��(��0b�"���0�{�=<|�~�!��8|>�UC>CY��
U"]䢛�E�JOV�M�5/�xeKNꛚi�I����2P�G�i��H3ѩc|/�O�� �j�^gggj n'S�ް���H$�V�5E���y}x�C��}�\ ����F#d2T�U�vUgf<�x�9ɵ�w��
3��t%���l���� A䞳B����>�����'�����ݵ��n�Ŋ�<�t���.A30L��#��l�������h��+�w��`�.%���H���F�"�"�Ȕ�,E�E��y�S& v$g��]��������s�w�A�J�����#�`}}���7*���K�k����� �,�nd� ׃NQ�x<K�(���?��o~�4�%��0F���J"yHP�P��+~$_��]8�G}�P���m�b1EQ����j~�Ҷ5�82K�f���!S�=�~7����m�Y�����,2��ݻ�H$�z�p��$$���|���������{l�N�	�ƫD�$י�L�%�\:P�P�h4�4����z��|.�K�9<lF���`'�8��L�Y_�:�V&�V��2�̬@� 酟�}�<������v�:G��Z��B�TI���0�8ϳh.rn��q�kG��P�Lp%J�v	a�wQ���z��M�'� �f���SNtxft�E�]f�t:�U�L�<7��5{/����V�.,/9�Tq{ܘ`�lF��0��ְ��r�$��n����T�����h4P�TT�+��R��5)��=�v�a��^�-k��b1g��R���a����[�9H��Y�L&FLn�������1<x����Ca5���E���*���1}�\�e\�$����D���ԭ
�F��L&�L&��b{{�hT�=�`|���@ ��3���nW��1��9mH ���z�D�$���$*'���������׿~��x��V�`��b��|�Yj 0icg��B�T����7MXo�?��杇RaD�2�eaĄ��T:ށp˹|>ߘ��H0�HgF3$�̝N�WlY��C��.$&T�ߺ>��M*�qny1�1�e���C�)�^��^~�CUfJVɦ�J~^��Δ�n���3�����7��	�#nJ�8E�t:�v���ڂ������.,õ����f���nWI?q�ȢPrr��!�?i�� o�+^Ƶ����D���BNy���!+v�$�I�s�M�@ |������O��>� �X�h����^W"��7蒆rm3AZ���Z����V\�Y�Wq�C>���C|8�P( ��!�����������Q�SIݑ	#)�+�*vnI��7�Ǣ����w�jD��E'3�kmm���t��z+��᳖ٝ]"�f ��𘼷:�����F��
�:�֛�y堭�o,��0��@H���{����"�N�wi9-iR�M8��y�ϗ���uO>'�� >/H�ÒJVѲ�ҥ�h~�r�����/��R0D Phz4UϕI�zV�zpГ ���mҫ}Y�_sVҥ�!+�0�5+�	V�D������Ҙ������
�0�L�>|���<�] �N��H$��)�w+���N��t ��A��P(��`0�? ����\������G��Ip�\�z�o�ךM�2�]]]���~���'?�	b��zv��_�֜���oEw��pv:Z���y��aJ�����������A>�j�P,�N�������lmm!
��H&fn`LjC$J�U�K�C��	�	��������K�-]1�]�VVV`"��:������t�1uN��.�i&�h��澔��vb�M�/��7�}�S�AU�����9 ɻ� ������׮��Lr��[v���x��iJ%sH�mf��V�դ�.�KoJD�����KH��ǔ��nl�g�������
T7��1����gf��f�^��V��đ��Y��
Q�F������9\����?ͦ�5��ҡ-�[���
�T�-u{�ܞk�c��%q~��h�x�P��#��LRa�Mih. 9�f��Mڒ��VS�v~�UR���%H��F����sD"�v����H�b�!Y�QM������ճPl���� ��K�i9���;?���!*�/�����)��=��U6���v��d3[[f�;R"�^��R�(�A�8p�T���@J��u�k8��f���<�������E�^h�����զ����|2����h4Z�������"��O�N�@��.E�g�^o�:f׭L�����-�U@4���	ˤR��"� ��'��*9�f:�\c>�^��0�֤Ԉ��UA!�`�D_%�����x���p���Z���)7�������K��"���f��������X,N�����yp[u��Ŭ��y\H3�\�ۍF����#U@U*���{��W*:��IT�����
������?�,������W�K��Y��!&��`�ڔdt�%����4Mp)����˄��D�:̨�շ����ļ�&���j���*���T7����J�Rs��%�����6����h�\��IU�v 1�w�m�ԦT��Z�4d����LY���i�[^l�0ђ-nR
����7Z���NR7�2s*[4ș% ���US��m$/����4p9]���{o���-z��d�Z�eK�(9�<�e��ʺ��O"�L<[���n���֝�P&�MI:��ť=���( װa��r8::��h�kpݳ8�e�Z���<���"�ɠ�n��.-�c;�����Y?o���u���Q,�j�P.�Q(p��}�b�)\)M'Q��m�Z(
8;;S�^�z� �pș+DP�vO�I�럯�'�?�����7i!+-+m��a�����.�d���겭{�!��(r��;��@��(�(�}�
�*��D���aTKË���~O�rȕόZϲ;�Ō������m�Y!5��R/Q�nc�PN�R3Q?|ﮛ_�nw�n�1����t�l6Q�ק7�ID�ݲ�^5C����eT�i�Yi%�%h~�_��bM�O�AGn����)W��p�ȿ�v�S�[&�V ߟY� �9�#˟?<<|������֝�А;E=\"~�2�{��>�Bx8��h��� ���V?��O�������5��d2���óg�������)��y��j���B��e��_;�����p8D�TB�XD6�Ž{��Ŧ�^y���h �a�T*���*��}�)��阹�d[ꖚ���.�bA�;��:Y�L��ʃ��ZR<�(%v;o˺���:���r@�JK����] T�������-�˿�����uy5�1/].�d>BT��~�~����$�d�׭/n��Ѭ��*s&���J�1C%�8���J�R2�J�^\\��"7q�^G�TB��V+�+ɝ�ۼf~�v��YI�j���1���!nv�\�R�suuU)K���p3�B!8N�}����b�b$��p8���t�$]f��C��;���IJ|�� �?�_�	��Wj4w�]d�Y5���v�j�`��2��A�0�J����k�z�
�t:Sh�cv��N1fW�&�Ƭ"�ϣ��#�ϣ^�#Nq9�x�zq%���Α��֓V��g�ғ[�q��&�+=�w��c���5ӭ�y�����ں��.Ӵ��������W��;`2b���0ΰ���O,��nwr8��Kpop������n*�RfS�C�������T9cd��g�)�kW�VˍoP���Ái�t��޺e���x�l�����h�Zh�Z��SV��`�Z�w^pZt�kށo��f����=f��V��lE�/�?.�'8�N8G�˒�x�����v��F��
���t����v��H"Y�~�z��g{%<�D�r"\WQ�H T*4�M��[�����Qi��tP�T�������tTl���E�y	�gx���O/�/�2�[
���x��!%��4��3�\�yq�����$�3fZ��.Z��+�>��;�{���IS�>���zR ��l:��.��#f�Tf�,��d�+;̤��|~���b� w׍s�ϗ�C�R�ϰ���b�32��D�W����l��A���T�#٢��������h<ͯ#C������tF���&��%����lmm!��C��l�!�ow��evP����i�����z!y��N�A_utĔ�-'��k��{u�o�����`0HR����J����I�.���ǡ7&攋[���&���|f�o���v��G^V��C�Z�����M�f ��!�ו�-�y��j��dMZ�f�� ����rm06H�JG���Bz2`&�g��8�R��Ĵ��Ҳ�ݖ^��f���|�~W/�'}��)��6=�"�2ԑ�yq]����;�o3ɝu>� ח�V$��l6�h4�#
�8��t���z��B�w���w(�W�^���))G�v��aN��#i
$��iw�VK��7��������}%�.�Sg!�����7�M��v� ��x<o2.�p8|�nq5�M������P_�Z��p>�O�`�ZMM@3�0�����y�GVT�Y�K�����og\}}+T�ha<�a�D�-+�&��ɯ���-����ذ����������	.bm�I*ݣ����;�y'-`�{����3����ч�$�ǎ�l'JC�4����(W�(W�j�LJ�P7���D��Ūu���jj�`�k��-$R�"���k�y�eWDv�f��r.���(�>�$M$8�T���p`2�6k���DQ����L�t�z��&�(��2X�(�u9�2&�	Px[�B9�zE/��(V��_�#�<Y�p�\�JU�������`���p�+�J���,�ժ�I"�Ȕ�4�*"�:����=v��xR��gM�-rn<��Ȋ�I�tW�&eb��t`�݄�-.�0��R�0L&�A�o^��a�X,��m��T�ּ�ЊV2K�hQi0=h�3��1C����dr)_�v)��tK$W&����o2�܈��p8��gd�����h4�l�`��� �ē��8�,i.�#(�[�̌�8���);V��dK��TR�K�7��R��Z�,�w��9�3��>Ob�g&�h���C%�V�q-P"o0�ǔ� ���ϢG��	�n�����d^br��1Q-`vVeAn��Ћ>;�^.�e[vҫw��D��j]R&q�/�����a8�N��m��ux<������������n�P@��F4E8�RK�Ů%U�x^P��.K�=�LFrz���w^ˌ�V��UK
]���������˵���~���}W-x��������a�0�s�(�y��f���5�f�f��d�f��zp����q���ަ���f"�*a���qN��N&8N��)
�l���+���`0ZV�W�3��V��"�Cڐ�F\��j�Luer+�xOe;P�)��)�6����h6pg�n�Ikg�.�Zf�f%����7�ϓ�3Kn�]}�D4|����M�u��gg��]���{t�f��HgC�f��,�um]�^/����w��7K���3�[�v�����v��	i��SQ,�����p8w`��gģn��,

t���R^~�_�X���t:�t:
ѵ����h^�7��ܠ6�,����˹9ɩ`2Ńj2�$���;���h���p8D0T�M�׫&��K$��j��h4���a��I����l%'��j�P��x��?���QW�w�+���p����-��v)^����n��v��f�95�R# �A"b>Gb�߯zV��0�l�.�j��cV�D�%���Kt�	ף�?:�P>Cѕ��P&3�v��N1g'y��f�9�n�J�����[v�,���卸0y�����9�S<�0�iw��]p@�V�M&�L�$�|jF�9��p�i�KT���|�y�9YQ[�	��~�{�z�"u�V��0���Ou���Hn�ZE�P����n�T�]<��Ul\ɓ����|�~_Q�~����H^.���<��&�z��h`e�C&�<���1��&j���T�͡4�6^��<��r�ݡ��]�\n�h4�	��p:T+��>��D�������$�"�ĳ�y�6���J��VJ�Xغ�5 Ż��u��p��p9]S�%��N��z��߿��;�^�����g���*��F���^����߯�%������.�.�h�Ph�+$:�]���á�"���D�d��	�Qv�7;kt^�N�bY	�"�T�:3���,�}��t>��8$���Z�*	R���0�9 �#��V��[D���)��a��"*	dp�{8��pO��(ʠ�=�C�kl���Z��V� Y�R&�	:�J����gL'��ǥJ��N����jw`�} �Q��IV*8�ND�QD"�ˮ��:������k�}ڂ��?�r�d!qɃ��1%�[��@�TB�VSo��τ��n7��6J�z�^�����-	����yr4���u���>Ղᢨ��V�h4
��V��V�h�ZS�G.�Y��,���"):�d��V�ZݖS���I���a�s���Z%g��"yq�=��n��=�r������mw�S�D*$($e2ݞg+�^2���"G~�W�����|>�N��@ p���\3N���e<�R��Q��cv����s���f-�E�۠�������U��������j �|��!9��ɔ.[��=�C���|2�R��[vG�f��)�����hx-�Ϯ��z���<�߬Sb����e�׿�4���ut��)$q2�4�!]�?�j�hM����4y��̾NNN��j�q.�S�~���|>�=��|.���ΠB��՚rp�v����O#3�%t,+w��V�C�zR�5
]'���D��l���-p��h8&��@�U��U��I�D$��R�	��E�f�z�3��=�6�.@n6��/��*��_��5��fxHH!|r\Y�q抗�Wk0����d�әR`�^^�BdVo�J�\y0.��v���q��LE	����<��d�3H���J�Pw��،�9+@�:�穋��Z6��6~�nm���P�bL�~2��~�EMp�q#����������j8:]IvGY<�y��U�ƣ)W/�bCw��Kۙ��6�\�3F��3�a\��.���B��U�#�
�~?��.����h4��V��]2�5#Y*�0��D�DT��󌉮# z+ר����v���J��Ʌ����`�k.��D�x0�}����x<�X,�@ 0�6�L&h-T*�F��b�xW٬�����J�2�k�}�x<��X__���6��	S	��B�fq���~�w��<�W?H偨[��A;�$K�G j3�<���n7� ��gϞ�^���p���`�
��_R�KFDm0��Jb�zq�[    IDAT��?;;K�j��B� �Ӊ��5u�:NS�χ�?�P(�`08%š3�):�7+)���uŉyE�<��y�M�J��bW�`�d��T�ם����k-)A<�d�O���*&9�N8������r����&<VVV��>4%>��%*�8�*�z�P��,�/�6�7MF���#/�F��G��PJB���I�BE����D�ZE*�B��x�J��r��C��x|~~�B��^��ޙ3N&5�C�R��L�n��s�b����������LJtO���Jr�������H<�����s8jzZN`��ut:�d�Ѹә�q5��G�v;Y��Tr�;���G��Pj�蒚����l��g%��]"U���#�2����<�س����,���}$����	�Uk+i�m���4�`;O����T�`��=,�%�d�,�f����~n�X[[SCl��?��P�<��h�TT�*�̒�y����l��ӭ��@ج.�]I=��ӊ>K6춨�Σ5{62�R�a��AƮ�T�g�2ԥ�d1
������=O��n��M6x<�>ǋ	�,�|q�1F�P�U�~%�@7o�J.oS�-�5�B����K0�yN��C�P@6�E8��ʊ��:�U���6��4vvv��`���kq���G�a$S���*VWWUn�.r�g4�� ��`�F�6+n���SG6�I�qy�r���a(�����PC7��H9Eq��\.�z=\q��h
6��b��8�ϣ��)�'0&[l�B!�B!�F#\\\�*Vʡ�;D�$�*p�vJ}��i'I0s��I�$�ޓ���'��t�]�V0P,��z��7�������=��'�Ӽ��}�BFڬZ�PK��m�l6�<??L�ە����"�{'�d;�45%2.]��U��7��ҕ��y���2y�˺v��ՠ��>Ytʵ:��8O���r�i���;�[�j�F�z]Y�˽¿�4�)��J��l=�6� ��\+�آ����K�C�2�N�Su0)���d�ս� �L���8��e`<?�����_��_�x��\_�~�m"��?N�Rh�Z��|�F�*�k�뚱�n��e��f�V�T@2���yǼv�\ L�(*�vo��F.�C�ZU������pN.�C���=;;K�-����Q��L�EةmK)�@ ��h4�x<�6q�لaSS�2X�6��es�f8��A$M&��{׭��=��ӿ�>u�.��-�b��z�Ή[����Kl�PơM&�RnKZ��ܺe��v����� ���< $G��`�`��?]��g�� �+��ڗ:�w�Xx[�m����ˌKou��LI͓�(��5��Kz�mجV�����2�a�M/`��0+�F�w��J����:���\��9�8��K��E�VC*����9J����.)1�F��K�J5�r��T*�;�� ?����R��<==E����ʊR�ч���!F�p(��Z�*����U�iVV�f��\���ʤkR��E�PD�TR�E���e�ʫ8�h4����$����r�N��8�ɠZ��{�̤�A���h�F�r�<�)����&Ne���R;��Y�D��8.�N��!���Lc0A�yB2���\�P~�_���~�����ܵ,5p����J>1��n�kf9,[�7��J��ggg�����b��r$c�v)9�v[i0�#�|\vq8�,a�ɝ�Z|���f���o�C8k��`3�i��q}pJ�I���QT�)#�����_&��m�Zp��ʍR)��c���w:0���y�d!��%�v������~�Kv�8��t2�.��
�r��:���K)1"���f�g����j�z7pvu����b1qzz��2766����$��g���V� ,���]sKw���1�L�n��4�8�S�V�N�Q.����d�"
�N�����a<�f�w��v���G�j5Y,��']r ;��j���(
H���d2�t:S|9���n�c�`�#�1/9�;�&y�V�-L��p0尧#ADJ�Ǖ�]��7�qW�x�0�'�|>9/����~����?z�1�+H>�-أR��L�R�L&���X__W��Zr��ݮ��z��j9x�.�|f�K���3���w8�\k+'4S��[�����
�.;s�φj/2�5d&:+��\�f����urr��O��z��n#�������db'JRҤ;�L^����	�M;}���M��E~Nw��)R��D�RA�\F��T`C��UN�@�2w�\�T*8:>�����/�����+������?�t��R� L�{�^8��:�8|�p8�n�=�h�,��v�Y��j�r�P2�mr�Y���\NM�y�^5�/'^�z'''�T*�;)������t:������HM���g+��	���bGGG8>>F�\V�9��=�n �[A��W�8��$��L��<�� j��}��&Q\�/L%��`��*��T
�b�v�o��x�K}P39�R2M&��(�~�:Q(���c{{���J9�����*L&0��0M)B���Zn�ZSç|6f�֛�af�o���DJ�P���)���Dv^b.ٲ4n���'pzr��ܻ���j�G�F=Q(�����s��wvt��U+H	�3ܓf�[>?ݑn�3��F^f����$� @ݟN��Z��R�����K ��=��ױ���Ӊt*�t:�l4O����&��f�U*���T*}�J�����Ű���DF���pw8�z��������f�J���t0GD�^��0�7����.21KjFʅ��v����v����`0P�f�n�[�R>��~�\WT��d�.�����`0xbF��h cssS�1��P���C$A,���D.������4�B8�/���>��܋ vQ`}����C.W_D �ƣ�u�����l�����T����prr�V���^�'��O�.�Yrkv�K�SW~�M�{vv��v�O�HV*��a<x� �x�� �Z�V�A�^�#��r�Tr���GȻ�ɺZ��h�e�(ٲ�Y��y���Br;k��o��<[&Kf	�<c�w1�}��U�Z�>�f�����F�X]]U�=U�Ot�&�ló�B��n �ӷ��V;]���p�"�Ҷ��l�T*��R�B!սc�<+��R��/^ ��%&�ɓ|>�w��'������}�0x�^���aeeE�XIi@��	����g0����.��Z��\Wgu���s��vZz���I�}>��Z<��zr8ꍇB!ܻw�H�|�B!�����Q�T*����O2�L�����pX�U�UT*%��q��}<x� ����f��d2p8*`���<�S8�M�Z�ј�9�\��8�R���%���F$��ue9{�eGo�He�K1u�˅h�Җ�P( ��$,�|�`�^�4Cru;J�}`D�T7��a_���r����VWWq��=5p!�|�l��i^�M#'����AE�I�E�K3:�"���v�BxӤ�n|��<Z}�,S���7�"�R����<�Ɠ��3���%���dEZ����Ej^�ZM��}eiJ��U�t��Fҙ�!���Q�� Ǭ�+c�'�ơoQ���\F�#��F �*�M�ׯ�� �cee~��+���x<F�T���>����l������M�����^�I�RI^u��v����;JVz<e�;Q.�Q*���vU�+�F�a�8��[F��D�t�$ɣm4h4�����P���������x<�h4�80\T;;;�w�*�
�?�����_|���5���j=*�J�W�^��n#���r��j!�������%:������M.B�>�1 �%}���O+��������ڜe�0��F�	��h��h6�(�˨��SH����u��;���9DN%�DD=
bkkn����8>>N���'�7`��O&�)���$B�l�V@��	��s^���/�����������)�e���1n">�O���e�R)���)�>_�,�ٱ�Z��^��)�d�{�����ì�_4��*�vHn+�oɕ'���/���X���H�&SMD��w!�g��d�^R*��b~����l�*�����	.9�rj�����#�����Ɂכ&����y��$W?�8�ȸšl���j5L&��˹9��yN��J%|���H�ӉF���������r�D��x���GGG*�����S���#�D"�L&��r8==E�VS���r���^��V����x�
΋�&�Mɶ�mT*�� ��T����t��x�D��j;9�u@K���rr8>�{�{��y"��?>??G�����������qqq���s��e����Ot-�Nc�TJ�'�B��-�(���w?v�f7h��Kf���h4P���-���קZY�_o2�(��p8T���G.�C.�K�'{{{j=�J�d8�u�݊�#�T���~�
��gxOi� 9�W�����"���ӧ�\.�$��&;���8B��52M��Rr�S�kkkJ'w<_N��{���p���x�������r}������2�,QA��׾�����0�����z�2��$�.�D;�>w�\O߅8_.�e2���ŅB��b�����S�*����iLL���wuֺ�s��������e�%�{J��p���(
h�Zo w,�x.��alll ���t�V�����8::J��'ϟ?���,����R�����<���s\\\ ���\YY�2����h4R�y0T9���J��J��^/��.*��Jne�kG	�m֎����	��~�JE�W�~?��K�\.���3���`mm���ʘ�H�a���ja]\\ �%�������_��G?��U>==M\\\<I�R�l6���U��qE��* RNt�-�Z����}|����r3j�h�.rH�ղ��f�W;�l�3��V� ��de���nY$��f0�)�t�n7��<���0|������_>|�����x��t&Y��G�P���`�+M��	n��y������7Y*��x��q*�J��elmm!����5��H�>�BG*��\.���Ǫ���N�0�׽�5k8���3Ͼ|������4!^���m$�N�P{��4���+\c<����x&�������;M}�嗉T*�8�N��ncuuU�g��>��K^�p4|�� �Z�v�H�r	�d0T��)�|�y�Bή}�w�6�~�x����H�ӊ�@e�ӹ�1���i������}
|��'�?����ׯ�ӟ�������%*�ʓL&����C�P������:�� �~�*��E���*666�v�Q(p||���t�]E����(�J���h4o���u����M��R��z(����k��xP�V���s��aD�Q�����e�V�x4�a�7�����F899���N<x��I6���{�~�I�7�|����xrvv�8<<���Q�Yr�h������P(�����~�����aB��oM�(f��~��d�,��F�n�D����6\��{'��E��تׁp��{�}J��qi�+[2�j���	���������L&��x���d�+7���a�@ �n��|����6��o��[.��r�W�T*qvv�L&�ĺ9�b�ek�垲_��<��J�1n�ݮB�tUY��յ�uf��m�X9�-�w���Y VSVB����Ik�/�=�aY� �m����������}��'�����C�Z�>)�ˉV��f+�n��#l��
.:5J�q��DMQ��˲��جkd����ى�V`�M��9}�Ɂ:�7v�2���(��(>|�:��9��z�+G:�2�2����p8|����_~�נ�+��$[�֣L&����"����j���4�hT�c)���v����������AT*\\\�EgO&�	��&��<�ŢJ�	�H��YE�{YAL�8��h4Tf�ĪZ����kkk�w�r�⦭�jO��y�u8??���M8�|�P�ۓ��D.�{r||�888���PS��z�b�V.������F1��N����boo�rYD)&������p7k}�%��A�uÇY��D�a5�V+++oXXN&x�L�Z�kr�4J��	&h-8��rc���}
x��D4��z�ި�h(����Bt����C$|=�B�.!�CTh�����%qvv�$��%�����yD�Qlnn*��[�Ӂ�?�	�Ldd���)����Juɯ�����V��,��s��������9�~I����h0VI�>�|�!�R#���N����z���"��'k�ڣ�����|>Q�VP���Ur��E��g����3E�>�n�^/��!�*�
Z����V�Vg��&=����r\rk����Ei�V���
���bX]]Us�fSQHH� ���"�J!�J�R����$~��?���/������lΒ���F�W�B!qxx���}4�MEӈD"Jۚ�*�1�0�h6�H��8;;SfU\Ln+��*���n<s[��������m4�5\������q����W������{�aeeE9��"f�b8&vvv����?��.���o�\�I:�N���`4)�dʰ5�M�&Y[[���VVVTY.����<��BAmB>"�f�<ݬt�AW �W��MR��#�i�ie����w��ƣ7ֻ�q�����F�����D(�D��b.+s�����<��B���ьsG��Ø��H���%̮R����z�������'��4��&"���8��  ���F�G�S�L2��4�`��z�VS�"����� ݶ�p;��a�s����.ɼ�j��ƚ��E�4�>)��x<t�]�R)�b�����^��~�m�P(��R�$�٬�����.S�!Yh��K�BvMȇ�lg�TR���s�c���j����᷵���������m���ceeE9.޿^�W�S���@ �X,�f:J����?���'���_���m4��O>���f�����
�ķ�~�T*��h���U5[A���p���8P
�����p8�n��L&���Sd2E��h5[((

����z��ep�[7]�<�x���5��~�7�
®�kx���譯�cuuU%�X��f����CL&���������_��'?��$��^�J
�'��牓��C��q����V:���|>�T[��� �J����8>>VI����x�ڇ��N���̂��d�L-�,x.����CO4- �VE���N0e!�p;��8U��l���)������j�t:�r9�z=U��aeD!�Q����|�R����#��W�
�B���<���[�V2�N��U,SRE\s|_�f�K:�����ˁ�j��|>�j�:���J�c,�֘�ahe8��w޾�R&Y���/3� �BZ�,�x��5o���k��H���$����I���A�V�=�f����t:Eٓ�|�I�1���C&�������D��Qr�T/�7X�Hw�N�"�&����fT}?�d��c.�Sn�DrI�j�ZJm!
)ɫ�x���u�b1T�Ud2<{��f3	 9�L�6~����OtS�T�Z�>I�R�gϞ���^�����#Յ@B'�(cj�W*�������ZMugZ���"�<��>�~�T�Ϡ��Y\t�[��"af�pi[����y������J�^�|�`0����g�F����Q<!rL�б�j4x��:�N"�?�����_����;����׿N���=)
	.���-%CmV�(�:��v'''x��9������	�,�T̾g�akDn��-ܤ���DG�s�`��18~�G����:�%!�q��ݮ:@����� �	�v4׹t$����o~N]�LN����v��p��vO�����D�\�U��H�e4��t:��,�;�VL:*��V���~��b��R��4�R�ܬſH2g��]�����V����$ķ�0���HR���6��Q�݉>�-/)%$�B��}>z�����l6��W����~fw�rY��ׯ��V�����c"��nW�`�RJ��4p�&�<�T#_v���B*�/
(��0�$X���3��N;CʳΛ�$�V�kŻ��1y\Q#�p8���CE���'�l6Q�וZ��榚/�T*�d2�f��ӟ��B�v�    IDAT$?���������>��z�*���}��׏{�^����L�[[[���D,S]J�7ɉ���X��acs.��j�����߿T��@�;�J�jU�A�R��>��bӃ�M�������a�X,*�%�������?���N��d2jғ��x�����1z�^"���믿�����g~��;����^�T*=:>>~����l�pXU�S6�W-+Z�2��H#���ٳgx��9���
j��HpQ�ǎ4Ҽ�3oz�6��.lz���l6�l6��77���x�W&|D���f�t:�Z�N�:�y�ih�xSsq4)��;+f��!��6��k����6��+�N���w{�^�P(�Z�b8"�!*���{����/�4I�p��f�bQ�0��5��I90��M��֘no�*����l4��\�m��� ����Zڅ��.�tM�`0��H�Хy��ԝ�� �$�nw��n?������������᭝W<��t:=8;;����s�(�B!E��>#��\N�T1�x�p��j3YeA���/e�<^�zttD��)�%;��,��&���y>��@iH�jƫr����.�?�я����H$���m9�K����5<|�<������W_��>���)��_�%Q��~��W_=�����B��������\.'������� �N��j����Z+n�������PT��55\�sr8"
ass^��\{{{x��JŒ<nw�SF����=_П��ɰU_4���Uv}��F8;;SS�?�����T�DD��S�J�Ad0$�^or2�<>::�m(�l{{�{��f��d��|��f���d>�G��T�m0�d2Q��)	kkk�%R��U�:<<D��R�K"$fF�~�Y�P�Y��m��ڟ��g��Y%-�^O�W��e�k���V����������q������S��:��ס�
��h4��ܕ�+b"�Dr�8��F��n�^�4��!���0�M�F�L�`0�j;��4I����x<�x4���Jn����*5	���-ZY�����E�˦O,:���Th03��{X���~&J˵Ƣ��/��,��c��t���^�7���������?�۵����{･�/_�L
�_�j�D�RA�\F�р��F<W��.C��i���p�1�>)���w��C�sI�"2�D9f�Y4��7Z�zG�&2u7킼�u��j�nyLաl6���}E��D"��ں,.�.��9ۂ���V��q��~��O&�R)��m|��Gɏ>�(����?=88�m ������N󗣣�d��y��d�j�d:�F�ZU�>R�vcc�����'�ՓjWR �!�+���c���V����`0�{"���:v��E�*Xv5EN�h4���E$Q��h��o�U��/~���Ft'�N���!� �V���0#iFr%�����~����K蟉m*�z�h4�'''����x<���
VVV:A�Ln#������(���f�x��%���Q.�̓�L��䝕p�Ez�M�����mQ[%�v)�W�8�|>x<��������T�Oɧ�CX����3�>���d{8�0űk�Z8;;����.�J�
��MJ�m� Kjk����%*���L&p��
��xw>�W�o�Z{."=4� ���t��]���u��v?�n�r�.9�>��P�Ç�jIC~��>�uJ�����]r2�$��������~��W��+<��ؘ�h\\\$��n��q�u:�q>���v��\.��Bh�����UZ�ʸ N�����n�n�N�S���H��,Ѝ�%�Z��^�Ll5�� �s�K
�U8K>l�b�m��E��E~��ݱ��d�҃T������v��Z�����Z
���{��0!�͢Z����������Inmm%���㯾��i ����>\z�{5P��h4F�Ri|vv������r(�S���OS�ۍ~�J� ��y�Ӆ�zXI�V�U�ܦR)ՙ�63�-%5oQU��Cfo#�ꋛ ے���j������J[�?�G�b1����
����P\E J��"��#�J��Ç�n���/���i,��|������^ ����F��r��8<<���9�ݮrv�Ѯv���P����3�ǃz����s���D)&�#���p��״
�V�aV6�V��V�j�8Xf�	b�ZU�;�����3rG�d��Wr�dA&�Dat�te�*�/�{���dqâ��r9��������T[����V�	L���Ǔ1�'�<����:��T�V��t�ef�0/31�z]+;�ժ_$v.+�z�yŅ�!7��e��K���=v5�p�J���1�0r�����ظo$u�<A�#W�Q2&�ͦ���L&�~���OC��S��I~f��_\\���$���VK�윅B!uxK9<��!/�������x���r�UusCGC���V�RL�v:��u���!�N�0U$�9I�Oj��DJR_����f�/;H�0�_.�_F��N��v|��z�Ӊh4���Ձ�aP�XT�A�c9|����b*��ׯ_��� �pW�������4�;��+��p8tM&�����Mj���n��\_�j��b��\.��Ϥl�e��]�c�����������6����p8����������s'��y#���f���A�n���ϛHm�P(�t��?�^��Z��O>�?�я����2�L&����@���t
�j%�F�WF��~����px�m(�׳gϒ�R��˗/����ŅJ8b��
���a�BU	�\���|>T�U�ŋ888P�-]���8�M�,)��ٲ�*[��Y%�2P���R�(�/�߯l��N'<^����!�"<l$�I	2�-�J�G�*
����[���&[�Dz�^�R����J�������
9��ht�`;��rs�I���H�RH�Ө������5p����A���ߵز��<4k�L�"�Sf�f�@p��HZ�,���J4�8�Z�7f���*$DO�ͥ�(����ڳ�p��8�v���aL����uj}R�H�R��d�E�O�f���@�_8�N�~8�@0T54 b�-�	
���k'uJ�GH�@�����n�awH��@����k��f㙚J���n�۸�>"��Bh}>�ͦrt�T*p��Je!������ￏR��t:���ꍺ�{��5VWW�������H��u�B!t:�d8v�B!�������|N>C�o�7�^��v�=~������K����^��H�w�.g@���aa�� ���B�P���	^�~���St�]%0�h4�{cwY_��ք�����$�Z��H$�^���������e���ŋ�*xgg�H���J�RB����S(pqq�`0�V~rcc#�n����=�F�����mNѲP��G�\n|~~��j���L�nW颒ŅC4�����t:�D���㣣#|��8::RF�#'7nf�n]VB�V���</��z2����j���x��Fe ��&\�l��a34Y�qe�J��TH��� 9�R6I�}a�b~��l*���V�<���/��p8�D��A���V��T*���d2��'�m�`ߴpY&Jz[]��ꀶ��/�n�^eRif.[�\w,��En)�~��m�5��*'�O�hy�s���U)eGf�˥�^f%�܏:�B*�0��I�~��K���$�e3�@�ܗ���jU%�|��F�T
�b�r�ZMь$g��JN��Beo2�._Cv�̾W7�����N��.y��8�#�r�$�L&��r�L&*Q�d�����ښ2�a��s�j:��� �X;��i2�*�
��*��~���x�����|	��D��V8�΁瓓��m��)-I�q}}���p�\��'�$�E�?�.���,@�"���C!�ˡ������v�	���fF�('���n�jH�|}~ ���n�����˩Ej��Z-�����ￏX,����čh���$�x<F�XT�puu5�����j�~��ٳ�kkkK�^,���p�[(GGG���8Y�TP,Q��T@��|
��ly��h����@M�j����=Ź���+��������dG�j-�j[�:���$G׀��t:U@b���z�wMO{���5(�_�~��K��	.���B�8��'����V�(+mz1������Q�H��2�/M/F�jqz<�]n�Uk��(�H�R�d2��jS��:Mc��h���Mg�6��NwmQ��e�G��ɶ���)	ү��|M:z1)��ev �V���Ɣ&�N��Pn����u{S�#��"�V���P&2���0�C3�]�eKҐ\.���Bn��#J�-����[���:�~���M����)���i'[Y��� ��}�P@�^W4��x�x<��������j)�ov'Ha�>�����>_�VSϋ<���!��ϕ�9-��y)�r2O�g��5�-�����������>j��:/��z�y2�LH��x���� �B.�����\�T�fPd��Zf9���̬\���,����E�����-�~�r9�����j��j�O>��ￏ��U|��Gʭ���a�6�W�ְ�h�\.�����A��%��`�J���?��O�~���^�0�I
Ih4����]�˕�M�^G�RQ.2�`PQ2�~?���K�]˅˅��������2������_#�N�R����(N��%,B�6��.�^��̵c���noZl���,�և䤑7J����5վq�\�=p�]S�TQ��=�.���|Җ�h&��V��b��Y��A(Q2j5�
]O�$B�%�JR���e2���v)��l6���C���(��P��׶���M�nBwX�K�y�4+�"	�m�������r�q����R�G��I���Rs�窣��"u�弦 x��w]t�nJ�>���p�I�Ll�!F�/z`6 W'��:?I�	�p�\h6�8??���	�Ţ�R#�^�3��|nV�!�3�.��j��K\�������8������r)W�f����cU���m���?��Ɔ*B����N�T���J���q�+�����[��P��,9(�uE��>�K�G��I� �V�A	(�N���9����r����8>>ƫW��C��}mF$m�gŞY��Ά)�iY��<���&�7���d�P2:U*��/A���'�|�>� ~����Sz� [�t a2�l6U˦P((���J2$�����e�d �����a�d��
�lm�zv�\���Jg���Oi���� 8;;�˗/���K���*	�.�}�9���v�[;�K�Ԍ���ꐝe;:��5�0���^O+����
Y��|�:�=ܽ^�%gv<Rh�L�9dk^Z��+�,羡��g"6�����'&V���ԑ��@�6+9]�A&>��Rw��E�Z���	��׿�Y$QH��"�z&�I8gQb���_6Eᦨ�"�<7=���v���� �s�8J
�aG9�Ȅ��.Y����>�*�d�������&�7�TR�d׃3�KI7��K& N�sJ��	Շ��<��2 (��v���JN�s��
̐1��=J�f��7�?�(h���ܳ�Eϓ"L�}>==E��A�RQ�iuuUI~��u��eGB�LP��_��U�����t)�����r��ݗ K0Ty���k4�.�U8���`0��_]]���b����� �J)9<�ߏ�`�r��r���g�m�:VC�z�ភ�؝�7C�A�2i ϑ�>e5&�	*�
����FG.RN�%��v��,)LDyhw:�Z 'Z�>d�D�2������
�*ˋm
rQ��D�Q%�
�TK<��䴼|�''' �p8��f.@��`砳3�5/i�ZGR��|��,��E[bVT	��I�b�`�Z���;�����P�=&�V���d���ӌ�&6��k�	 �!�~����F�� P�/@YD�I �%�<����$������akk�P�b�^����
���>�Ѩ\[$�ZM�m��/�>a�^�(�e���-�/�,R��&9�:�됚޴�&�T7Z�	��w�p`4���c��:�V�#R�tKZ�DxYt�!2�}�?��1���>���>j՚ⳓ[?�P,qzz��[�/��ˁ�Y�b,b�����.�o�x�v�v��iF�Гr"�Ըm6�8==U�#>T�g��d�sD�x��|J�Q�c
�ʇ2_a�"�'o�k&���I
�A�a��pLY��!<��lll`{{[���t�_����>��.|>�����G̙�恬r���|d�n�vм�B��	.QM&z�/���h6�x��5��,>|��?����j�*�V���p�^�+Y�N�&ɛ�j�I���L:)��.&D� PB�r e�&�� �~?VWW����4�X�Z��������888�h4����J�9���@��������2d��!j�ا'�2i�P@��E�TF�ۇ�w��sm������zLj��uu�K�N$�\*)GC�1���ɧ|fh�����Ƙ�M.�T[�f�v��/�����u��aD�Q%���җ]����ޏ��m����#�"ʋK�A�^�{�찖�"�G�Jv%f%&��#E�&�1��u��L�������~�4(3Jp��=���(@L��2D�,)�^OM���i�V$�4�J�h
z�kũ�s�ܦH��-�%Eiw�Y�Q�{xv�!B���T.�Q�V�����(=u&�~��V�v[�dB�z#�2�Y��b3���\Lb��ʁ�IhI/���Ut��E"����.�����������X,NR��b�E��\t�̋���n3�kh�,W+TN"�|��x\q� �@>�WH��e\4�����r���V�^WUV+r����u8�.QX&��>Q6+Ia���,�MG���~�H/��l�l�\�\�JE%�~�_����̻�v�y��Mօ&2�Z-P����a#+�Uk\f�~��<<���'��pX&��'%�x�I~��r@4A�H���c4)�Y;R�k�d�\�\�&��N�����W_�믿F��P\r���X{.�p{[����N,I��}�{}���I�'�򾸜.Eâ��乁�t'��%�A�>-er�ح+/��J�Oy�4�r�L�YR&�L92Au8�K_,������p8�Áb����(��痔�[4F�]��b�Hō�$ʷ)(�b���ޛ��u\��;���<��Q�LY�lyl7�{aC��C��w���. H����v��nMQ�X��X9��P\�}�"����")�-��H�2ω���k���,����b�B�����H0��\���ₑ�������
�B4_�i4��r��X�\�m� �)��B����+t�K!�A)������`0(�#�Rs��.�.4D�
��e���i�B�cѴ�m""*
�r [�j�諯������ަ����ۣ���T*�}��lR�٤N�#bU�h��(n2.>��|>��h(~.OЁ��o���-6�ь�j0ϧ��"�ɓ'���O�nW�ɥR��Hx7�cyXa��k����S�w�e�d���b�Q�Ë ��*)�{JF"�F��jU�b�if>��?7������ϱ�?��`��:�����6/ϳ�-\ ��hD�ŜӅ`uq���c:=9�/��}���tzz*&��Z���,ߔ�uz<{�{�I~[%����,�<ԈY
��y����\��9�I��|F�EH�[xf��d�׸.mbn'�gQ�"��u�<�a5�(BwqqA�V�R���y1||||L�?���#��Rf�oJs��/~�m`�A�ق`n-ƃ!�!FׯV�	ǣJ�B<�۷o_���1J$� �,Hdp��n�+ӹ�$(�8��&�>�l��
v��A��v��������b�CLD�f��#9��V⨳ٔ�������@t����^Ǜ�TL��A4P�{{{��d�P(��|O��]n��a/h!����f��:g��L&��v)��8���O/�W/������={���V�	}1g ��Z-�.M�M�kWy=~�����Ъ�����z/�� ȟL&t~~.�a)`K��0E��Cf_niq�R�uz�z˞�h�r� H��x�JrR�K�    IDAT�kc��y��"�^`��|>���v��>}J�?�^�'t�h݂}��7���$X�b~߄�aY>��S�~�d8_�(�x������a���H�z��xvU����������%�l	{Z�h�7�t:bh(�(ԯ�����������0i_�]	X��9����kh3���yiq����>�����D���F�z���m:>>���=*�˔������D8�]n��u� �|ݢ����j�?7�t?�11�N] ���ʊ��j���)S��R3�8!���R\^����!yk�k3����3���@�t:)�C����"��*]\\Н;w�X,�ԐL&#d �nWx�A�X,Ā�<�����k{���u���r�=�56�Ʉ��*�z=������}:<<�:3H0H�Ϡ���hL��e'�u��2�[�	�96�#������L+tVp���?�zI&�Bn��\��!�/'ZJ��u�	������F#���z�N �s0�ԁ�0����x<���1�� �kQ�>������DgY���@7�����ʽ0���G����		ޭ��8���xU!&\W������I5�*_k�&s�@����r0�N�㲝,
�D��jѓ'O�o�
��e^�[�y�
��}ߴC�M���W3uy�[�YuC���)>����žW��P�����U*�|d�� ̤��	Gy��:���b���DD",��t:�^�G�~�z�5[M�+F`� ��d2����[�nC���yqU�j{@���tSr8��;Ee-k&�va�Z�...��)�.CeLy��8�x-��(�hUn���F�q�VM&��r�
�p�}�h4Ć��_ ��r	��y{N�)�)4����O+��e3x/�n*۴��֫������k���c�
��ݥD"!,���'3J�~��}�bmr{lV0�F���R�����x/��%g�Ѳ�k��<�
0t �g��k�B��V������z�����jö����>t��e$
���e���/�����B�3�E�c��5"�<�f�4ǥ��(Hn?Հ�N��C�h�����_� ��n����rH�R
��������tpp@Dt��݋x����8|x=g���T�ve=��s��y��,?�)8^�X���]\\��8tzz*��!��١��-!O��c��ċ0n�s�k�E�� ��_< �x�:���x�j5����������qUŠm������\[���kR�
��je�*�5gggT��(�J��|>O�lVhy�1>��X�[- ���o|�D���xODD�lV0{�PH�!������ժ5��{"��P(���|X`b��%?vD��N���\	t�4��]���׆̄��l���4a|��[���� k4�	�gD4˕>��]�6V1�K6��~�Ї�C�m������\g�?�p8�"�HǓ�` d��qF��M�ZS��4�n��[�I�:խ_�ߙ�����t�*�9Ӿ����ƞ�T��� y�~���6��mWҖ���J����w�p����ܥJH��&<��AU���kc�R9��J��!�I�8w�����￧gϞQ�^��ks~��R��vm�(����y����ٕYw�;/�x,2%���E�r�|>O�LF��xo�N�w+�&������
��*���4���Q�բN�#���g�|��v��7n�����W��*S�:+2/ �}jqay�6�`��*	�м���Qw��}0�P8t�ւ(�����[9ABqyy)*"��!B�=��]��8��x��&�	kXfc2���*�i�!�c���U?����F�D$4�D$t�[[[���n�"9I�ӱ\�hT8/A(�	7x���[�q=��y�5�`��=��@la`W��PN��r�P~m������e5c*�a�L�����9DxI�l�q�a{���sr�t4�P��̇���N�Y��f|� C�y� ޫ�od/_�^$�p�͟Kq��k� T������j��Z-!O��[�h�C�FV�_����bz���a�3d� �[>4�;j�|��}�F���+��`�y'���r�J����b�82X�6�M�_8`��,V��y��F�_�mA�Sd��A���K�.W�ޅă���0�� �Ft||L����,L+l�x�� _V�ZB��p8�^�'�R��rq7�z�Yc��E�j�Đ�0�_��U�<�D��m->��e]g+L���� C��~aKw��}�u�X��XL�N����왩�� cz�!
׊)���W�*6\�*W�N�� �CaJ�BO��t������І��
/vu��`6zS�.�	hڰS� ���:��-`������� ���8E�
��Dawo���\v�A'�,�*&W�v�;������\��Ð4 t�`^qv��}W&>����c������<�)u?R�fU��x��%�31�6R:"��;�$�q�̻��4j4B�]�[s�Db��������M��� � .
��*��'��ok�5w�����pS �DMˋ��p������PP�����a�����Q���$��
Y 6!���	�'�P��~�E�#�"�RB0�
��CiH_�BB{Y�׭��xIl+U;�.�Z�
�U�[��ߐ��1&g����}�T*.�-lPܧ��&��ryͲ��������A7� ƕ%��ŕ]g���3gkg�����碝�8�F��b���|~ӿT@b]vv~�9]GL5����%{i7u���Ml�w<`r���bk�'���ҁ�1��oy0����"_8x�����]��p8L�X�R�M�S���t���|�-+!�k6�tttDGGGT�V�^�����~	?3�H����>��.�M�2K/��\B�{̓��� �V��b�A�a�QxF0�$[2r��yNj���2.eW�n�M����Su��k�(܄E�pk�*�����j��?ҸN��'lj�85W+5��P:�vU\�x\�^ְ�z=�t:��Ǣ(��9N$B{��`����y�M���2���xlz��e&�m�+/vQ����Y��Z�&l���d2���5�3>�uk�=/�/[�D$6+l\r�cP���f3ZL�$����ۿ��P',d�!Ϙ��^���i�̶�����h�y=�?����`z:����Xu��ɐ�-�{`�Ǉ��gr} &>�_#����� �BX��|������ �8�8�YR"�2���p8L,�.�����^����)Q�^� ���αƯ'�.R�Mq3��/��aٽdY���N�����`��؆������T�up���F4�H��s1E������ę$6��vS��&����I{��Z~^�=݃�7j��е-�y����8.;$~�0��&^Q�x}Y�+����-4��c��zhn�$��Y� e��uZU��o%m��ނ���j�.[M{���lv�T�r �����P(D�^���Ё�W.��q�v�Z�8�)@D���)��� ��*�$/h����FD.=y���1�j����p� �kF�:��j�Џa�D.&�6�����*{d;�m�3��2���$���CV���~���8ח��,�`0��� ���Mg����.��x��:*�𕔂ܡ��:�#��Ad@���1���` �!�Z�NOO��l�����d5?-b��8\vM�H�e����qX蚊	��Ŏ��ɓH�Z�Cp��=B��k���D(�H��P��b���cN���d���+N٦���U���4W5��c?�7�cT�y���>|��E����,�l��ߣ��/,R����d2q�t�X�K1l�:�if&�uU��u�e7d�{ٜ�M ���Kz��9���Q6����M��ؠ�x,����1��Jg�cA�d���'����]xp�D����l
k�f�JK��u���
m9�D�ɤ �O�֚p�6�eA?k|�ޛ 
�t#L$²ݴu1\^���0�]��`8�9��<7����}:�
2�?o	�����-����!·A- sV1��~�G��h4*�:�¾qqq!�nx��B��)@W��
v�+�*��v���#l�+�ϳ�p��^��ζ�
k�wW�{|�1>�&��Q�'�r�#��������y��[Ul�
�NR뚋�i:�4 `:t����e@�����v\�!����_׎�m$���z�����2��W�S��U1-�k��7��������֖�')����G��/����65�M*��T�T�\.'�ah�U�J p������Uמ;�u8��#�#aW�o0�T*E�HD�|���txxH��th4�p4tE�"�\���D�Sܪ����*���I�Y��i�0YE���؀n�3���mf5r��e	�ra�s�PP�D��0Ɛ����A.�Qi�&�>p�/�Ч�Y���r�n��tttDϞ=6M(z�>dok��Y�l"�tá�tJ�T�H/��Wwq�m����ٜe6�U^ϸ��x�����3ª���s�eܛY�ql�h/��g��(��6FvW
�@�_�٫��#�Ŝ����`�FY�šZh����JT���F�ݘ^$/�u1�
���w�No�H��Q��B"3��Z���>Rl�ͦ*�d2�ǅW��=��ZElZ|Ms����q1�ã~�}:�R�ݦ��Sz��	}��t~vN�ˁ�u ���jБ� @�ej������'��t%t�W��mq����]�@��3�*�uCl(���MgD���,�JS0�2���`0!"�6�`���i!��ȭ���>9I���ˡdt�����J=c@���<��ǧ��"��h\I��x�j�J���T���σE�oW���@&i��d��ܑ��Ѳ��Nn��*;B?� 6��.�N֠�@�KT�^C_�[������u��`E��(��5�����i�6T[FÏw�&͆�e2l���b�$�Ԧ7	�̮�m������^��6k����� ����b�á`s 4<x �Q>hx[
Eں�~��0���:M�?Z��������*���)�z�kÏ&oC�2���U ��}�u�l,�t�p��]�� X��s6����m���c�>�ͮl�/bE�W��|`��|�s6��d:q�����
��`��L&�P1�C}��Λj=�C�<���gggtxxH����j���N��mc+c�	��*̦�;!�����M~R�L��FO�{�� c�Y�e�<�!i�À�{j������~��fr�����L^��\���6F�a�<,��ʡ�]@@5UF^�� uYد���^5S�&�}���ݣ�m�'�e�;��6:99�H$B�|�vvv���ЮR�%���a�A(�V�!H�T�4�^�NNN��ӧ�������|.,�L�EU��=�)��)^��*C�~�M�E��K�iS����D/F����)�m�/�/tl�;X��� �xJs�˻��F"���l6�����>�N��Df�d*|?�K���C���tzzz%�a�0������Ƕ��(��{������鄉4}V���u�QˆT�9�8�U Ⱦ����G��Y�U�y��U3C�v`�u�Ъ ���.sC��D�^C%2x��IX�����A�ͿjۣU*/�6��7	��>^kƯ��뚩�sy
{>��V+�!��@���_��lyį,��F�n���o2��=L�w:�t:�6vD�$����n��u�u:M��X�~��@�����^��T@\�3l�����5�	�0h���
�"_WTBG @�^��J��Dk�y���@iP�lV$Fq;GH�4l���=??�j�J�ZMXI��*0U�m���u�23�*��:W͑����M�2]Y
���L�����5�Ǧ�m�)��+�������<�u޴U ��~�+��4��b\Ml��[gz]�"��x���f���V|���~���
p�LĤ͆!ol���2x(pe%6_P0����r���!�J�< ��=�aϭ����C���k�`6��l7\��"�ky�֣�lӡR�G]q�u@�X*���Ҥ{�tM��m�\5]ojw�g�[z���kZt��PD`��|m9p[����Q(�V�%t�x.WH$c(M�=���cN	�^O��� 4g���W9t�I?�E.Nt�Ҷk��	�.3ܶ.g��S��>�^{�j��[�� �pG����Z��ެU-���pl[��5[G�M�{��0oښ�un":�v��U��8ȹ5\"�Q��O�kg>~��p���a�gA���t��rkr�.Sys��ku,�M[K�
��SU�]&��u>s����uf�&�īf��쯶8�gbn�~�p8�n�K�lV0��Zή�$�u���Hu����-� z9��!6Y>��a���4�
�`F�{�:4�~u��2co,5uW���A��P����{����U��4j{ή�|\�W�&u�̛�a�cټ6[?<��֫-�'�u}�i��&֘IQ��k��=צʇ3Z���\D�
�˄�!-�]�74�"�Z-��CK�'������'�E���5-���k C��V���ψm�H�~xQ����e?�g�U1i�UV�*�@�s`�������#>d�������p5�/n��e=�x}V�����k�,��]צs���
6{��S� q��H�G��y��׶�O�YU�ï/�n��d�j�~/���$a���f3���~�X���=d6 ���[�S��I=�i�T����)H��!�W���˚�Z�˶?���,_���9�4�N��2� �/����`�ƣ�a�������'�$�����c�UC%*+ΊɀWW��ֆ��������)�g���������Wr�&Q�;�֡;e�
HZ�a���V���|�<8y��x4vIn���a�ţ�!��"� M�<1�fq�8�����4��>q��LN>��@ݜ����ܰ�&�� ��� ��2%ݿ�kNu}���MϢ�yl*�u"��&�:��֘����%�N��4��еY�~�ST����L�M�S�z,��,[p��ˀW�a�Q�S�������i�V��@�"O���_x9�_]V��
g��xjLhs&�v|���K�^������^�N�'�9�T����&0z(�8�L&]-o�� p��$"hk��9�������MX���= L{=���^=<�|4�l:3�p��Y(�p��ŢW2�f�}��~��Y7�z�u���mB�F��7U��M��*�n�M�u�{>��j�P:�~��}��+6���#������Q��J�^9��]�~Ӯl^��r���� ��:6�ϗ��U�����قT��K����L������^�L���Q �ܚ\&��˷Zr9x [̙O�@�
����V+�!��n�4*�4QD�3����h?������m*�J���;�,�8��	���DD���}W�י5(�8K�ϋ��|�ۃ����,��&�ɵ�\��k:�Rh���եR�M���ÆI��{�`	ݙ�LG��ݏ���:/^�9�.=��a�E�a&?^ܶ^�~3�D�(%���*�U���ۤ��I`�JY�'���u��X�r��2����lc�{�m׀I��'���쉊���2[P�G���YU ��	�����O�֍�&�6��r��㞩ܖ*�H���x�D"�J��Wj4�R�1���P�R���ʯ5��`�����p��L��"4 :j b�g�0���zo�C��P\�����dO����9�V���]�u��[g�UA��V�f�V�&b��{n�m�D�����/�FȘ\t,���k�K���9�c����^�*�&���,��Y��UmV�U�|��@������h^���d?ĲE��&�Ɩ�5D���CR��`m��\�a��p(��d���_U+e�ƪC�3S���kS�����x<�(�_8@�R��R)�/*�ܡP�� ���}"��t:M���_.�-��tJ���b
V�	    IDAT�k;q���>5�M��ͦ-�FbZ���<t�]���t%{q]�J^"į���i�!/��zW.�F<�'���#�6�P2���+�Ce�?�
$�3�l�1���A:^��K�%��C��t��}�u$������yS6�6��u���}pm3�Wa8M���p�W��-�k���ˏ7�����P>�b���q�Xf���N����ڬ_[�� ��V<�VŸ(�t��拗J��")	L��2ϩ�~��w�C�V�z&M�%�Ͽ�N��X,F�D�r��Er��%	*�J�����ɤ�,�A��I���.�����`SaŖN�]C}\�� ]_�U4�M��r;*����u:;;���j�Z(��c�o�j`jU�V�G��Q���l��X���`�/�,��:�9@j�u�^��_g�u���uN�x$늑7�-�����g���	�_?ii�:7����[��!/>���K�m;�mi�J��L�[Vki���:�l[I�::���n��iJZŬ覎�~�Φ���m�[�0�Zy:ߴVL�_�F�\�ρi�\������T,�P(P*��6��S&� ��2�ȭ���1@�l��5��Z�=�ˡ5 ��<M�\ΥمW���f������NOOi��V�	�/�p�9��ۉ� l����q_Yx�b�l,�P���\Ȓ�e ������ڛ��ˮz���5}�U�X�����j���n�O�ʫb����o�^���U��B��YJ/FX��u ��,���.�����#�g�yp��[?�겺�U��e�F�k%k�W�B�������-�Ζ�
�rp˭�d�ƃ��<��Lf���W$�l6K�r�<x@�oߦr�L�\���,��i�~  ō���`e6m>�M,������i!A0�L&�x{�d"I�hL0ʓ���~�ܝ��}�6���ѳg�����tttDB �Ǔ�V9@m:��?׼egW�М�U=:�+�Eֵ?��^��&���2L�@b�\�v<����t*��g���l|�_������e������gd6y~�zm��hX`t�
p-��Y��P���jj���bm*�e �Cp�A�2�V-�L;�
�b/�el�U�lsdk��� �ޡ�Aw)�@��� x{V~^l\3��RL񼦈O�ߛlS������tJ�p�ǡ\.G�R�vwwiww��ݻG�����f)�Ɉ�2�J"r�;�߼��]8+ʋk��D".��g��Ž�vX�G.��h�`g2�T*����Ǐ��/������z4��f�q"�������{��6IX��X���6M�R�,��b6�	=9������_����Y�e�v������Z�b��H��4i��s���u�s�3�� ���(ѝ3��Mx��m��U�t׃���"P�{N¶��k��Z~]LU�<�b�F���x�������m����:�l��v �¼�I&�P]�<���c'��k'w�O�&��<���l��M�Cg�
G�!�M��˖K0h�8U�
�mmm���mooӭ[�hssS�kq�~��?4�\R���8�8�[pn�C}�i��
88���8C�����_|v�7�@�:T*�T*����q*�tqqA�v[����Bk����h�y_]����k1<6��`����{F���]�l�T�˅�N'�"��>���ٸ��S�G�=��x�|S�	+����q���a�����+��ᅅ���-ՁV�u�lqaK�鼖m�M�3���yU_~�U��M;ۏ��vY���d�"hm��Ѹ	���6��} l,���+���^���olu�U������`�B��K��@ �.햟�l?��o����@+�˴��K;;;���CT*��T*Q:�`v6�Q��w ���D�l�\!&
� a�a`_///��g�0��s
&�M��31v|��� �����F)��ѭ[����H�]\\�����uj�Z.�/g��l��~���@)��@��B�r�E"����W%�Yf�֥Wڐ3�A?�Md�Ҥ�d;�tx�z� n��ZU��z��B��ד���^ƣy��C��u>�U	��Č�e6��\ �,?��˂�uO!.�@�&�m}������e0]ܟΥ@��YvS�	��b/tŋWKO��pI�p�V� {	�(�y�Z�Փm��O�c�LCw��\,�{6��P>��t:M��ݣ������.mllP:����S�� �� ��
�� ����s0����{��l6�D"A�b���"��iqu�k�y'��5ץ�i*�Jt�����T�������������NOO�����n�J��+�z/���h���ָp�Y������P�8��E��<zI�T邪=��~{1�6��8d)��S����� ��=���xu	m�"p�#�l>��sۏ�FNN[Ǚd���-�=������j��ׂ��/����$ �豩�l�ӄ�MK�V�c�{U��׀��a�	�lî~C����c0��h���怆�WUl�Z|r�2g�T-)<�ʁ>�|(�x<N�b����iss�677x����7�1 &�L�x� ����0���K�Y�� @;������h$>���;@*������ؠB�@���
�7�@p�Uf� S�^Ȱ��?g<S��L�����������4i8^KF��*ς�����3p�A=�^\GX���b8��H���uTI����:��D��%Nl^�/٤b_����\c-�)B���mX&��dkiӑ\�m]g��0���M�0�h��kk���W��A�Z<o�ӂF��^Wڗ����:2=6��*ޖ���,lk��u��޷n��F�a; �b,y+�Є�!��.�$�Z�.[еob�Ү�{t�� �����d���޾}��ݻ'��|^hM�Ѩ��/�8&�I]���9є^z͎G4���jQ�Z�n�+�-O{+��ܦ���d2I�B�
��E�f�"\"���8�ߗ�e���nv�؍D"bM���x,� c�e21����E�nݢb�H�@���&��u���B��]%��XU\�2Y 0���|�5�2�3����|�`P �@  �����bj����'K��"�_S+��m�ޫb���Ժ�{^ݰu؆��A�Pغ�xS�_?~���vU�g;$���y��K�u/����g�-�U&bob���R���>�/j��Z�6ZU/���]U���7��t��K��z�`� ���@�d
��	b�z�����s	�X�ʯT*���I���Mw�ܡ۷oS�T޵��?x�*���|.�e�dۭ^�'����9���`k�ݮ ��>��-nE�Q���@6�L�����; }$�X4F�hĕĆD�`0(ޓ���r4�t:-  B/b��j5�V���-Ui���n�/ �~�O���� w^��b�������� ���{�\��L� � ,��A.�.����
wPI%�I��%Ll����*ߴM�,���������a��չ�J.lH(ӳ�e���}pM~Z~�lZ�^���ŏ͗�`�M���ņ/��XG����g��`��UQa�q�$)&�[Ujj	.4�u���n�x���Y�+�7��i<��U���:�4�����*^��1m�6 XB����)��q��ݥ��z��޽+�vvv�P(P<�V|~0�r\1� �z�N���T��\�
r��`@�n���>��}�<��
�� 4 d(r���kj2�P�ۥ^��Z��Ʈ�n$z%�����\. �L&E���8���I��۔�����.6��t:�1�J�V~�P������tqqA������3:>>��$��LJ��i�uF"��`��z���=o���L����W���rN��q>t&K}l�,�sAe�hh[UC�Jg��̱���#:�/y&�)Y��ǽ��?k��������_��g�O|���)WxY�?��3I!L���4L2 >�#kܼ�E/�U�et�]B������+7B��8����ʆ�*FO��L~��£me?Rhҹ��SlbYu��2�r�:
���t6��t6uy�rk% 0U�]�[���dm��Uϯ���8��a,�� ݻw�~��_ӻ�Kw�ޥ\.' w& �����w�@hC�Ѡ��#z��������F#���B�ˇ�.//�&�?_p@;̵��7�s��L昷��L�6�Q2qp3��R)�}�6���[�� �N�B:�����:�Co������d2�z�NO�>�l6K������i8�b��l�ugTU���=G�]=�.�6>�)wmp�Qp��s��F�Q׿3%��.������*�ȟO�@U�1�V�M؋W�L�o�k����^��Ư��֥I��6�^Q/��d]jK��W�F�4��`��$a���2�v�/h��L��>��U7�o�\�v�fq���-�y�	��7|nˡ��d6o�ʚOk#�~����o�zġ&ݽѥ��2%�(�e��v���s�?_{\c��;�r��֢Zd�G~O��P	�tww�<x@?��O�'?�	mnnR"�� ��#���b1rGH �OOO�ɓ'�����_M���Кr?\�g�S 3^ ��#�^��į����� Ϻ�
Y��}��aoo���Ç����s��E�(c�p���d2l.�r�L�L�b��`��<y"�-�fP��_5�����9]^^R�ӡ�pxu-�h��V�D�5sY�L&.�5o����W	nm��<��,�2�uP�zI
�u�Y׵�9 ��㶲	�$?�'����gx�bi�����˄J��A���òh�v��͊W���M�����/���ĵ��p��z�Ϲ���f,���;$h!�� BK^f~8h��]���˭6h]�U�@�ژ���%
`�x��o��22�Hn�� ^��f3j4�h4(�҃��ޣ_���������(�L�"q��r�4��&�N�...�X�'O��������������ȩd�gĵ�L��@�I���"�ܫ�dB���&���w:j4�l6iggG蔓�$9�+��0�W�p�H$B�X,(�LR6��P(DGGGT�ը�l^��/RŰ�5����=h>���)�4�8��C������<�������O�.�k�������i<��JәebuU@Ֆ��J�2�s�fK@�ޫe�l�~�`���&,��b@Q��ޤ�-S[z]hM ��%�6)~�ӛ���#o�8�98�-O 8k(3�6�:�����0
�B�e�#V��Eu4�����`~���.T\.�`^�p� \�OfIuL��������9���mO��<勇#�b�������/�K��OJ�����fi1_\9�pE@�F�\_�j������o��/����c����@ �����aGl�*�ÿ����_\�^�G_��p8>>���=��ަr�,�.>s(�q ˰���T*	�:�)�Ɉ��+9�i}<�M7W0��\����fn�%ƞ B9Xx�90��>�&�������2'{��]�w��L��mj��3�G�$��	�͖���c]����K/ܡz����ꀫM;Նa~��� �r�'��?�M�q�p�&P	ɂ��[;���B�p&���`?�S*��s0�O��n�XM�X8]���:DAR �9���hq�=����7rx��*k��V�8e6i` G��Ѐ���?�_�����{����9�C��T��r�6l�B��C�V�tvvFT��i0�a���c:==�k ŸFx=�C��Vцy��q�k�3�|Mp���hD�n�?~L���S*��T(�Ν;�q0�x���P\b��b1��ަ����"@�\.��_��ƞ�=ĴV��)}�ы"f6Cp�D����C�a���$���3cӮ�ρutuV�Q�����_y���灓(^�]�,K�T��jp҅�l�l�
��=]'�U��u8R��,�=Xw���[κ;�{#|pבfacբ��z������R	���{Ζȿ�=	�MT���h��\'�u��@	���d�<����Hr�n<�d"I�hD�r�Z���΄	=��S�5�?l� ��&�D\�Q 0N�O�a���g�Vt�ϭ� ��Z�N�b�+
�/~����~F>�w�}�vww)�H��+���>��?�������ѳg���ӧtrrB��z�u:�'	Q�9�Z�;^mJ��=]��+�E��k�ۗǡT*%4�gggt~~.����ݽ{��}�]z����޽{����˓�d7Q.���B�NOO�����?N����h4h6�Q,�c��g�� �:�Lh4����]�L'��(�JQ�P�?t���PЩ@�,�ᅾ�A��5������c����Wa��?�1ɀ���n��[%��:/V�{){g�û[�aŏ�̪�ԖU^s�e��"Nn�a}U���s������z��o,[=�̨3���RU�D�� 2���+jn����AѲM&��тu��L� lP��h�k�-L|��!�^�N�B�����ϑ��U�*P�N�[FW�˃X������T��׌�T뺭��5��ǰS>����-���G�կ~E[[[���A�DBEA:�|�z�N��������������?NGGGz�p8,�B��+)+���L�I�h���Z�i��H`���&�	U�U����Z�F�V�:�����T,��./Jy�'��m�`0���c��],�h4h8�U��8~���x$����1ͦ3�D"�N�]��^�Jf��Q�o�:�/@�eh��w�0�żW���}(FP�rj�{~��:��Y�p��5����?�l
i���z�׽u��-c�LGjյm"��������[yӒYZ�����p�:�js�c:yۍ3ur���&�@x�h4*�����1m��X��u:��._S� SY��A���6t2����-�f���h4ġ�6�
ܙ�y�e�絸.Pl�/�pC�I2\���g�Y)~ �zy����zmJ*F�O��B!�f����C��o~C���o����"� �]�arp���j��o���?�����z��	�z=���I i|}pv�	/F�&E翬�'t�W�\��~x/1���~�OGGGB����?�1�r9Q B�*GZ�:�C�r�B�������&�o��ɯ5�'~��m<�t6�h$�j�r����l�xSg�m��kF�${�1�^?K�oe]��oT�@Sj��� �<�$�H�3�'�qF2$<�r���vr8��I"�����}�>�~�N�17��l��u��=o��>�k��յ���]�d	�.�e>�W���m��f�[6�pUS�<�Uզ��@�6��Q�\�d2y��{� �HL\�V �g�-S�����ͫ�����2x`����>��#�*�����U�Uh��K,�T�~c���9��g��s
.�C1�HD�SQ �~p����>�3�L�u����SYA��>��8��i��ؠw�y��{�=z��mmmQ:�iTr�-�`0(����;���g���':88�'��V�i:mQ���:�!k3�dr>��Q�J�֊r��d��{���}Z,txx(�E���y:��\.�*�d�">{8�l6K��ߧx<N;;;���O��Ǵ��O�fS{�s�=�[����K�.iJ2�����b1�,���O<��ž����:_j�t���PͲ�������bs�x�;�
O�,�Wv2��v��	�k0��P6��Լ�D�"v�DBt񸿱���^��	_� ��-u:Q�#�{�l�����ᦘ�䣩h�%����Mu4mp�_����kzm�y��bيۏ�o �.h�����ep�D��q�A�(����$e2���T*��q�k��y<��q��D"�F�DrU��I&���� ���%R��ͦ0��>����!E"�FT*�(�HP>����lR����<謗��f�2��k��`TL�|1����ωF�עM����O���躶��Y���UE��|mB�p��=z뭷�Ν;���o�� �� ���������W_�_��W����:<<k�}Be���ip�Ip�ʚX������/Xe�<���W؅<z�����B��    IDATr�
��ۣ��~����D�/����+
Q�R�t:M[[[���C��������Ϸ������2�
J�Rb����e[r���TKe��ۗM�Q���TH/���=�K��cVU:y�vd,���k���A���XL$�%	*���[A-x=�W�:`��d@���]rHt��!&`�A ��z=j��b�r2�P�բz�N�j��������Ъ8i�A����M�[�9b�^X5L�����j+�*�k�y�׆�dJŚ��{�M%�N�����wG�ț3?8���X,h2���l���Y�AJ�R���N��N�]������<u:ᒀ��.؝X,&$	h;'�I��١\.'��=`�dM�ix�o��w����0������4���{�C3P\�e�k}/�A��?T�����r9�я~D��կ��ޣ��*���dD[\fD�4�t:�f�I�|��˿�}�����O�ZMX2�ɯ7��*P`ړt��Oڴ1�����\y�����\�OD��v���\tWǡ��G�C�_�!� hF�9�������y�F���W_�n���^�^��4�N�p$;M��`Mq��zƴL��:��^�=��5�yY���"�&qpϋ�x<.d+(*p���(�p� R�֦�irG ܭ�-*��s�9�L/�v�^��!���z�{"��Ù��d��P(�nQ�ץF�A�z���:�[m�^
�i�O˝S+jk3j����L'�M�BS9;���ի�	ә6�	>���������5�#%[�p�V
�J�P�B� 4��w��T�A)@׌���;8p_]�O0&�a���'�HP6�W�բn�+�.��^H��ަ��J�Ӯf���X���N7�����k3� �b�p7���Uz4Θ��ɲ&N�nۦ�ȀNf
���`0�`0Hw�ޥ_��������z�-liA����M?��^����!=~������Q�^!��<�O�w�!T�Arq�PDٲ* o:ظ��k�U�j}��x��mڊ�"moo�g�����z�z�����Ľ������N�EY�,���f^ǜ���P�],Y��!��^y�A�D���=��T�VT�^?Ŏ���Ս�����`n0�l6K�|^���!���t:M�l�r�e2WᄽQ����*<�9���::}\�/�9 ��~N �<��/BDb���q*KT*����R�բF�A����v��� "��r����X6tAW��eUu�Y~���0�ߙ$�!3]G܊�5Q���o◗f�OK�4@«v�G�_���� "��E+(��P�\�b�H�|���,9�#tvظp��A.,h~�ʭ;<ȼ��Z<U�o���,,��\.G�^���!��}j���n�EB�y�v[ǥ�i��ۣB���[4a!d����C���2E�tT��g��d�]�\�}�Wi"�@�{�ʑ����m;]�6x=��P�vvv���ߧ����޽K�|^h�p������C��f�J���ݻ���%'�l h�6���7spu���p�R�P@`ӭ�1���|ve#P(�P0���ȶK*]%��y-
����}��pF��	R'�����-a�pϐ-����ކ5 �֜IG��dpmv*�zq��"ї��*��)���g.��z|�˶d�f#�ӹ{�<��F��i����`Y���x��ܤ|>O�t�R�������w.���q�9���
�}�����:�?�^�el(� �����f�P(P�ݦV�E�Z�NNN��lR�V��A-�Gۜ)�t�W��7A$r6U%[��/��dp�)!�!|y�6~��i3��N��ê�؄��VQ,�l6K�b�
�U*��r��36|`L^x2#�7�\��7p�67���^\�R�f$���v�M��U��l6����~�O���b3��ؠx<.@���h�a��s�%�,[�_�����`@�p?t �3��p/�b�4�Mj6�b���l6ր�h'j�-N.� 8	�B���G|��������S6�6a��Jg�l�b1��ݥh4J>������`�9�[���'p�f��๐�QT���B�:�D"����Yg-K���O�ˮ� �m�ǡb�(�Oe|���<y��Y�E>��|Ȳ�Uh��p�7fU��V�Ѩ `�H�≸����5u{�u牋�<@1���ּ�I�� �HZ�.�܉�]�d2I�R��٬ �(*�S�ݡL&C�R�J�mllP6�u���������K�z#��/� � �`��%�:/(tv�b�Ţ1J&������jQ*��ڶ�q�A�u`0G���*@sY�zկ�*要���]��m�?,������6�ѨH�A�P(P:�	Chp��'�e��?��P�Ѹ�����&���s�Ψ���@  &���,��u��jB��j���l���>�r9*�J���hkkKT�pW�ǆ�XF6cS�z�8WL/?,y�����=��şCG��f�L w4Q��l9��*�+��k��K��cr����藿�%��?�=|�Px��@�=O^`Ɍj0�R�D�|�~��]���~�p ���%].��8���d2���fɀSfKe��J����IPT �j\?n��#w���Vn���J���,i���=-�t��-�����M@;��Cv��Ů �������D��q�.{��Z����ˁ>��~�O�ˁ���`^	���m��u��Pqם`0H�B�677i{{���$�j5�v�bŽ�������H��>�CC��:�/��}0�=c�TJȂp����Wk�K�f�u�]�!�d����J��{C4�b�H�����%U*:99��^ݟ�)��pY����e$|6r�!���*��7��bS��R:��)�Ru�Qi����ף��sa�@�N��@?İ���p[)0��p��?X�Ӭ�z�������_�d�CU��bl�N��ݮ���T\�%>8�ńO"�[<ӳ�pX�'Q�R|���*ݷ�&�k���IW�x|������r��В�|>'�q(�����&��iZ,BC6����P�Ѡ~�/� ��,|�Q�v�!H�PY�P�w�y�~���������y� �h����:]�G��F�@���q8�`�4-���lz����8�՜��� 7R0t%��SD,/�������P�[�.�2���!7���%ޟ"�@^3\z �"�C Bۂ���t:M�������5Z��\ W�i�Cd���Ǻ��ϸ�5�U ^������s���ZP�^ ��=�z��htu/CWS��HX� p�Ys�s�Y4�2��ܺu��ݻG�RIt�`��	k�b�HBʐL&����N�y�r�zq��R)rGs�0�A� \.��LDIf7�����3�n�E���J���<A#�}~]���%έ�޾*��$�2������n����&6�4��z����M��k���o*W���P��i��X����K���B���@ဎS��N��J�D+2�Ɉ������D0��"���w��}T���f��f�ٌ������l6�V�E�Vk�����|>����Q�ۥF�A�N�Z�,6"|f�qh�E"1�](h{{�����ٳgT�V��n�����+��t��}
�trr�b��[u��2�Ľ�ёu��G������xL�h̥����y[,֐�������$�s�Z�j��B�`0� ��U㌣�WT*���~F������wߥb�xdGC�>qp�&aU��\��C�/��d2����D#F�T��t���%Pց1-��"���\k��<t3�^^�<�#X%��Ê*�/��@)��{I��ٽ�=���W_}E���4���	<s��H ,����B�w6��Q�㹑3�g^�Q�E��8�x�H$r���Qf�����\�k�Hɮ':?x�T�o�W&ߺu�vww���q��)e2q/K��E��r�b�A'g�qV� +@���'�ɸ�!��u��|��d2�G"������a�3�0>�=�v�ٌ��>�Z-�w�xo�N��T*�����SA�Ȯ2:|?r7/ɨl��������*��DB�D ��F�J+����~�JU7��}ڀS�"���Ѵ8tz^Lx����䠥�}�6U*QU�͑OCc���[`ɔN��X,R$yDDg��`2��B�����#�:��GD���}����l8�~2��a6�}Ƶ��S��u�'�'
���V�`a���#��� l������3.�$�溶���jHI���$������T\���˫�)�g��~>
$�J�l�x �X{�tZ �R�$�N�#<!q��5�I>��8ݿ�>��z��!U*�D"��]����?s*�
`CK'k��#�^�>��cT��.=�t(�t�2p�EUۤR�ڿ:p�����Q�0WH�~>����rvv&�4X� ��*w:Qp�U �`
��M��Ǻ��&�>�K3x|�ʏ\r�� �kqQ4bp	����Xӽ�!�d]7f8J�U*�h��766�^�����&��e��'<�;
/��W ��T�����d�q*�
f2�P<��ř������g�����x<Y,M��///)�S&��{�x�N�����n�]z�J�B�TJ�����T�ו�^`���n�$뀶���n�4u:m�0�в�������o�Bl".�ы� �?#��㠇����X,FNҡ�sQ���M�L�%C���c\���q*�Jh�>���;�L�ӡx<�����}��#"ztqq��x<�(��Ǚ�B��F�ч�<� �����7'<��0�E^� �8�F
�Btrr"Z�|��9��Xt0o�q ���9�0kŽk�0�� h8 �&�P�Sud0
�0(��8����B�^��ܕ����";;;�����<x@�B���ͦט3�!M��#D�J��V�a�%���p�bOTIV���2�dI&�i+��u6 :�ty��K>�;���i2������O~B�ᐚͦ�+`��Y>.�8����)�Zɸ��ݫx<.�> \n5��`������׫|�}�x�U�v:Qh�b1� 0"��}�I3��忋F����R�P�R�R�D�d�u�lnnQ�ף�bA�R����<\n2�
�eX:�r9���f��ǙL&�L&C�ht%@+mnn
B�V�}6�L>�F��@ 0/
-�!��e��d?ܦс@����U�3��p�+�b���xhݳk���)i��yS�AG:�zM��tR0Eߔ��F"a�{�B�.4� �����4=�����ܠr�,L������hա:�T*�����B�O"�ȧo���#z�_�J�� �j��:��������Ƈ�v��5:??�<�����o�,�ݙ����t�Am���ёبd;!����3{`���=dCg�5� �8�yZh��ns=�>�hf��b���1�5�w%t��D��5�Mj4����1� ��t��߿O��ݹsG�y�[���D"��/(��[�¥��T�'2C�۾�si����(���]�����(e�U����������}�hZؙ>����ǔL&�P(P(�^�G���4�D�/y���]C[��U7�\^�@S��)O�e�R���H�b���5!{PI0d�<�k�eYf"��^�r�?�]�� �x�Q��IY&�ͦ���R�����pM@���\.�9z��|�B��M�X�T�\.r'
��X*�>gO�Tr�=��Ï"��$|4�?DqzzJ�nו�H$\�:��� m>��P8$�g��� �-�
����:nb��&�[����EA��J� `��]U�ab)t��m�����+����6�ϓ�8�Y�	�=���8
�<J$g2�H4�xkk��!_�t���?�F%���h4�������ϟ?�j���W�`�v��X,(�N]�?ڙhŃ��f�\N �ئ���1� š���haB�\l���.�@������r|-׾�5��)[]^^��A`& i��O6��~�O�z�NNN����NOO�Kg��񸈁�d2�؝'�	=,;����-W��D<{�D5�o���`���-f���xU�� ��`@ `��~�\hq�k`����3Ր�I� N���v��@�R��Ɂ �������J�hgg��z뭫���C�Ǘ�X��aQ�!�s��*j�_p8D�I�Ζw���'T>Ѳ���Vt�^>rk?<�D�%��z�x<�b�q>�{�Wܻ�M
��m�PZT�0� K�٬�!�+���L&i{{�vww)�H<"�����#�B������|>�*p�E����}vyy��b���ŏ��������ĲP(D�h�(@���y�n\666 ����#��c��`�u}��X K�Y�N�M7l)��&|�T�tk:M���d���d�o��e�Y�u����>lt`.!C��ܤT*�(��}���>���~�&�۝�Wu��������?mll�����j�� a�f\Wʁ%�mYk���Ύ`m��h#q-����q�2s���q&�a �<q�k��c���=9��=�F�+o����F�ȍ�e�1�3H\b�
��;99�D"A�l6Ł���
�W����Cp��$6�W�y��r8
��l.� 	P+�o xp�=���1�]$T���R�t�d��tp^z7�a�۫��
�Z�:&�]�aQTq����M�f��J�\�x�r����	 {��p1�ngŇ�Tg���0�u�����V.,��p�2�9��x��٬�%�3��X���4�F#!gh��JI�iH[=��d�,��<��?���#��d2)�x�T*E���t��mJ&�����'�b�ӽ��7��R�z��Y4�}4��h4��Z�
��`0H�@�U�"1E�HUL$�H$�Z�R�ټ�*�+�&��^A6~^�ֹhp�y#��<����K��k�d���I#�<w͛|8`��i��@���@e6�'�T*���666>��r��о��>���ϫ������s��:�·ggg�l6���R {0D��E�}1\
�(������f3:99�F�!Rup�x1c2+��m0�\�����@��$`ox��� d���PAܭ��42"�����;e�zy8���L��T�V���Lx��m��j�h4��^L;��¦�?��dL�F��ժ����1��v("
\���p��4��������,���g�R�Ā\H����$��y�4��!3W���x1����%�R�\���]q�y��=b[���᥍F��e\��<�����gGq���di��@p/_�a���M����V�K(0��ń4�f9�ZE���ʰ��A[[[�N��l��\�p�Y� �9�R�R���]*�ˏvvv>I�ӟ޽{�ua��ٳg_^^�)�����B�`�y������w�\�d(P�aZu��B�����ϼ/�k��)�l(�UA��a5i��mY]��æ���~� ��D��i�9���V,�`���2moo��8��B�?����������ۣj��i"��}"��C6���ɓ'�ss�S�Zơ§�!�t�'''b���*��gf��67�TJh��N���- #?�9��Z�|�l-��A�.�C������\#�$	*
txxH�`�NOOi4]�<B�������=���Z��h4Ve<
��t:�D"���p����C?�#�V|��H<S&��L�sF��pU`�/�ՙ�/���@.-������D"B���;/��"���t��薀	���|*_��bM�A��.[\[ND� ��m hB�ϣWuޛ�%���5>�(��ϵ�\���+���B*P���J�v֝Q����7��
uy#_3<7�l��۷�֭[�L&�R�O���?��O��ϟ{��}�����].���8����:U�Uj�Z��$�+<���	��r�,,:�t:�k.8:�er�Jn��\E�`��d@���^���U�Wm��0��b+L7�kHl�h���[S܏�'��`���l6�\.'l�����QF"C�N�igg����R��I:��tgg�nU@�����x<��P(����Cj4^�Y	    IDAT�F�QJ$��0K� �D$��>::���d*d8pr���,e2ђ`�.�0X�\���j�E G���@0�`���Q�CT�C��7���?bH��t�<�)P<�x".R���=���4��z!�X��q��}��w��_����ӧO]��=:�� h��k
��f~�܋��[�\����������?�!,>Y-kXU�J���t��*;:~�p��[�\#�F�����q�����l���6�z=ᐢz�(!�c��9�\�OhY񹠭G���p ρ0����ޮ�vܯ��W��z`U�2ȝNG�-�?��e�W�*
��� Lv��`+�פ�C�޽{���?'��r_�����V��1��>��!�J}x~~N�ZM�e�R)����6��D�ЃD8ɳg�\nA\�cꖫ:m:W�c��a6]�ǋ���L��sTA^����ߔc�
�7;��'^~����r�ڄ���jj�&� ��%xP����\.��'w���9
��>mmm}�8��߿�wl����������F�@��x�"B��xH?�������r.�4R|`F&��C�I^�%�����%�&����EPP7�\Ch`�D��.�Q0�\�ʵ��1�?l^c�/�(
҈F4��DK�)�m�Uk�h6�����ٙ���V����ҿ���_��:88���3�	m�s&��e���+�U���%���`�����#Ӟi��x�hU���~�����;t��|���}��;�C�n��$�	����.t����U��(���-H�;���|��v(�������,�P��� �ׅ��手x�yg@ �zPH� R�e!�"�}�S�n| ��� e����z������lww���l��r��wwa�Z�~�8Ο������8ǚ�Ig��<�����@����z=WꟍL�&Ta����Ɇ��ܗ���^�����(����N���6���|&� 	����W������ұ��c�慝
6���g9�C�b����d�߾}����� O�<��2������trr"Ҏ0�D\F��y�CT�x�r�moo�ï�n��~\���@G$��ȄD�3.x-��6*�һݮp� K�A1�|����г�ѓ�6�6b\
�9��Y�E ���ɘƓ��c �X,R�X��qB��������X�Ϟ=�?�����_З_~)l� ��DճΙC���L;M����*6Y>��>����Ӵ�K"k�Uz~�ŗ���c��]�9�ٓ�++�����ҙ+�q0�����q�FtrrB�}�U�U���.wဖ�w���Cir�0�����?�{����*҅��r�D�|�3E0Xi���k�}-���|6���e�	OE��~ ��LF0���Hh���`ȹ5��^O���r9��ۣ�w�R�X����������S.�?�^\�1���T*��޽{�l�h4Cf����a��F�t��-!��N�.��.<��w�%	5���9�_F�-�]�e��d2[]�_-�Ml��=a��#o] ��u���#��ҭ[�hoo��٬���)�\�Q�R�$���������\.��h4������GGG�]GU�P���R��R�]H`zxK�I��%�]p����-�e�ǧ�� 
T���E�C��版D�� $p�kLn��gq%gK���UY0$
��x���T�:��j5z��1�B!*�J
������o��o���O��H0�\�l��s���4�<�&y����	����
<��71����i5��q&�__���<;;�����4�L�^����.9�C��?~L�}�]\\��g�ޓ\�S<��3��;&��p��(��p,'ޡ��kq��z�;�9��׃�eC�T ��9�ް�d34�Mi2���U�s}4��&"aE�"{
�`�=�E[ ���z��!
��S��'�]Ν�k�o���㭭�?�b��%	:99�� 6�i�h4�����n�i�X��񱈑��^����Mnj�L7��*��d�#lp]x]�kc����]�=�����.5��=��9�L���b؈1��Mӧ�b������`0H�B��y8��;���زj�3"���ӧ'��?9����Cyɣ��1~Ñ!�L
=Y��zO^�pYI<�T��
&��}���ޛ��y�I����w�M��(Y��ؑmd21h�	��#��| ?�p@�d���N[�em����}{?��7����@�,.�}/��UW]Uw�f�6*[����z+24��hu�9c{j�x���3C]t��=cU��,�=t�����*�I��q��Y\��p��}T�U���p8d ��G�l����mj\c�'i�g�OZ�&I�&1n {Q��$W�Y:�i�3�>笤4�o{3�m�hmupp�^����c��������gϞo�I�c ���=����b���9�y/V�Us�p�������gL�=��l�k1E)���[m�t@ʁt=�aY�n�������A�VC��t��Ed���X|��ï�@�F��b��@ ���-�������_E"�?<o��S���������D>�����72{UR�����mC�	����idޛpT�6�dK�ɼR�Yn*o�wV��yht�+^�.�v��/�2al_�Z�P��\���(
�VWV�H$��m1��x���(
wS��|��?-�ՃC ^��������b��{{{/M��~��
&����T*����`�\�d�l�$2��a]Ɉг�-S5s�+b����LJ$15�th���[mѲ�6V�?��#����ڱBa<hFVm������� �I;6�5��KL�a2�������Z`'��n@w��iV�<O��x�:��,2h�!�F�'�(Wʈ��F�=��dT��ŔP㭅[�GAG���F���ن�N���2\��ϸ6����\=q5��{����N���f�m�f��F���v~�h��R��4E}�Ă�*;)|&c����p�ҥ��d�w[[[��{Ѝ7�>z������P(�i"���Ύ!�B�k��3��Ţ���~�E�$�1m�xvaӢ��t���Z���yK7�b�\�E��y_w��O�M���ͪ��H&�H����x���u��)#Y K@p�N�q��e���ލ�bKpk��믿���z�����8R���ۓl��r9��>�kjkc���,
�b���l�$E%ԯ�}b{��F�ܤ�	Vmn�R1l7]@]�c��0�)r$2�6{������GuI�Gn�\v�q��<;�ծ�g��������^e3�t��m1.B�z��1]�uP��XL���
pm�Lj�{�6[v��Զ0�%�x3�Z(]7�y#h��x^m�1����6�k�/�`���Y��
|�R� &>6��>�:�#��Pok��P[��%d�ٻ�H�O>�d���޾������|�ߎF�����>���A��0�Z��z0D�XtO���f�b���m���������ï��,�}��Y��0���̳�+��E�LC"�@4u�Zէ�l�P( �I��:(
acc���w������/�˄��?�����動���{��O�@nP�v�kI�h�P@��A�T2Zh`,9�����UG��r^�Ŵ3�y�������Z�f ����ΗpM��e	~���gd0�chG��j�'�GJ=B���.��L��,A��w	N�蘧����Hs^���z3��v�{9���"-�i�a�C�<j0���%��{@HB��������|&� 8���Tz����d��I2�*g�{���YU����Ć-�̊�8�78�I��C��s����`��ϞZ��#�N����_|����=H��Aw�<y�����g�^�=2
vj�Q4E6�5����A���׵��y���Yݱy���Bj��~�ՙ���w�Բ;+1�E���ڐ܀�4���������tI�C��:�&p�4 $I\޾����;�p�wKp;�����޿��V���Dⶦ~٦�h�N�����H�R�V�F��N�Q,��f�n����d}؆%���>�n���q��z�(���b��\*�_����Q��V#A��(��G��/�>۝@}g�2�Wn4�ƥ���Z�EK��\s}vx���n��E�����ym�l<��g�M�l��ܳ�K{0K�խjG@�	�X�����'��`7u�}�����-O�� �ͩ�g��"V}h	�����u��A��?�*��3�g����ښ�@�t:�,�J9 ���2߯��E:����VVV����/��<���F�_�F�Ϸ��?m��(��h4fX���$A4�R�[�������ȴθ�̫۝����Y�$&�^�#|��j��
pm@��&��@�y���=Hٸf���eP&�_�(_Z����DD�Q���bee�x�h$�{��.��0�kE���;���_��؀��q�ƍ��������t*sh���`�f��@?`yN'�I3�����J���M�����c�be?Wd��ᰉ|�v)_���F��8�?i�`?w��4PBY0�����_ �IRn�7��smC�B!lnm���V�9�:�M�]���YZ��(�7 �� O�G}��$�uҚ���C�B�S�x"����)�z��֊ �h^��F�F�x`sHJ���z�<�R"޻
���B�\,4�S�����h6�f���.��UL�����C螡ϑ�D�r՜{<$�I��h4���-��m�5��쮭�!�����Kp;����w���r�___�tgg'''(����v���	������'GGG/��y����LZ����u s�N���Y���[��E�%�b��]��2�7�ZP[%�a�V5a:p�6���
"���:�`0@,����y��R���h���c��P(8����$�PV���L�n�X^e2�3�&Ս�#t���?����N������G���h�@0���C45�W���Q�{��޼Gi���?���z�n�kbT��Un��zUЪ�N�\__G��A�ZE��6Zb5�'(��Rk^r^v�U׶Ik�a��.؋X2����	?/C�(�v�JlK$�ՊD"H�R�S�1��T*�t-������#&C�zX�Z�"��!Ɋ@ �R����۲��r�l�V�|~�rP�$�|�f]S
	`��h�@�N}fm=g>ߌ����aٻ�P����:VWW����}�����)���5��
�kKF�3 ���h�ۨ����z3k�l��u^������&��ō����&%�����#Ә�iV9nӬ�m.:L�Ѥ#�b��R)�E
�i����N�q��
���`���t�7�.�C������:��gd+����`pl�.�.�\�D�4`8�hW�j5 0L���(��׳ڃ%�I��ĘfJ�z����]u�'���fȥ�O��}�9��_L~�0B0D8�BV���Q�`Jm��"A�K�'�읥33�M�y2��Zb�OsrX�cd����6�y��r��+��V"�����#�H �N#�N��V*����)��a{�Ѩ$S��Lĵ���0��"���Fͳ�`�;H�V�����ZR��ϭa>��N����	�m�k_'Z���|ckrc��q�����f�w�^��677��������?��O_lmm�>
}:���k��v�m��K,���8��"��>vww͐�:+(�ԉ~UY�Y��y~ξW�akg��sG��#�]7�e� �I�_[�@��q��q�v�|�,�.������D6���H$��gq8'�� �x��=O0�������Pj/���L��x�D�,J�D��M���2�f����{�:~�C��$�p!��bH$����B��_�T�@ue x��k����u4��ɒ�Qm���'���@0`>����i�)���|�.]B�VC�^���Z��a�t�V@8�N���Y���ދ���K�~���KU���&���$�u��՞��Ұ�a��n�P@&�A86��,�z����ht�V��!ө�~?m�ly��E�Ր1eۿ�j������f_H&���rƱ�̪�g��AU���#M����fǺk�ž7�;��k,>�[�}������p��7����?~���~??M$��jf�]ix����ɧ?�F���։�g%^���gb�tt����L�63|V����军5�<�(y��E
���Ŏӭ����϶����]�߿��pd2��|>�� >=880,�F��A
Fh{Łn<:E��t(@Rݼ8x
���y�B�&�M��^���I,�t���"��-[��Fc�[�X��-&(00������1�(d~����� �����F�����=��o�;A�[-@4�J[���dA}V�}�i s�6���nW�n�#�����t:m�uy���KG>W�\�g��h�T*!�H ���b13�� 
>;���}L�=�)�#��",�����.]��d2i�c���z���6�@��?�v�콌�&/��&^�Z�qP�y�{�R�
ǵk��~��7_lnn�>�H|ztt�j�j�.xt�d�`0@�^sX�N*�_��o������nQ�v�"��<D�ڦ��T�E>ܘ�I�,�A���N72���d�r9�@����N���f�$��ꔲ�<����<}���`��^��)ۆd�	*��J.,�k[��q�*Cp�k[�tl7��8�B�[��w�5�1�
W_Nz�z�����2�|�����p��h��P=��3���i#�`ee�YI=��Id��l�-t�{�R�V"���1��G%$t��EeL�
@'���e��}풨;����u���#�����yT3�Ö�.�$𥟴��:3��ms�)�!�U�^>/�Z,�|>�R)�4sM���o��6l)��n$����P�a%Ń,I�t\��r �L����;��Վ[�nݽ���P��#���#�j5�Z-�=���`�H�*��C����yDठ�y�t��,��E>�\�4�7�T�υ�=�ߥ	W�	�f�F�B&�7�;j��}�T
�x��%�=�css�����E$��H$r�����=|�C ��Ƹ�o���C&��1N��UBܤ����P�:1��	X��` hZ�~��A��� ���A� T�wi���{tX]]5Aܬ�\�$�"އ�
���$U�}�n�z�1�ZD��C3;z�L�Tq�9���"VD\'Y)�U�5��m�Lׄ�M*�y���P�6}>XpQ^��Zd��0�.h��t]����f�����)�6�ꇵ��.?K(2�.�St}"8�~��Jm�$5���-�s��X,�do��q��݇~��xns(Ҷģ�-
!������"��	?�k�"��<��j��M0[�O[���V��,|�Y��
�⦕�vAi�Q���:���K04�+�uJK)2��p��ray=ǻ�{��o�����߮T*fAQ�-�-� �k��jR�o���F���ii��VB*7��.[����z;�cF��\s���F1�p?�a�����^�E��Z��$�@��l��1�n��B�x�}s3�ԢRfw�;��Z�h����m�X,f�3�	�hAşW���G ��e�:�b'����Jc�f��21�m������^�R�n���~�E�L��E�Qø6�M��0���{��.;(�K��]�����?�]鰛F�� �N��l���8==E��5 ۾�
Dyo��uG\������������?Ob�����Xjo����|�x<��z���ժY�y�s��/.0��r�d2h4f���ϻ�M�:�<�g����IL�Q����<��E ���ˢ�3nZ�&FM�+���p���Q4���r��W7n�X��^ӑJ���l6��o���4��g�͗'� s�{��F����$�dK�y�h4:�X4�������fc&3�Cu��n��M0dN�RΖ�Z�������(����C�H��\.�&.ڵZ�Rɼ�M��5��i���Z��ldqm�    IDAT��|>�J��W2'�y��2�R�V5�i��.�˨V�(�˨T*fP�E��]Z>i�`w���kQ&H�ۮ����|�����C��W,��0�L(�,vix=��bc�}~Gܶ��,X� �vww��\�?7�������}By�"��VJ���A5��F�F�����󬅪����;�h�wK���?����|��_E"�ۃ� �J��WXh� aї��prr�v�����m�h뼄�y��͒�N#2�����j:Gn��4�i���xU�;M~q�߭���Z6����2i����bw�Ē�}������{��}���~�:hճ��i�ۆ�!cik$ɴ���E���"Ya�s�A�X�DLl3I��X�k�����C4�M��ɉr�Qc��4!�傪Csc�2:�}�������V����������f��T*&	�,�[����I�y�22�,@8�L ��Q(��f����������!�!��. ��5)h�Z��j �S*�ppp���C��e���`��fj�}>]���)Y����s�6||C��-w|���R�JV]�Yա7�MS��0r����0^���C�J%SF#Q��>���a�躒N���d�.6��&��`cc���j��yvU��bj4��:��sj����v���A�.����B���B��-������C��㵓�H$������n��=a;��5k�"��g��.���H��,����,_�7�y�V�z�*��,�h�'��8��ְ���X,�RgK�Q��X�w�yg�޾�#�H�!��^����Cǽϡ.Z�A���j���pm�P(�A�ƶ%��;�mx���2RR��	�~�������e��Rnt|o��K��a�h_��&jc�ɫ6Tۢ�H�U��N	`�9x�8-�IP:�>��`^�:okN?3�!�����g2�������@,���I�#�U=(�{��C�L\?t-�i�N��r����=���T*aww�~��]�FáW�(�stV �v�Z����q"xH&�����b `Xjv�T�=���~�oBX�&w�]T�U���/��C||��R.D�{�\F�T���j��X2����7��P(��\.�d"	�o�WVVA@,����삾�ڮ&�eG��^��ؒ+�:��z�D"�%����W�������U�X��b�f.u��z\>,tI��\�-4�U���m�?�0�gY�\�E~����E[��E��Mѯ������iuu�|�X��P�V�ht�޾�V�����@�ߣ��mխ���fD�N:�*�`V�̚O���jl��D6����6VT�Y�l����=���
�y{�"���~�m�z����� �_�f��b��,�9�Vh8E<���	���'�ʦI���g�&��k�J�������{�y�&����D�H$�����/چ������x��*�ϣP(�ҥK�T*X[[C8Ə?��~��G�h�Z�`
�)�����1�@���" �)���U���p���$��P�m����"���u��	2�g��x��� �������2�L���{{{H��(�X]]�իW���eZ��(��&E�~n�,m[0��Q˭�>�ܷ�a��|_moo/	��|D"�?��߮���V;H��U�t� �t�x�J���Q4O�@=�g|(}v�Ӽ����	pE�?g����'�Gm8u˅�i;�Lƴݸ��*�BH&��_^�vm����ccc����~��os����u�:u M�ɀ�v�`u����z��R��Щ��_[ߟ��wM*��[����u�^�%c���l����~�h	���M�Za.��z�l�d�4!�-�`0h@=���h4P.���4l�R�����x�Z���P�Ռ�իW����>��K��K�#F%z�# *792�,�u*�CR�~������뚉��
[���p���ч��bM��n�9!@S���9���l��� Fc!ȹޯZP�ܑ�T*F2B�k,{�x�����z�n��G�amm�J�z�����rX'�I��e�Wఉ�g��m�[�負e��~��ϏF��/��7t���;w�<y�U�۽}zzj<�m�bM��D"�E��������;�s>�8o���Xm���k����9��?�"�y����� ��ms0����h-�g�d�d�T*�|����d^�vۀ
��VK'����p��aC�y#��a����C�ٳg���XYY������ahC�G{۞�%��!� �n��{{{�T*H�RfhG۶��U`N�S��b�@ �J9�m��S��d�J����ҁM���i�W�:6��*�%�f߸q���/p��U$�I�Xۖh�p��>����&�f��}� @T�b3�ߏ��*��*���qrr��m~]�m!i_7��)�	P�m������|����#,:C���l�z�^��iV���IP�6`JV����&P�BH$�#1��J ̓����z=S�$�I
��6(峣d����sĂ��+H)׈D"���|޿�z��`yCG �����m4��5�k�>;�^�`�P��e��^�:�>+�i�-�@����� �y���4�:�b<�2�%Q��䢢�7:�ʛ��=�`��i�`0x'�|����F��Y8�]���
ہ:���`�����Ȓ�T�K��Z����Ԁ���}����C�G�!e�������f�u� �o�9���"77q�e9�D����p8�X,f�k	��|6T��������"��KDga_�qY��
���"677��{��ƍ���B*�2Z�F�a��N�k��XP��[��7�d�%�""�˙!��ׯcoo�~�-<x�����Ү^�c�N�r���>?�˥T�@���,$ ���:~�N��Z��A�Ht�EH�R�.������l��Ė�M*��0�jϞ=3�n�����6VWW�DP,���������u9��2�D"a�9�������
����ԝh4�do�౶�v�믿�2�H��}l�W���S�	-�܊��Ť�3F��-��kZzڢ�T׮��-��k�HgU&�~V�_RL~���ֆ�\n�dR��~���bqY=��ckk��Ç��F��Y�p3��A3������%�.T����������X��j;Z��Z�J��*�z=�{}�T���!(ug`�W�����)���N��ٳg&A���bss�t�l��HĴ�	�ժL�(��ل5�"#�ɠR��\.��2�n�4�ꟗa��������F����_��Wx��������d2#� �̈́+��7�//���K]0��=�2�Pm8�,�����(
������8==E&����1��[j����m㙷�e�]�xoi�/� �NS�eڱ�k�p����!4M|?�G�� ���&��΄�OjϥE
����p�f�� �n�vS��6��K�.�;?�ӧO,�_�B�|�uQ���W�3�֢�������#�J��!��<����H;B��o���3�ã�+yЭh�I���Rrb���"��y^��`g1>�=Ϡ�<�x�e�<i@���:�d��H$��#M�����T*�d2�D"��'��#���l�6�ܦ>��Z)�Ҝx���&�H$����d���P��qpp������ޞ����d�:mn��~�R	���,l;�I#t�ř���*���x`:�������lll����X�!����j��A�,$	�W*����y�n,��ƖJ%�|>\�|}��������alm--�#=n�:6�ɠ7�8@G�1&��+�J9l՝C��ա����l��T*8==����O�F����YE���I�Y���<����Ǳ��>�}����^84�Ca$I�}�Z�v6�fw�@�ω��`z�\6��"B �{����h�}o�B����5���=�n|�8���>g L���t̽�∱��tz����#
}�D>��r�����l��K8v�;�֣�Bo�S~^���p��k�����Lw������)&-��)o4[�ɪ���d�����r�D"w���*���o��F��k��Cj���ڢQ�Q�����P( �H�V����?��#>|�R� f*�:C��dB����v�j�@�wJh��N���� `�t:���3L�իW��f�����.|/��0��L�%���3�dRc�n���ka��M B����~?�\��[�n��?�͛7Q,1���p�����B���N�c <}��7��h��F��`0����'��5'�H �;>#5�h:m�
���}T�U���bE6ySk�=�Ţ�A���j�b�<c����u�
X�ժ���A��>�v�H�uYm��AKƖ`U[�|�&�Zt���g�`�~��r�l��|�"2�L�X,��]�b��jW��h #���|>o�	�Q���f�H$wC��r�yK{����e4�MY����}���:�x�v^�0��Ս�7�F]h�9�󾉟� �Y ;�Y3���l
=.Vd��b�sB(�W(���o�H$^��p3��)3���2b��S�L����j5<z���=���1Q( ��,n�dM[����S�B������h����0d�Q� �îʹ��5 ��&�X��7�4���h���������;4!�P�"�PPiG�.�ϭ?O�S�ǃ+W���?ƿ�˿����G6��5�-�N-&7v:��u�������R	�R�H�k��	�������(�XYYA�X4l���E�X����Ѩ�
�����R�t��53����c���
��P���B��7xM�SI�������726a#�A���-��.��0VWWM��6�i��+ȶ��Uʠ�,�j��{�sVc���a��j���622�,��>�C����`d�fvK���z�9�����}{G4+� P'�V��[�=��I��uiq	�9k7~k<dO����9[��{a���u�D)e���8�ɤ�r!�Ɩ&M�=ϗW�\Y..o�P�/���Z���7^Ն򞢶��Z�V������1��b��˗/cee�p^�׀ ��	`	(��0
�`щZm������\���۽��ق�`���c�.���b�����sA�u��r��~�}G�C�ɠ�>�v �0kAf���t�����?��|�	>��C\�t	�Ph�#�n9��yϰ����8>>�ӧO���c<y�;;;�T*ƪIeZ�������sÎ������:���q��5\�~݄J�k6���ZgE�Q\�~�n׬UO�<q�j?k��!30��	l�+˩r2�����:b�K�?~�z�n
%)�۟]�
�TM��#�5�GYZ�/�R����V�v�R	���ƃ����F��Ō�/0vi!p�}���M�cK����/766���[<�����`�t:}�\.r�k�]%��c�2ɉ�MYv�{�Vp����c���s�Ӓ�� ���U�e45�g�����x<�t:�]>�����>=A��Gp�-V�=�*0��Å�'�K��Y�|�t�!ন��j�Ł�H$�Z����iS��D�ZE��t���!�Й�%����&)����]�Cd�Y�8�ơ�D"�L&��oҠ�k��#8:#:�I�/?۴��y�R��$C����?��|�	>��#lnl"	��Y湧�b4���Ϟ=Ã��������?����=�z�Rɬ���XYYA�P0:L 8>>���a]{���,���������O��t���ɵá�9c[3
!��ᗿ��a��!vvvZ��nm6�mh�Ivܰ�<�䋟KX���/��8::���a6��i��S�z?(8U��:cA�6%�ӯk\�����p8�`8��30�aeeŸ��z���`80�|�=� �����<�t�����-+++w����/��mF��N[���y��^p;im�6���m>��`����P1�w�/���<>j�|ئ�{�qZ�|��-���$+��&���#������p8�,���w2��G0}nt�N���ޒ�}��+�����z-�4X�Uj��{2��o6���A
}�u��Z�$�ժ1��V��}Ӂ"n��Z��>�	���g*?��AlX}�n��������Ǳ���[�nᗿ�%�����ݞ���P]'�={�o���?�w�}�������������E��i�r9lmm[(�U*b�����v�����駟�E�R��ﾋ��-d�YG��A3*	�B(�F��h4P*�pttd��!�E�z*{�23�@��[t�j�UBC@��=j�Y���&(P��/�[��m#6,~$lο����Me8|/�4�'��k������<N/_��g�\�/��:P�{C�m�������[%��rZwm��a�^L�^�,����E���~�9ɪU4��q�����"*`4tc�? �D"�����T���_���i������nT���-$�ǃZ�fl����ש���j��ƬL��1Nd\uR��8_����n��(e��2��r�`�%��]�%	����8Z�Jд�ަ�F�z�rٸ&�5�$��Ϡ���ӸV;��f�'I��� ��"�\��k׮	@��C��u�?xnF�NNNptt�{��������ܿ�?�`0@2�D6�5�Z�X���._��+W����ˆ��v�888��'O���c�������X|��eT*���6.���������|>� �6���屽��Ǐ�o����a�&ܳ���C�z���ӵP���^b�,U���z��9e6�z�J�L�s��h8����Yu���u�~2�}�<^�y�}#�T������^��J����D�Q#��7�{����E�p84�V���_,����)j?�CfZT]$�v�0�����&��2���i���'����vsP0��ya�
��h�`w9Q����ރ�H&�^ժr��:'e��Q!�m�V��R�d�	'''��E5�^�]tM^<__����F�4,p�%������r�=KL7H�DS� ���h4B*�26`d�5���*�9�&�>�|ol�E�Q�	i'�Mj]�u�܊SM��r�y�&>��#\�v�d��8�����p���C|����_��o��?��NNN����B����-3,��d�������E�r9�R)c5��z������mc�j�\���]<x� ��_�_��_8<<���!?~�>� ��.�����@��~��ᇈF�x��C.�l���ߴ9�p�[��R��5�㇮����sK 
�+x���� �J� <~m�릫�c6��g_a���H��9o����U��\�h��N����C����H�ӦCD}&� �~�<�����CGCCA�/�� �x<�%�r1 ���r�`�V륢��%m��"�v��W˓2��-�z݂|�:v��N{�Bx��v�EW���B(R+#��<�UZ�.��ikzI�R�l�=���������S������ �r^��X̀GD�_,7rnX˔��!7m����M����x3◿�^���V]y��4`�M�8�cC(��x<�F�I�+�ۭp�f'������q�����ի(���|h4&5�N���޽{�ӟ����������7����/Z�]�~� �B����ud2��`0@�?A�8���`ss�X:u�]���cuu>��|�>|���Cܻw�����j�裏L����y?�b1�B!����֭[�>���5��M+��n��o��,dx;t�ϯ=_� ���f%������������;89{{{&X�������LZDj����iv��{��"�p$V�=��B���]��������w���Cx�H�x1������s�|��rcccI�\����}��z?K$�9<�>�>QW�I�PQ�%g^��<@�	��rf�y@��"Q�g��P�.�$=��x��(o@.�:9��	ꋸ<.�}�G(���3L"��������ҹ���ظ$�I$�I��孛;�bޠl�2Z��U���+LӦ*�U��D��
�    IDAT"a�����c���4=M7b;���������a8:�Yy�m��mk�H�	N�q����B���Dw�(�J�駟p��=|��x��	�ժ�~��G��o~�7nK7���먮.
!��~1������H$�w�����h4�|>���U�Es?��&�e�Y\�v��cz��8�=�5��l�U��p�?/����=���v|�]�t:�T*8::B�T2N56s��A�� �熌�])��gP7�l6����sN���=�M�ӯ1ͰT*�q�<��p8<�x��'�7�U�!k˒`� G>��s���/���m;�vp�}S��$Y�5r^b�uc�i��y����-��Q�n��h�Hz�-�)j{gy\������������Tʸf���K��F��χl6�T*e4��~ߡ�U�j��(�	R��v��׿�jٱ�zr��F�޾�H#���	K��F6����x^ ���9���( �?n:C�Y�vh�OS��J��id23�CP�g�l���1~��#K��>����}��wq��-��׿ƭ[�p��%#'Q���1mÔ}�x<G���X,�˗/;����;��o���1<x�+W���͛�y}��-+�U�^��#�ÂL:#��q�n,���Hx��Ǭ��;���k'���m{�j���w&�$ ��͡3e_�	Gu���v�H��f�"��Z-T�U4c��h�Y��=��Է��~��A��|f�w���Ъ�ב�+lk[ w��_�#{��(1F�����\�q?�� �Nc�9d�H2��<�F�.z�M��
vd��jږ��
m-܋���i���
7mAq��🀨�l�V����Bfs��&�Y�n��q���D&��nZ(q!�,WڲR`�^���T�!ٹp8�t:�͍Mt���͕�Z�o��Q[3ev�&�.>ݘh�J^ϋ�P(d��eZ��F#T�U<|���_���_������1r��^����u�����/~��ׯ��@V%%�yx}����6�h;�	�B�����H$����\.�p8�����8::2�=e�X�1�]��>}�<0E�[�4g�Il�ar}/6k{P� ��7&�����5��LǄz�n���@ �h�SBP���vþ��CV���V�U�R)�r9�r93��������rۇ�� "�����R��t�����U���m���8��;��V����%}�?��=���F?/�L��n���4Wnm8;��?�2ߧn�6�X�a! #�fG�c���96`��N��Ry<`�h��0�Δ�\�pu�WZ��tk��ȍ���q���5�n��t��9`���-0NU[]]��ё��O$db04-e�;�����l�,]֤���%R��\��+W�`ee�@��,�ƺ��������?��NOO��q��5|��'�q�._�lǼ^/����}|_*���NvQ�������43ڵ,>}���moo�
���}M�t8���:�\��G��ѣGh6�/1��4n��8I�
�\��S}Ψ��9��p�7���JG��Q�������#סCJ<؟��s��g�^�����T
�B�h��>�j����ĭ�������C�7>?z�����ܳ�� �T���g��$����0��X�d/ϊ�Ϭ�W�����J>�;IOf� جӮ���
]�4�\���ߗ�ż�fv<Ϊ�S��C�\���	J���9� �V�9&�څB!cwD� 7Tn�l�꽤�&�L�\�	=m�25F�Vm<G*�2�f|ύF�,��Ec�V��V�h����yϹ���R�yZ�ô������"���ڵk�v����I���{o4���������A���ￏ��{πu�`pG(r�tv�[����V4���qd2\�|�0����888����������-�a��P�@=.?�;＃�O��6:�����Y���K\[��X�>�rMv�e�^�����`n�7*��;��+@�:@0zzz�j��X,�B��xcQ�,ݴ��h4P.�_hn�ͱX��X����-�c��7�z~�����ﳇ��z^�~�����׉���}5o��_䤿���ȝ�Ļ�X�����&ȱ�G���Ќ��C<��bѓ*CI�T	:8O�R����c��e3��D�5�"������}ÆRIG�z��BQC2^v���X����j 5����t�x�r3��'��ŐL&qpx�F�a����Çs�slM_��y��]����ad�Yloo�ҥKH&����9�T*x�����P.�����Ő��T ��-5��*Y���RuҼ�d��HR�IF�C����L���h���������qxx�����ʕ+fxKeS�����S�EB���ӹu���v����5R_S�Ke��3m4����3�X�%�)[�]���ӗ��������H��(�y�#ߋ�"�����h4��Yp�`�Fh6�?�Tc2��]��f��k�%��y}�k�[��M��iC�o��򻝐i՞[��E���1�nB�I����9b�f&�l:�5���/�}�e����mj9h��F����p����`�\kkkh4�t:8::2 ��U�,���L�ޝN��i�������Yk��i}s��Y�VC6�5��@�`��P"����������z��l1�7�co�/��v1t�WOP>/��6zR�έവ�LkkkXYY1�
�'����x��?~���#3�
��J���d��f�����Z���0 ���԰���d��y�h2];��-
�~�:��w����>4����"h��$�Ncuu�|�X�Hh�ݝT�O��qkҹ�]eN�J\x^�5����n�Z/�$�E�?�p�n��M���S��֜��}�D���L������*VWW���e~�z��xv��hT+��5f[���L�]MJ��Z��q����`�Y(���0u�	��/ul�;m=t��7c;�+a�7����ބ8��K�� w��/�݊��mm7[�j���-.X�ۋy
�;������h4�M �M�����$(�-��Q�F�X���x�V�VQ*����C3�c0�Գ=�6�n�=�J$H��H���x<h4��aܮ��G����'O�gQA�5����|(�J�f���^���32Ō�%�H�7����tZ��n��M[,m��`0�|>����R)s� �̈́`�R�`ww�؁q��]���a�}�CtC�{���3��z�nd ��8i�ʕ+��r���5�����W�B8ƣG�prrb4��X�1�b/q�,�� �� �H���<�t�}�w����,*�$�c��^�����Jű�SO�R���u{�f=~�*i�Y>۶ݝ� ]��H$�^��j����Cd2#�����𽱸�������9Z����&�#W�-��%��X���ʝ�����2��=���L̺��ऎ�<�>��^˭Kb�ɷ�}~��i��<�H��n�H�.��Ν�	p$(�u��vх,����i�,xZ��ͦ�	��Q�����1�g�X�ժaU�m����Ѐ\n������*��FL���6`tu  �~_E��uĩ����O����3�Вmä �MA�P2���wW[�p8l��D"�0��B�L:�h�1rw{{&Y���"Q��P�T������&��ٳg�t:�35��bgg{{{ƙ� ��"7��D"��W��[ڵZ� .�#v.�&�1*W�κك�n��n��ʸ�O��s��'J(��\޳�����U��D���F�c��l���H�J�V�>���.�!�����ʆq�0����d���=g;i �^����`0�*!fX��m��i���!��>L#޺D��zL���1�F�\�5��a?��9i�wy\<�߭��v��{����l:�u6y����Q�T � �V�e@.��|�v��؈;�J���*<���Җ�����<8����Q(��:::���)�����d��q �,ӳ��e��#�9@�Tݺ(�.��bEm1�������� �Z'''8::���1j��� 666p��M\�~[[[����&|��	���{|��׸w�Iۢ�E�\6,�����c�����?�͛7��փ����i��{�E;L�����n�
v����\���׵]$��g��#���t-��*�������^$�ё�@�p��z�5��Z����s�k�(j��f,�����Tx}���{�퍪��afѸ<����in?�F��=48)��u�����INK�{�e��iNXQ����2|�w"�s5{������'��X~���E�ܨH���S��~��u7W2t�q�k2q�N��U�O�Wv
��j�h9�ʹ�{�f2�|>d2�1әNa4|��E��<����`��_e
���LP1���A)�_��Y L�A�f��D�Q� ��f����C��홴�\.�+W���w���˗��f�`!�'�<x�?���>=zd N,C86S��1� a<G.����Yg���k�h4B,C>�7j^Wu�P��Vtt|p��ڙ�=��
��d����t�$����(h˖�6ڹP�F>��#ߋ�=�"��`Z�	8�!��l���].��a�����q�a\�C��Sv}ۺ��c�L��|I�\\�N�,>K����ϛZv^R�y��d	�u��Kv���y#&�Ncy�l���7�ͺh��R�{�.��j��L�j�m��M�������78��f�*���P�M���M�ml��,����NԔ�e���`}}�\�.]������i������5����&h�_� 
�CZ�y��:(��N$����=8�F�VC"�����q��lnn��*��� +_�Vqpp������nwl���+���x����x��1._����5�B!d2��M߳],�u\��v�/����� �i1��`���:R�J�SA';�,pȓ�6���Z�u
��RZ̵P=�ʃ���V�<ۋT;���0dra8F<w���zm�bq������Iի[���*ٲ<.&��D��uő�:�;H�y ߢ�Y�g�@���'���g����I��E���2�ua&}�,vB�̦M$��˅��x��������#�ŕ[R�1���0���Y.��j��vZT�In���S���jԾr����jùiS�I��}��z=�����ÇH&����F6�E:�6-�z� �9B5`� �0�����,���0�5ƎQ��yA}��[R�'����z���Ƴxmm���/p��M�����2�@�0!+��b�]�:QzB�^��T*�ٳgx��)VVV�L&_
�����TNj`���k�Y�x[��,�f{��k����b����&�y�$����}<� �j�L�����V�����b�^G�Z5]�fG���fӤ����ӁE>���@��]�-�[˛�����v���=�~��ԅ�P�b�`��}�,��m㘦�x[�	�.��\&]d7&V7�V������8� w��^�c�R��DeT�1�B/�e\�{}��%�Z��?n2���0�'�%� h�u��\u��NF��4����6=zd��D�L�`�jձ��������%�n��0vG ��S�nk�nº�/�������5O5ӍF�Fä~moockk�B �W�Z�� �\.�B�L��)�H浮��8::���j��K����"���f�RY�-�`��F�R��̳�i+]]&x�Z'�ia����*����T*���5
�|>��u3P�r!�����Du��9a���������^��N{�v��]��Y�v��F�a�)��v�P�% ��_J.�����z/0����d��Fw^2�U�>fu��Rݼz_�q�Y�/B���!�Ǣ���I�'��-"�	��d���o�����x�A;
����Ço���|N�a���tN�7�f�Z�b�Tʰe^��vGGGh�ZH��㤡��������l��n;Z���F�6�����.n���rk���+�J�����n�.�i�n0���3�á�~��~��h7��(�����us�/uJ]T�
��3K���@�B�J�v�D:PS�g��o�u�v����?
9�7��X�q�.�r�J�Zʹ�m�K�F�)� ��u����c��h4�b����M\�t	�z�1����Z�I��P2d��N#ꞠmZ�}��y5y��Tu
��z7_�~~��$՝���ռ����A�����h�Y��=��.'߻��6�n�꼯�y��E�j8���ydG��[o�899�}����>|hB�x�S��6���]f��C�=�n:\7�ޫⷳ��݉����$��p�]�W��'y����.�[^��hԘ�s�hy\����|���ns1�3�'�
p	)E��J(���
b��� ��6�岣����ƀW�B5j��H(��{&xP,�Kv �6z��0j�ɓ'F�KЭ��d29�89#~9���v��Hm"�e����7l�3?7���:�E�������Fz��C�h���v�O1���m�6ixK���EU��]��1���
��ς�k�`0���!Z��Ѩ<��l3�dee�$��M�Y��I�nw>��!��lf]YG��}j;m�HQ[-e�yo1y0�L"��9Ot�R�E�� SKf��N��1��v��h4j�(�C�]%x�|�Ѫ��%&*!���a.��KmV�������`0h<�}>�Y{��W���@�$z�;��4��6�����HW�,<�Jxۭ�Yg�P&U,n�=Io�ĩA������q���]@�u-&�-�RO������Uc���zqrrb�Q:�B!��!t��T5�V��`s	�Tk�B�5�=G����#�}�NN�~��"���C�Z5q����Q���K̷��S�A�{�`����m��0�?���!%{�jֽ��Yϵ��vK�F:��������^����S���#�LN�/>���,��<S�`��%:��itt��Is�;e��(�!�;Q*�c����QM �>���2zWS�Ѩ) y-)Q�.����@ ��ک���];�Z,���^�9Z��h4j�9x�k���i��	��4lvVFwR��2�E�����]��>�/ټ,�q^ ��z*�geLsx$pQ�x֥��ܨ8�����B�Bf��R�Z��4�M��Q;�O�)�ɂ/�a=_V@d����:�}ڹ�d��TM�>+��K������T��������8::2�4��Ά�:��f���I��;��9~�t�#G�.�.4�����nzh��b���N4�N���c��p���.>|��h�L&�����ys�T�J�Y]�Mْ�Y�m�h�?�X- Ȁ�3�p�>�	d���0��6����DLQ�J�P(���j"w�={f�K8��,4Y[�$BY�2p$A��8�wur�[�j����U�a�����r��@C�������x�*���Y��y`�E1�$��_��\���a�:���Rۈ��dF�r�%�����b(
��qee���� ��W���J�M͎� �D��)=O���>�\.��n�S�k�B�{��7Sz�j�=�2��!Áѳ���n�
6��r(�-���g�^/B���ܧ��8==E��0��d>�� �[�SV­���zem���5�9u� [���ŭ2�|��&jˤ����g0 #�͢X,f_�op�\��qpp��O�"�T*O\�,�*����j��+&�D���scF���ߵ��ֲ4�ܵD�aZ��0��ՑC��@���X�Tʤ�q��h��L&������5��dm�B/i2m������V[?'Y}�����O]ez�x8x����I-�tX�lt0����䏹\n��\��^��M����bF�r5�#�M�k��U���G���r�?+�E.�,@>�/���6	�r��pe��~=grow:��,�p4��!�������x0:[{>�ϑ
�L=�Tr<Tx||�N����T���b1#j�5x�u�F�f�YD"cie�r��"0��Wj�wP    IDAT�"� ����)~����W�U�@�%Ռ�$�N�+�h[�h!����::��x�EO72�,���d�l6Q�Vqrr�z��l6k>��W�������Se�,3���  �8Dh��l&��l�\.�xX^'�j����j�ێ���SG��&"ف#�`�sM����]��<�\c��b��<�����q��iӉh��(��n&�^ڵ�z�&ҹZ�������S>�����D�~�Ԫ/��M�lW���}�{����ڡ��Nݳݭן2:��s���/��p����~����Y�$�v���u��X
�����?m��yU*
h�̊m�I[W�S�PC�./�P���߿��ɓ�	F�����*�f����=V"�{���f2�T*����H$�Lo(�`�iV��w�����D�[:r���0��������ZOMk5qj�zO]`(���|(������0ٯ�phZ��l�@�l�
�yh�.y��\�����D"H�RXYYA�P��?����#��N�MЃۢM�0�J!�J[�f��h%+�a���Ӥ���b��NNNKh�zٛD��������oUo�y�H�uJ@g'>j����f���ՠ�pӡ�P8�p��p�iUϭ�/-��%������T*�7���������0���F�`?Gt��k1җ]��Y ����|r����>7ꍪ]�&Hj������v���`p��́@��q(��p �ʼ	O}�n�Yd�֏i�T�$��t������$�<ϊd�`�4z\`�k�ﬠ��q ��/��K�8����p�-]����p8rX����v�/6�N����F#GCx}^x�C}^ �|��� �������v�~��x�t"��aq�>?��>�#�t�Aߑ�6O�/Ձ@�Z5�-#�`
����s����,���dE'y>N�6,jkC	 T��L&�J����qxx�G��ʕ+X__7	Xn�0����$��4�*��d�b�f��?=���ّů�j&�W���z.'K=+7WuP��m�Ɛk��U�=%ԻV;�gZ��pC!D�c��T��ԇ�ir�@ �t�T�<?��K���qzzj�7�|?�`�F��I2�2��CW�⎅�2�rS����
XY�i:��\�q����3u\�[�������N����V}?��^�g���rKNs��@�<L�\{�d[�J w�r^�v�6c���i��}���\�)[�Y���60 P.����:��|���ޮ�j��V�ORad�d�^/ڭ6�(���;���&�L&szzzj6e�U��u�h���p8t0C����jF֠���@�� �sGIaSTn�,��>�w(�Ԕ"��{$�����Pj[��	������.ك6n ����ς���ZJ��TM���G2�D6�5r���#<x� X[[322-6��B�t��^�����@ ���ƙB��	�s�677q��-���;H&��\�����f�������b0�s�a?&*3�a�h4jΕ�'�v����h��su>�#sU��g;؆�j��Br���jЮ�þ|y�5m��<�+�x�����E,3 �N���%#�H �NK2�H0cS0R�l2�[e���uO�,���?�;���?�<��A��J�b:\�?�f��aS�ұ�u���R�l;-$l~����n��_�b�$
��^�N��Mc�ra�2I���E�=,y���� �Je�ý �h4�����>99A�G<7?�p8D��r\?�׋^��as|�� ��(���<I&�F��hV��e۳V���"F�V�U�$@ J�r�lZ��jQ�i6���#��F�cM��EG���c�T���LS~2��	k�Z�����2�N��~�o��5&�#�M���[�v;Zk��{�m�T*899A�R1f�ʀ�z=���d�}��)��.��ױ���b�h����ع)
�v�~��w��O��Z�:�V<�������`ss� OBj�sF uxx�Ǐcww>��.]���r���^z߲x�F��4�I	h��Ƙ�_����l����1��`�)�}�N,�:�B����a>9��b���Ϙ�lFv�EAn�7v�p"��hd<�Y���aG��s��s���BF�¯ib�$�J�����l����]v/�qrr2<99A��0�>#,jx��|^�3k�k�h�y�4Bs3kcAu�9�MR����z-]�'�B����"�Ŷ$cI9�D B&�R�,#�����t�F�F �H�l�����{��c���*��!s�D8�lXW�0,�R��e�-�p��fʹ��h����Ŧ7��_�V��a���9cl	8��d�؎��$���l� �V��V{z���m��v�״v��sJ@�N�`���_*���bH�ӆ=�R����}�P(��+6��ߏ��-D�Q���bkk�?Ɠ'O����r��N��B��[�n�׿�5nݺe~Fϓm9�Z-��Ç��ف��Ç~��7o��ի�f�&p��:����lZ�|��:h�"W�.��r�^�m��';���<�Z-#5Y[[C*����3Ҍz�nB1�yQ	�_��7���v�f����&�|O*A"�Ԁ�	f�N�o�G(k�����ڃ�>��n�R	�t�����?��%��~��ӟ~��s���{��%*)�s�����M�L������:����NP��4��6&��&�-���˜���F�P@<7�N��ݮYdvvv�����\d��Q�T��J�~�h�px|�G�x_0B��Z� V��/���l�2�8�z�8::2�G�8>�	G'''�V7(�@U�UÌ��k�`�.0#���Ð�`>��B� ���Fs-�H ��"��!�J�4������dib��õ?m0����^=r�W��ܕCWun&QT�LY��7�A��n~��s��|���~��R�|�e{�D15;Wu�s���������&%�,�a�C���yֳ��k�g�,�ժ��)Ҁ��C�H�H^�w�6�L�����@ 0��`9����������ױ���+W� �����xgggh6�X__ǯ�k�������ץ�=Ry�4<�Z��D"���}��ylnn����������.@Y{fjY��z��g6�0�;��д��2�dk敿gԤ�Hcj��ݝ�����n(���2,����Ƅ@'�i�YK)t����v�h�F��o��4��� }|�Ã���6w�s�'�Z-�E\�~}���}��Ӽ���n>������4��	�H����AB���s!���"�*����Lskfi���qQ���qQ/�Yw�$���1�80ٵˮH����).P����]�O�:==ݍ��f�Y����"�!70�.�v�}���v.�V��Ѩ���������e7N	�G4�'�?O��~�,�EPk�dW����#-C>��b�� h���fI�36ͱZAk(�MZsH6��SG�2�,Bw������i�X�v�eSP�T�O��]#Y���-���Eaee�h+++�j�jey�\ ���:nܸ�T*�d2�~��X,�k׮a{{>�o"C��k{6JVx<����x뭷����o���Y��02�F��Om�f\Ќ����(-0��ꪀf��v;�����W�-�/��q�����觯c�^G�R���@4Y���Rn�g�s �����a�7m����%�h�������N��F�����#�xO:�1����|����7n�Y^��h|�j�v���D;�ԛs��*0�}?��y�Y ׬��X�3ʧ��Eӟ�E�63�k��λx�A����m�`\���s)�x<od
?{�I���-
c�j�M�s�YZZ�����	{�`���|�L�ߏ@  eJ�X�zj�Z-�����7js����m���a3�Zr�`�O�G�����,x�n�N{��j�O��F{<2k:�r �C$�M�Ʈsjy�ͦ0ze�*7�����N3��x�^����ʕ+H�R�d2�V��f�8==���6�y�����s���G���8y�kkk�Ec����͛7�)��vZGldjȈ���8~��G�J%�������x������%�=2���N>��1F����af$�ʋF�mW�c�u���D0��g��m�f��B����`���b��L&#޶b`o6�4�CPf�����Z�;�h����Ze��P:�ٗ��zec��д�26��o���hݘ7��v0���	���:�V�����J�� �ˡP(H3"�2��Y�ce��l�%��������V�"��4��9ӚZ���/�b�2R���2@�,@;K�k,)��^�'�4�w�ݒ\e�Z�T�F��Ӱ����w�Z���'���E�@�eQj��0s��LU��C:����T���8Ҷ:f�����b�(`�����ӱ� 0���1�T��9��sR�63��	���fz=]Vf�6���qL���P��B�VC�TB�ەF�tYY۰�x���|`�u��G����V��X,"��"�"
���M������2���ptt�P($v\�b�t�\N6/<�f�9�i�.R��pD$,�I5�����aS���)�<y�����vܸq��>666&�����c�V�	���3�j�|V��qQ��
_�LhK8cC�n.��l��t��i���M��	��rY���ڍ�Z��qй�b�HU��R�����x9�ͦ4y�^��~���̯�OX�r5mt�����dy�8�V��;>��n>��*��Y^㋲�b�(�7=g�A�j8�O~ʊ�4+Ɨ5!��^�
���^$��2���N����X��j��h	E��i�$�A�����n���_��l~�l6wONN$AJ�OnX��<�2;��~~��^�%{	�B����x<h4���Z�Xr/�&����˼^�TX��z�p���,5[M�=8]Ι�W��#꺴ק~i�1��y}�bS~��o��e�b�j ��z��?����"�����%�^f�W�?w�da3�677'<m�l���4���m4(�J(�JH$���X__��.-16=i ����Y�]oN�B'�I|��w����xoܸ���-x�^��:�Y�8��y$�I����X,��nK�@G�.Bf���fF�F_�i��ڛXK�=�afL?�GV��vK�	�C_W�˅d2	 ��\�cֱ��� �f�=Kp[�ץb@������l�K[�q�&�kP��F�R��xn,��Z�T�ը����zodr��U�Նltt����1�lJ8VX53V�. _eE]'��"�[�i�g8`��v#�4+�Ӿ�ׇv�ߙ�f�o�cm�5p�d� �,w\�ZM&(&Q{Y�V�N���x�}����f�yůL&���d�f2�J%�|>Ytӕ(����Y\nv�}��0��l0�\.�����'�n�;u�0ɬ�TEO���k� ȢF��	�~�\����fo9���Uj��V��~�>���V��֕�nh�FK�]6<&��.�k6tڳhIF/V�%��6�?~�ۍ~����Mx<��'�v���4���g�Y<y��N�\[[[���XZZ��'5x7�R��m����J'''�����'''X[[�?��?��?�`
������j�����ա�n�}�6f��fD�N�# �U �����j��v�����Nh�f^3�ds)1�=����ʊxޒ�������L$�1�L<h�3�C>z���,+z���o��ɺ�"��zw]e"�&�Kpk��aw�7�xv8odr����?N&����7�|L�7�{8�
[o�ɦ�V�ɽ��ޚ5fMk"���^�2z���{2:���*6�z��f,�q7�'������'�x�l��Bj<�5�n�jUX?	x6���������M蹆�!��2����5����'�Zm�P(H���a�Z��u{���m�U�	��t��nD�Q�z=d2��yai��&�~?l6�~?���d1e�7q�qg~�V���AB1���0rL� ��ǭb��lD �����8����}I�Z^^F =b��F���L6��� J�z��$7#;��/�<�^Q���%�$h��z8<<����D���"�*���bA,í[��1��h�V�����z��������7p��\�vM�H:��� ǒ��ku���f����w�T���>����o�A<���ǻﾋ�>��n݂���j���,h�����!���;<}��dR�x\��Y�pYyͺj�\�>�mTx/uH���E/؛p-�$@gy���%t���r�#��d��oC�#z�ݮ��9�Ή`��8�S�4��\��f'�67��d�^/��h�y}y�z��c��S�9���>���|>������ޗ�n���7+ī�����S(���eCL	eov�����6�ϣX,JJ���ޢU����`/3��HO�4o�yaf���Q�Ӛ�~N]}��5˃�wb�����X�7�(�J�ѻ���~��R�������x�����7 �����w������S4������#�}Y\�Ȕ�Mu�E���}�F#���)X����p�\�(�-a�ȴi��`0@�ۑ�0n��^��^�7aS��T/�z�� �̑�������nW�8A3��lN�eV8����K[�i`3-{܌��L�f��Xtvv�H$�l6�R�$,4��z�.�Kk(;��>}�R��l6���%lnn"�L�i8bmmMJ��K�%I�"ciL��n���*������cܿ?��NNN�����G�Ν;���F(��W�k�(�����{|���H$������ϴ�A�c�M�Ԧ�gF�o�E�꺊�k�1E���/�˅z�.,|�VC4��]���p�l��]��DH���tJ9�`���:7�s�L/�M��\����f��̭��, F� �ArJ�̞�&j}u�X������
����&Y�վR�T/�ɠ\.�x�h�TM�do�岄E��$�%Sxb�ȴꆰi�|���YL�4�����4J���.za��h�<�,�Z�T��cs���ݛ�fC��@2�����u��oX�W�������ݳ�3t:�� ׵$��F�^�#��>�dF�|�rf�ѐa4ŕ+Wdc3����b��t�W*�	c75�~@:R�XU��,�N}���c����Y:.���1�T/�Z���)�r�;f�X�p5sk�%5.�F�����qv�]��ud2���"�H ���5��[YY&�o��A�RA.��f�b��r��J����mlll��i-u1J��x<�o���|�<x���=�|>\�r��n߾����qb�bA���tS�q��}���Ń����yցY�
f����Ct��L#a��v;�.'lvۄ?0�z����\d�i�V�T���%�97����"�ֆ\j��R'>kF7���jO[&���~�|>�\�;mG�%/��e-��3����T*�j�"��t:�7��+|�К���h�v�(
B��	�uJ7_�m���S�IU��]�?�3�=��)L����ۜpؔ��dP���
��DP.��h4�$5��f��t���ד'OvR���x<�r�,��N�� �^�K[�Tq�[�^�χ���W�iG*c}}�V�BAJ���d�u�dp	�T�U�|�o	<u=A�e4�c���ߛc5���<�	+2�����������h4�'k�eѦ�~�ۛ(W�;u���$�������p2���׮]��瓆A�p�A���
���A8f�V��ɓ'R
___����_��� JӢ�N�"���boutt�����o����۷��_��n����
�\K��Ւ�Ѯ��8>>ƃ����B� �Y��yK��뮛մ�-��3/VaR���p8[;��n��Y�[j]�W(��쥓�x�l�ԛ%�e��Q/����Z���P�V%��Ϝ�\p����L�N/�2�_�L�%5:��Inh�ͦl�����x�ZE.�C x����W�X�=;;��\.�T*�	�D�#�s���P.�'$k�Y��[�`l6K�4�s�5�-���p�!��dLK��@u�\�t:H$8==E$A0���2r����Lt�Nm4��r��.��_�dr7��}^,w��4 �B��	YY.�6�m�f%7    IDAT�� �M�{���� �n�t�@�j�
���Y3˕�m�!�����,��dr�	ln:�@/��}9���e�e��>qOЩ[�e�l��.Yt����th�Z���[�hK�i�Y���ylz��j��H$p||���~�h �G@	����B8�[o�%��t�b�R	�T
�b'''(�ˢ�f���*��������Ǜ�0�j�P)W�6�P(�����)��$�v;~����ڵk�s�~��_�����f�A���ŏ
7Ul*{��	������d������,�eq�� !�)��z����(Ǎ��|����,ǰ&(Y(�p8҈E�T��a5_���a�d��e�!7@zSF7�2����s�f��ݗ�Z��s�f�MJ���Eb8"�� ��:�7�ϫ�~Z.�w�Y��'�o}>�� ���P.�Q(P.�%��8���A�&!�e���yY]3^�"y��U]�W��k暰�o,es�%�)�J���X[[����ꪀN�N����t:w�ᇯ�ܹ�f���W�\��P(���q�z=)�k�N��ʽ��m�fNt	]��$16��J%T�U����n�c}}]`����	��%0���,����d�ߋ�)5���%����^��Hd�]��m�43F����@@��MD���p4�0���f]ʞ&����2���V�$1�n����y}p9]����0�T:6$ݹs���Fs����pxx�D"�\.�r��T*%	o�hTt��PHbtFP*�P,����[�����&�{�=|���z�*���p��U��~���*�n�\O�>���2������㼚=�9R[�i.ǝ����%z��fV�56(��3���4����n�S���t.�C,C,�\���c,��� k��n��9��y��gƊ�����C�	Yi#�mf��9�RVr ��z��t��a���&�����_���䤗H$P,1�Ģ����� ���N�\F:�F���;m3�H��u����,�tQ�nd��@�}�/��hqk0��/z�	�0�D��(j��R������������
����ؚ7��K|�$�ɻ���(�J"Хbݜ2m,�g2�,5Q�����k\Ju���d28>>F�R�{ｇ��MY�YzՖ^}���&J��< ���qJ�f�X6������k����z�f�)>�d"�@�n�=�?#�ԍOf v�&ۨ�Ջ��o�
��y����T*!�I�](K ������mIkK&���bF�H��ea�s�����i���Z.��^]�r��>��c����E,��}n X�֍*��do���Ų����^�K���{��*c�akb��=.�`��`�ڤ!�U��$�նYZ���%v��XL��ds� ,V�ij�>wꔛP��݌:����O���lp"֩����5cS(��f4>�\{*�
�"�Ȯ��{��\����vR�ԧ�D�fS����gz��j�&�L6#�E��y����!	gI����|�՟i��y(��:�2@�yo���!��-�����	��M�,����� W�^E8���z��񸔇].z��z��������������ض���ɓ'��l��T*��L&1��G[+i��S�t�l&=��n��\��m�=gq��.R�NOOa�X�h4d1�V���Ljpi�m�Ya�d���e)^���p8��Β)֌.cE�kK�L�"S��<�\��.�5�vv�n��@�i�g4�g9���m�H5�/4��uҿ�F�R����c<~�.����b�ft�`f<�G0;�H$���<~�'''b�φ�j�:����Ȫ�nmm�����;��o����w�y�����nL�&��7�H�����`ۗIB=µU7>dh�x��vQ�TP�V���˸A�Da4|�Mm�LHg�<�k��ñ�sZ�)����d2��bX__ǻ�;>&�}b܈�b,��:����j5d�Y�䦍�n�5(���6d�@YY�ZMY��-��Ī�1|�5k�t:Q��ptt��z��Ç_����o@�K���曝l6{/�N�$��	\�q�� �2�H$$F��v���~�j�y�YXl���<n	F0;������h6�}�l����N�n[�{m���y<�{/�ʉ��J����~�:������-��ё`��:��@ p����ݾ}�Ƚ�V�}�N�w?~�J�"	'w��\i�&�6�Q�Jy���b�;`�X1�3 6�a�oll�f�!�J!�ϣ�h��rayy�XL\	�^�4x�j5�Ѣ�Ok^9�t��k�[�p	b�^�,�5|�9�|>a5��@�F=Y @�Z��Vhc�F�1�Y�]p9]�ƛ�R��r�,?7	���Ƞͫ�iq�Q�d���*>|(��o~�\�~������9�����ի⧻���\.�t:�T*%�Q�z�J�z]��x�G6:�`>�7n��/~�ܸq�:� �:i)K��G*�������O�?~<��m��z��ʡ_��p��p8��t'�b�鴄'D�Q����f�X �1����;���3�Y�rn��wZ��f������~{���X��h,W2�	�Z�^��f��\.�L&#�n&	�u�����x�|>�l�#�M@ı���)�ce�V������'�s5������t:�`0�k���aq_�z��f�������}4�M��ay^t����8�x<���S
�0�<��ec�Y���t]�0�������y��������yLKO{Ub�i�30�4�eI��].����*<B��������������������>���7 ��������I��wS���C6��rEwEk;)݉L�`d
�HhF�b��f}���C�{c�Lݯ����A:�F�RA�Xb���4�H`w�É�j�������� A��lvӚ>�/>?�|ZlQ��j�併#�n��%��h�+��߇es]�����5fv}��
�	� +���=&�r�
��H��O�}�A��mmm��l"�� ��NHr��ժ�~���7ڶ]�zW�^�fE�W��d=	^��T����k���Hc㼅�e_�p��Oͧ�8��K�G�Z�4O�%�ό��z�:����,A+e��M˒�U�����gn�BF�A��x�s�we��>nj{������R������l�#8禅	ʤ4�b����L�r����3��y�����kkk��{����L&w���l6��H$�iF���z<�CT*��i$�I���ȗY��M,{��&������E#��*��1S�y��<���������־J��i�Y0=0�;;==���>VVV���!�r�h�-�j�p||��h�s�ƍ{����ݼy��]�H$v����Q���t��$�����h]��@ʃ��!�\���x�v�E'9�`�s�*�\�f��r�,MF�����f�Z_�K�ZJ�ﱔ�L�� �x�BG͞n���.u�d���r#G=��b1�|n�_�Ր�d��'�P8��Zf��_)�4�C�j5��╕�62d�)	�5u8c���e�Cloo�`z]���F��Vxx=�Lܴ��OpK=t<Ǔ'O��������,8�����t���E}:�&�i;���%p�V+lV�TE4J�ɍ�^�tPA�����>ϼά���d��f��j���R�#��T�V�%ϗN��~����g�XV��כ~q�ʍ7�:߃15�� 9�N9�r��q.��x8�_ o �9�m�\���w=z�L&#�A�IX�r:��T*���8887�ca�T��+������4l� �WE�r��´�}։�B̯;�l��s�=�y`�<�����AQ#�f�����D���i�m�ِ�����CX�֝�ht��������xr�>|���d�e�ٝ�O�N4|uw.����q�׍)��革n83c��gdT���H���E�E��b��b��盰��z[�o����&K�l�ь��ln�	:���!퍸�j�ruJ�k����y1�H�1$T��	�ആ?�36mC;/�/^C>��Z'''�b�E����I`��T�Ò�8���	��F22��H�Ą�E�t���g�<�+������Cܿ_6�fs�IBf�Q&ft"�͒�zX0�h"J�s�gd��j��01���	��.u�L<�z��x<�V���e�����"� Z��x��\�
��80PO��&2j֩����N�Q׵ZM���j�A�k	#��ך׎�-Zو��M�<�w��Z��t8�P(�ɓ'�y���'O�|��;�Y{x���r�r/��|�������r�yRoL3�NNNprr"����<�_7�8+��<���آ��hy�.�����)OX��k�[dq���"�֊�6�N�ѣG����B����B������"<x  ;ׯ_�wpp��[o��f�������h��D����:J6`����&YGzT���lN�RF���b����T�`�G���bC ������.���lv�{��b��n�eE6�蝽q�ǟs�ꅐ��V�U��dY�椪�~F�'N�M�*0k��3�iuvv���S���	f���%�H�e2�׉�*v:��y<|�6�kkkX[[��ʊX|�ʇ��@� ���f��b}@�a�����0tI]��q�$	��}��)R����yO�E}.r���4svcs���i����͂�&/�����Y���ar�)~F_XYr�͆%׸I�s��"�n!�Vp#Lm���NNNpvv&��d��N�h�#�Ȅ����n��Vi[3�����뛵͘�����O3ה��j�0j��N���h��]��}��Ç�����o֞Y�Pح�j���#�Hi�C�Hz��2���	`?%���(f���A8ϡJ��fc3 l�;O�k&�GG�Np�KL�a�/:��7Y�7�̍6un4x��)������o#H|+ӌ���h�Zx��	�N���wrr��իW�L4�ד'Ovr�ܽ�������|KKK��@����(���w��MF�́@`��lJ�-.�n��}ҒK�v����P(H4���$�G����td�?�`8x�M�l��Ғ0Gto�s��eO2C<V|c@�f�	j���[����pvv6ᴠ�qV	|�󯁘��5{?�E�k�n�q||�V�%,\4���nݺ��W����іK7��}4�_�Һ>��qC�� 40�����XB2��X��J�ޜ���s��b�o�{�R=�-}ެ.d-���r������m6��qH�As��$�wuc!S<��0��:��4Er<�Y�:ZJM��4q||�R�$�����z]d	�
(<VIB�� F����DX�Q�D&^�	�զdEo(87h9�Q����m}��@�������������~��;w�Y{��O���Γ'O���&6�>�O~������ppp ->���$�*����N#fқ�iD�"�\筸�K1��X�ץ�8O>�yY�9v3��%���(����bXYY���A"��	� �VF�?�����x<����g�h��D�쵿����f�����(
�DA�F�Jv�}Q�٬8lnnʢD*����pb"84�S\.�l|�{Իj&cpY��N
�+V�'w��T�8�mY�gCA��# �o���jH�k�X��ܔ�Z���d��Ce��,��3:��>�06�h�j����H�Q�R�1
�����b�(����*�^����,6���C_'#�5J(��̩�f�x��~��G|���͚�36�̛��;/�[��͞���� �E�^˴�c �o�'J���]����םג�Em4�N��G���Y����899-	�y�[��4�1퐬��A����sg�17�#<��}n9V	FYQ`ŃcZ3�d͍N1D�k�-Ċ�"��;��Tn���Ç;�x����)NOO��v������F��L&���3$�I�J% �ͬ������[ӰԴ��y��E�E�sip�M��]�4V�eA��i�"�3���Ƭae�٬�3�6$���M���J�����X,�+W��������tz�Y`0�X,�����;�v�����g7n����h����{����^<�����S��dg�0Pg�fN@�z�l�xggg�l1����)%&z�R��E����f�/�~6�A�./��GkY�a��t#��`J�#�ߏ��e��zƋb�ו2��l��ɀ�R]v���g\䵅S�X�P�7~��l��i�.�Q7n���j2�?��H���d��y,��K�J��@�Q�df�N�a���d�J��L&�Ǐ����x���߿�r�,��y-I�����u7���e� ��m	������B���W����"�t|�x��R�M��a@K>��j�) i��z8���s�gs�ٔ���PO���4sˍ,-��á4�q�p80������ב%ݸIf�ǭ�6�mB���N�O�ۮ�9�F��ܩT
v�}��l~����/c��W�����6b�|~�X,~rrrr7����i�B�n�ý��㹐�	g��z_*����^��eL�������Y�E���g7�i�����I^�"�i�#ȝ�3+e��r���fQ���l�ƌ;�V����CI�y�wp��5iz)
�gd���[���k׮݋��moo�C��t:�q�V���������;�?�LyH����vUw
�\=::F(���x/�8�����Ό7{�4��5�,!j[���e)��Z-�j5���ŉ���S�Ap  �f�^W��Y���Ah-�bp/���5�\@{�1��K�f�drb"7F�Nca���\d"����Ş��� j����{a�Z��^����%D"�8h&�x~f�V��a���?�c�R����O�>ŷ�~������X'ȭ��Ml�g����g��Y=f��p8D����"��ce�iN���,�˨���ZR����$Do�Xm��z��gCU�V��&��+2d9#�ȄՓ�U�֒�#�}c&�m�X�����	�m�3�%�f^���]8�t_��n��j�9�cS���S��f�\��y5�MV�v�������B������?,�r||�S(>O��;H��2����G�t��Mj*����	ҩ��]�I�|�t�����0Т��y�u�ߞ�|����E���i�=�Ocm��6����F��ghVMw��N��h�J����=i>y��w���%%�l6+�w��v<�p8�i�Z����_�B����d2�/�Z���R)�6��C'�i}�����Rف�N����4Y(��fEB��ө�����&&&X&ʧ���M�p	� �"����r�V��^�O��z,�$ʅ����n��F�����&'Z�93s�}�Cv��� `�Z&ʠ4���'�E�^λ�?C9�E�]���f�����moo���!�buu�hTl��;��vQ��� �Qnh����������sp8R*�c�fS�5�^F��"���GO`n�X!�:VZm��A7�cLc3&��ͫ���	�����'�.������`����E&���b�>hV�\.�u��zc,RM!�כ ��ii��d�0��;�XH�̹�c�d]!�G��,��w���1v�������677��@����N�R��L&w>|�t:-�LKat�;���E4[M���9ֈm^7�]$��u������ ��M��.�k��4_��.I;�^v!%��]�dW�N���h�����alll��ի�y[��E���B��~��ju���� ������+W��]O4�\n�Z�~��{�}����|^��o��(E��ݙ`o-�����l6+� n@��4"���i ���/�y����ECO�\��⢪�׸S���[w����g���M?d�Y�d9�.]B�z\���E��~��|>�x<�L&#cYw��M賒_���x���NV��jaoo�@ �X�S���=m�R���,�i���H%S�7�R'�C#x��2�e��cV���]���{�N�� �z��_���Ύ���"h�9\}��b-K��ծ"�|���QϷ�����K7��d�¬xP��x�v�����J��~V92�SzޱZ���؞o���.��*ڝ�4�ROO�m�/Xy�v�/��z=��e�?;�������?�v��?����w����L&����c$��³*�R    IDAT8�z�y�DJ<G2���
#.����W�L_v¼�43)�$
�A�����(;���a����/�����̺9�.C�9qZ,�Z-�r9|��װZ���o���mܺu^�8==��5��j<@�P�͛7w"��������P諫W��ݱ��=��d2�W*��d2���3d�Yi���`՛�XQ��j������nWlr:���,�~?��0��,`L�a��a��-��{�5��t�k��N��_������[=n�g7\\x�dƸ�ӥ2��%��&}_%K���\(p||���ST*a��|S}���=�M{�y�1c2�/ޫR��l6�׋d2���S�A��~�>%G����4kOp�FBڕ%�I��|����7�z3����Y��S|��bҩ� ��}<�|>/!Jj����'��F�	�����h0a�Z�$Ϟ=��}��dkm6������m�w|�x�t*��|��$A���L�rn������c�:�ÁF"uK$�V�X^^ D"�	w��|.�,�9�ɭV����G���	�B����?~�������>z�h�P(|����^��1Lo�X-��ι��h�T*IRǷY�mF�9��I�����r_�D�uX��sq0;���@��㢾��4K}3k�ӌ'�Z�����	�q��loo�i&���j�����r9\�zu��������ɓ�������j�*������t:��-�f��Nr�%HI��(
����1��<\.�xV�F#�B!�|�X,�Z�a4� �q�q�=S���3��v;\N��gn�g�o�;~���8�k�A��j��f��f] ǒN����l�N�p���;�r]	�	"��������I��=�;�,�f��8/9gQ��=u� �7��n�c�-� ��'�������Y\� �K�<>64�2H�)¼jش�^�4�s.��b���x�ud�A�Ղ��E,C,;~8�?��a��l�5VI�<@p�O��=��1������O4:�(P��J�v9�T5H�&��)c-��MqRyq8a�Ye>c��m����Q.����&��{��A7���<o6����eZ[�x��Ͽ��/C��W׮]��"X���n���$�����r��?�H'�����Ғ�M���r9��y�r9����9dڳ�*�w_��v���"*�H	3p�(�>7��)5f]�E�$�y6�Aƅ��d��v�]��q���6cmm�`ׯ_��㑈I��d�����Vׯ_��z������ree�ov�I&�7�OR�T�����J���H$�N��Rhf9���%L^߳���4i�I.H�N�LfR3M� 4��jv��+��@+9��Nhs}�:���<�L�eE�$.�\P��9�����v�����d��Ɨn�+������i1���Ģ.)�6�����zFg=����}��8��1Z��{ad�u<����"�^���">��j�6.�|`�㯭��~�<��n�`K����>������%��r���Zr���ޜ�I��F�V���T���Z�3���$3�ٕ>�<�F�!���z]��R�`uuU6��t7 ��/.����@8�`0@.�C�XD8޵���f����ޗ�H�h4�7t=z���f?�V�;�d����f�b�� ���)e���4eZ�Z3���S��|�2	P�f��}�Dtޔ���H絉��gM��^6h�� ��L__v���~�Z-�������ڵk���F8F6�E�ѐɓ���
���:|>��{ｷ�p8��o5��\.�K���?�|�?���t"�!L��FN�>25<P��ħB� ���y�^T�U�J%ٙ��~aW��0�ɘ��m� ��R[l�LȮp�ݠ�����r4A#˨,�rl���:?~�ff��	��@3b,���}yM	8�s1��zRy�V1y����,�s�"a&7� �h	���n�ō޸�on�����"d�Ŝ7��aY�z7�q7kA�s�u�Y��MQ�L8�q���E�4Ƕ1�G���,�/��e6�钀�ZZ��6����1&�cԪ�j��>��N�����f7mZ������N{,i)����YךY����H����p8<a����5^+V���&�>}�@ ���vw[��݃��/�^�Wkkk�@���`'���K$;���h4�X,�F�Rm���}>�x'S"rrr�j�:��ϫJ���;����ȱ^��X���n��R^l�1��,���E��,W�i��9�YZeT��� �^�c_�[����Ν;XYY���G*9n2�Ұ�����ӻP(��l����?��۷o;VVV�XYY��N6'''��\���������ˏ��T����Ғ�!08C%�T�K���֫T*��� �'Ǣ{��]�T����n7��!�+���&XP�s%[�nm�[�Ǚ�F7�X`�E�X�%�%���q���"0�J���p�f���,Ĩi�."8Ak��������X���y�F#azM�ё�Uf��<��,p;�� ��Me+l&]�`�od�fʋ.b�l������mt��s��&�r�J�ժ I2��C��Y�Ǥ���3�����D3q$8�P{Jk@�]	p�y|O~_�Mm�E @�t��h8�p4��R�y�h�[�f�8::���	���H�4[MiV�ݖ��v��h4*�
�*��YGB3FK�J�&L��.r�`0��Fw�n�ݽ��/���W�X�o�����>}���?��Ow������ y���b������P(�^��R����3����\n"�o�eߴg�,�pъ�y�Es .JJN#f����.�h��a����H�΢'�'�y���l����5��Wv(
����|��c�M�\K.���.X�$0��d�L&�w�^����k��?���_,//;\.�?k�����J��i:��|Z�Tv3�Q�դ�9�A<��tOp8̉���v�Babҩ���0F}e�כ`ƴd�P���f�a8N�B1�F@��y|��\:�0�h��^�i����& W�	��u���q��z�`e;#:\���e�Rۑi�c�5��f}�}�h4�aHǋꦟE�=�J������'^}]	R�-�1�W͒��eI���{�Y��xL#6f� �k1˪�cD�^q<h����fS��`��5A3��\� `d�y,�����g�ZJ}���{���WG�j��g�(�f��m���p:�ye�h4B.����?~�\.'�z�XKc�[�7�l���b��G���`�T*�N��χH$2��P�T0��6�H$�Ǳ���`��n���������,--���n�T������ѣO�����Ǐe�|�{5螱���H$�n�+�o����������v�H��TS�.�t�穐M��(f:O��E�wSw�I� pc0�ս��y��.��L�5�K6�]Ŝpk��>}
�ӉV������NV60�M \^^��jE�RA�V���>��"VVVv���n�Ղ������_�A����"���Ig�\.�����j�R)�r9�R)Ir�Ւ����pK���"�lP������=_�Z��ٙ9�j5Y�4;��������t:�n�q��lmmI�M��\N�0Iڂ�c�7:,�QC�b��n������G6�I���?��|��ZJ�}�c�OwU�͒e�`��Ē�>�d�t��Q�����,�t���<+�E��.,eM�C ̓a,b�3��`h}Yɖn�2:h-�B1D6AQK��S�t�����̌���C ����}�4I�Z��k�Z3�zi\�(����]�xv�@p�]�ݮ�j�-���#�'/�R�$�?�`x~����ðZ�(�JH&��f����ƻﾋ��M�b1�j5
y/����#��j�`p7��\��_�����;w���@7�L����OS�T�������&	d�Y��e�@@�������
�ÈF���|h�Z8;;���=z�ǏK����r����c�e��N�K�U�_�u2�<�vZY�e>���̨w�l�<H���"�f��N0��	��Yy�y>��_��W��y\�z���X^^���G4E��G�ZE>�[�ݎ`0(�l��Q�������n,��B������_�A�3Ss��b��2JJ�tz���~�h4��l4ý��O[���Y��d
�|�z]�9m�4�e�Pr㟥��(
���p��X[[�P�J��D"!�P(��h7�P��5�KKK��{}����h4���u8T*�q�l���9a�#;j;���z�0^cg����h=�hX�%(h�Z¼0U��r	s��ò*��) �k�iƗ����MA������ό�%[��F.�.K[�2��,��<�Ĭ�y�z7���f�9� O��i9��:�L/�4܄�A����$H����5��$Z�*���Ɂl.ϝ�l��R���F �+Qd����x"�@.�C6���v�1\���IFSs���r,�\�=����������ocyy���d{{{�f��V���FIX*�B"�����n4�u�\w���?|�KKK��|6���ūnLK�ӻ�^��j��K&��6��]��r9�\P��
�N�c��rd�X�`�V�D�=£G�ptt$����D��-��T����/2_�s�e�0�,	�,�����v_�����l'.����o��]��ܸ���B��B����-��W�����ho3�NOO����p 
M4�	'�LJ�%��.//��s������6���lR����/f����~���`0��y�R�����6�m�V��\)��h�^�KJ���%C����R���򖖖��vxx�d2	�͆��5au��"��U�E��5+9)�f�V��R��FG�(
�~����Z-V�cY��A3�M��@�j�b8s����P|juÓ�'��)��-�R<>Yar�ϥ\�].�D��%36��N�Z�z|�����*�Vmy��E�nQ�����g��4��e�$� �U�.��nO�=k�h�1�5�3J9�ϩ�,s�K���1���ϒ<����W��,q3����P�pQB�gD7��&U�.x<��>�~q������Ba,�2�L���*���3<�"�PH�c�&R1q��i�][[���i��v;�\K�sS�J�`��w�n�n�р�����n�����~���t:��u��K��|>��j�>��j�r��|>?|����v�}�T*	�B}��?����sC�ڒ\����ڞ����lNXzN��������r
f�U��|����,
��Y�i|0\t�h��Uިi�?�F��:;W��������bXYY���6��ְ���H$"6Z�4iN�E�pbs�����H$���=�����������鴊�F�N�3��o>�z���� �b�|^��Z�RI�us���	U�X�|���|���.Ճ�	ep8H�R�f����wn�P���B(��ƌ4�\�tg{��B*��ӧO�D$�rumN��l�bQ�WK�a�FX�����hV�u��0�
�j���$�$<2d���e����k���kZ�L��4S�x�Lk�X,X[[Í7����P($�(�T
�R�HR3�ilpZt^Z�P|�
�"幋��۬f�E��<�ǯ��!`X^^���h�9i#�l6��5����a�z]����G}��fG�k������f4�L{3���<�7|�9�r �g0�9�3�|>8�J%����V��u5tޚ�-�x=(����F��|������j��L&�?��R�}���!��ۈ�b��7���N��r��L&#:�g��z�v����� `e���4Mۘr�R�ׇ�=���u�岬���n���}>�n�}L9���2�Ѩثu:������O�<�g�r��f��,fz�`��U��?�M�1����������[D}����U��Q�:3�,!�"l��×����w�	� ��˸v�"�����\X�#�p8�V*�	��B��r��ݎ���	V���u8�"zB���899�R��P�(R�2>��`P�m��%Yl.@�wm4(���f�R�b��jE�Z������4R��ժ��S�f����������c&���1�q��-�b1��~Yh-
��4n酔c�f��
+�,,V�#�sp�ƌ.5��D'�E�8�i��VT�C#�d����tP�VD�Ɔ�vt:�J%��q�\�[8�ᗿ�%�ܹ���m�A��i���y ���0fM�f6Y�:�͞q}]Ѫ^&�]Ċ�v=?�W�>�|n���۸}�6����3������V����(���ddW9�0�x8���j�v�02�r|V��W�x��D�sh6����E��b��f�6�$j�==gX2(��;%���L )2�f��h)7������"�N��l�<���&��D"!֔������D(B(B,�dCjs	vy��АխV���벮���]�˵k㳪;�j�n�Q��'�(�X,"{�vu<�;�����ʊ��~�/����@�F�~s�r���i��i�$�"��9�,��}�A1��N��y�o[���@�5�^�4z3jsm�=͇����Ա2�����7obss��px�ñV�I�����߳�jMd�s"�V�bc�+�(���%��قE���/`ܙJ�&mx��L��Ц�;qj��鴤HQ��Ő�,�qA�Z���Ӭ�q1�ys���	쎎��lm��F��۷ockk���21��eY�uZ��B�R�h�\�G�G��T���Xqa��ha�L�~�!���T*h4	m\�8��$��8�����"���w����{��m�����N@K�angm��Y�M����r_V����Y��m�����u��b����b{{��>��D"�ȎF���3�z��j��H$"��6^�o�fN7X��#jPu����c�(a`S�Y�7�Դk;2�jF`��[2� P��P.��H$���S��q���$4�[��>��z]�U�<��l6��fQ�Tpzz���-ܼy7o����"����~i6�ڦ�Ǎ��`0�F]����lQ{��Uۥ�@�}`�l��  a�Y$	@	��fb��� O�<���)�:��̥��cJ��3�2�Y9�|�~�o�e?��7���ˎ�L}�Y�rP����dp�/Y<���i#��tii	�J{{{���x��)�z�-�����v���0�D\�<�I�j�����r��l��l�V�aiiI .K6��Y���B���N�D�ÈN���B�V{OX�FP��dP*�$�4��r�$�T*���VOr��5��j-�q��h�\�\�ÇeR�ױ��*f(�F�Z���6>�?z�?��hg�$���&1<Os2��ة�-���ܒu��h.��t��Ǣ	��������O���>���۲�Y^^�[o��l6�Z�&���Lc1���L����/"}�5��-lz|Oc�5�2�f�'�p5m��1vF�^��3�sӕ�!�m�Zp�݈F�x��p��\�vM�u���z�*���i��H��k9߰�T�V�l6�h4
��e3�1m^1&��@`��ǣ��uS�NP4V4�m鏥X�_q��Z�������&����8::��t�.n�m��l����{Y�Vqpp�|>�r��r����-loo#���v#����Ą�I3?x��z<�	��Ԩ�=tb%ߓcAGa����j�F�h+++�����M{&�����N�e�auT��"�ݴޟE6��\��HC^�E��5 ��?'�����y��� g��1nӺe��O�2�a5���,��%� P(
�4�������իX[[�K[1N��8�>|�/����	�uX�fp)��r5������E�E��?�z8C�V�l�d2)�L[^^{.v�	C/�F�X�4{ ٵm����̐�fC�^����qrr���3ܺu���b#%�Q?xВ6`�x=	�B��Q6���,6����c�=ϗ�l\4����r�b�E��F��q�~��࣏>��֖�v��!�^/�z�-a��Y���V�LӨ}S5��&�0V��i�͚?ϛ�c�hh�~���8�z/�����hK-�#�c\���q������xL�|�������[�y�&����t:�h4���D~��|PZ    IDAT���e�r��M�q��Xh���M��Mo(B4E8F �p�S|���L $�ac�t/7�WZ���ʊ��Z�D?��R�$�%�@>_�l���8<<�����H��jpx�q�G���̼n�冾\.����H�R��x뭷������U����;�Z���u��y�fF8����"^o3�5+ύ����3f�M�L���rH$"�c�%%q�fa>�\J�I�*z�����1ZT�z���Kap�i0fE?^�ԿHR�e��&��vQ�����E��$�N�&�p8<ѩ~xx�F����c\�v[[[Ҹ�sч�!J���}��%��9I�4ӧ��u\��66[�9yr�dY��H�V�A:�F2��]4�g)ŠΘ,��:]�!�ev�~]����y���F-��#	���6N�zSA&]7ԐY��q��\�d.�uo�,��N	<�L;&�t:�t:�R�$]�d�l6nܸ�_���x�����	��-`�n����5C!NOO����4k<r�ݦ�M.�ӧE��k@k���bcd���e:֨�,�f�$3��C���PJC#U���d-�|�G���6W�c6J,"��~?~��_�Ν;�D"��l6�,--	��è�j��f��j��d	�@�X�`p"\��[��d5��jI�+��|YQ�x]g�"�םNg��R��܌PF���̘���C���#�N�P(ȳ��e��c��r�$g[��:���b%�Yz�T�������M����&$
��x��z��忻ݮ�5�|��sC������Fb��&j�N��I��z�lVȣT*%8}�F�bpy����$�$
����~�i�eT��Ӓ$�];����l�En�e&�]���l�}�����7P7!h#~��&ZU��dR��GGG�B���l��X̼y�b��B2��;W��Nqb7�s����rx�XD�ٔ��e�r�,��nzBr�"�"��]���>A��V��z<G�XD:����)VVV���*̺n�����O�ݑ���^_����a�B�+m�t�������׌���/��3�2�R�2��t��|�S����	�Ϗ�`̒Q�Fm���:>����v1�?==fˌ��Za���z���Z=m0�����L���禀�#�Ӷ��>��xhg3-1�������~�]��JE���������č1�ǐ�U��@ �p8���5�������=��}��a�l�������x��B!�r����4�f�C��@ ���M��d�co�Z(��2�ȧ�X��j5��t|���v�-�T������^����J����? ��x��P��O�boo����0��񚛹n,*ۛ׀f���L+�[o��Ƽ^���,�����T��h4:��&дZ��B}!�O�{��9�Nج6�;m�;�W���l�86������8::B"��Ϊa>�G�T���	����:M*4+N�e��Ecv��,Ƚ�^��}��~��D�i7o���,&׌�6�5qBc�,��!|��kJ��O@��4w	������ԹP3a���MX�pa��]�3�B�bJ�o�Ơ�5x\����YW�e�K4�':���*@Sv�\.�H$"e�P(�� R�m�c��#�;��v`���`�ȝ ��8'�h��8~�iН�����/��Hr��Z.���eL�ՊA��?�ʕ+�X������5��uӅ��FG])��F*�7+P�a��?���b56�=G͘7^#ld�	��Xr��0Y\zwNǴ�3�%��E0F�S��'��z�X]]ŕ+Wp��uܼyS 8Ǟ�4Z����ړ�eh~F��A�X�D�w��461Q���n��;�HV�V'��hō��%ƽ�Ac������u����{�S�L&���S<|��ZM*[|N���h{3��8�.�&�r\h��1��r�,�@ �P($޹kkk�����ʊ�F��k
u��Ǻ��{BI���k��M$��R��q�\�����ӧT��lSV�7��i��y�i}<?��r{^�{Y��~�������� ���guE'"���;I5�2'�	�R��XHj�h�OM��1��n��f��j{䌞��p�}U��g�Z�,�؈E�Y{ƒY2�]j��c�����f��y;t��K�64>o6�2�3�n}}ׯ_����l8x]Y�g��Q�k�8ӛ �t@�G�-d\�=s��p8^��%���{�帮3Kt!�<	� 8��eѲ-W�����Q���RO����~�~��PT�o(�U�-�f��@ �!��9�������{�}�t5"�0d�<gk�o}k�Z-_I���O&�c���C˵k�((��j\J��d=��ylll�'?�	��R2HR�!��-M����u(���'\C�p	�m DZR�q�n%��?Z��HݶtD��t�]p�i���͜��>�,�J&�:�f�������K A������0�?\�M��'�	Z���!Z�NOO� ��!���ń��@I�,�9�`zqs>�Z::���qJY�pX��#��g+�����!1���V6y�@r�I{.�F����P(�`�'O�`{{[Hh5V����땴l$��=�)�LrK�RK1�!H����������x��)������3t:u���!A�(�,�L�u�ܨ~�>���ep�Z��"A�5��9�u���t�d��� ����̲�����@�����8�/7Yz�f�Hg�K,�I����v�?f�_tW�m�v�JNA���t��K6��%˥2%F_�_�ge{}�g�}�uw�]��i���n�qzz���-�,���2Yj	��*0���಩EO0�%~�l#=i�;;::R�Ȓ�z�5��x<�?���S&�����b�Y���B�����W���,�����P&�>]2��џ�d�M��%~鄡��Jp+��KW*��n�gcue4ǚ���H�!A����������/����C,�CJ�z��߿����
������zV�ݗ���P6\qm8;;C:�V��h4P.���B�Y�\�dQW���㜦�e�Gy|Oj؏������n/Yh�@(�S�o}>�]����J�:�{&�x<�ӧO��鋄ɍ����(=6K��R剄��Ņ����������\{OOO�|b��F��p]��S�f��+^<�j�I� �2����A�g>@9�:�jT�
_HB"�Ɔ������� 7���F�h���],�X�w�ݮ9�v�i2jb(IZ�-?�,!I[��d��h��p����&��K�|/���,�l�pM��:SG�Ϙ���%�.��Z���1z��?�F��F��" ��*���3��/�2PC�d=�����|>WL���prr��к5�\��}"ؙL&���0ճ�������xd�_v3ֳV��L�dtd���t���\�ܒ����dHu0!\���ּ���9�e��61��T*)_Z]_��(�:�~X6����}���5�3�S<x�?���n�k�O���ÒU&���3���n�\.�C+&<@�`/�+$��"�á��P��
��$�����{����j����s���*P���uVډ���
"	�Egf?��Y���r:���ӱ�]}I��:y�R.�����n��N��dW��E�Y�dO�z_��EOB'��~�=��w�t��Q�����º�+3a�<(�!J�d\WHa��6���>��9!}>�>���_��O��S%���U�`E��.{ڵ�z����)�t[,]��� �@`'����F-�)�� �A�A�X_`| �|�kC嵍F#e{F�;���������@���&���B��d���yS���V����c�fꏞ�dby��޺���믿Vmx���+��O��H��HgDS����3t�4���V�,�d�L��Ɇ�,E�=�u��D���s���#	�s����P�\�z�*��$yx���l��k��.����a��N����/��g�}���3L�ӥC�O���P!��ʔ,i%}i)�`S,K߲�)�ϫ5u:�*�B��Ucr��� K6�u:�<�q"��/��ֺ ���MJae_��B�����N�*��r��H����;����e�&���O��k��%@gɃt�a���Aq�AV�.y���i���9_�֤�Ҍ^�����ut�(_�5����7*��(��]����w��=�W��dF��S�/mr���)�d���t+}e%��k&��'�n�d[x�,AR����P�PK�.��k<>>F:�ƃ�'#�uj�)/��i�+��,1��:�V��1Y]��M5��W~�>��j���?�b�������?�\~i~�q�S���妈��x�զr*7C�.$5��b ]I�����f�)�_z���o)M��Q:��AP�kYv71���"�y}N��k	�Y.���>(��M�0���ɇ� ��c᫯�������MY�b4m�zP�����J�+�����JC�PP���9�A9�dD�\� r�I`�%kT)��q��'�ε�)�B��! �\�_�d&g��� �CV Lv~�ݛKk�`bOM{�e5�Ő����k���K�^��'�u�հ,�$���i���.K mڴ}t�&���n�kUe���;��g�锠Y��I+'�Ӵ{Si��z�����#��������W��J�t��Z�|�t����L�� [+7X=�C��U�l��d�>�>?�D4�����?�\xܼy��.S��t1}E� d����d�L+�Q�X>� ���|H���h�;^g���	��-��|�3���.���Y��������e)�8==��Ǐ��?��j)�L����6��D��/��)��%tӽࡍ�3<��*���J�/~V	���Z�H[U˧�Ǵwؘ`�.Ӈ�3�ť��*L���5��~��m}5Q���1�z���E��H��V�/�˦/�Q��!�����A�m�4�V�@lܶ���`�E�Ƶ@��	ai�H�J���b�S۹�ü�.>Պ8�T>S���#-eiR2��L���ҽ�$�/i�d
p L1�t��x�������*��*677����}$x0�~�_�y�K��Z�;L�G2���sH���@U�eD�K�ۚɤ-�j�61�d&������{�.��'�<Yk�����c>��Ǐq~~����g���[*�N"�X�C<���>o=��%��_[Z	#!��SәKR�O�$���jоk���YW�ۖ�Ė�����	wa�]��5}d$>.A�$�I0�a�f�A�� Ip�6Z��2ή���pH�(_��S&���T�
a�&��\ �u�쓞�ecML�:��b����a���}'hR>}>���`�ϒZB2F�2�U���Ԉ��釜�{��(K��`0�Ç���T�t�TB�TZbT�����a��3�u��UjL����-RB*)y�c_���`'-�t?�_�-js�ӤK�����=C2�����P? �6�w�y=YL69�J,��E @����������(�JƘհeO��[*�@�߷E:s��&N�$b�����ּ�Î��Ԃ��k.�U�:5�x)E��3X}�*|%����2�NÀ�(vc��"�5N�0��>c9r�YX4��l}���ʪ>7=jw�kA�Eٙ�Չ���̙i��2�}Ne&���m��A�� �Qv̿�^��������Y��o��ִ�D)J���6�=z�_~�%ʥ2nܸ�L6��\#5�&�y͓�DE:3�X,*��N���%M�U,Q�T�f��d�j������0����ėM|��^�&�ˆ#j�u����ej�d���R��r��"E�A�6^�����x]�i����c���u�2#��̭|�t*X,h�Z������1�� :���W�g��&�Ao�sz4��*؀�m�0ݫ�{��؇I�2��.�3���6�Tl�ܗ��\&Y�.��\.2��찬$�/��颼,qt��(ua��e���@#�����lz<׽����Ԧ(�]��D�s�L��A�9jp�e�m]+�Y� nT �sz��	�������S��s�2�����@jf)�x��	��?U���z]�0P��b�Z�z�F�tZ�1يN����=H"�J���R����i�둠��{����6t����v��;�nn)��N���K]�1e��|>Wͅ�L����z��r�l&X�������n���3���K|���8<<\�v&Д�]>�\�S��y��H�}уzL �uPw����m`>�r`�!�̵0L�3���.>c�ww�.<	�6L���'�5*���9��:�^�cMb3d�
�}Ra�t�IL�0 �V
:���!�6	��B�L�_�m. 4����yV��u�n}�\�<_@���[l�!�L[4���Z-<}�?�������իK�n�b(��3�f3C���>��3t�]��J�<;;�d2A�X���&666�h4�X,p||���ct: @��@�R���6j����<::³g��e����� �^O��i�F��i[�VK��$9�p�Z�~�t�b���T*�����n+M(����:��n��<n�$�Z����j
ܾ}�^o�QAgS�T+���A����ٳg����_|�/���?F��U~���5�6�L�cPS�O)ֵ�R�lG�I���.9��WAw�qU�¬.��Y˸�S��/rF0�	C\]&s��Z�����;����fl@�vb��%n���6��"�\]F���"�GGv���0�O�.}\R��S�Oi)�4mc�}���,ޮ$����*uC21),�4N`J���_~�%NOO��t���ڵk���_�i���SiK/�R���6)	�[K�r���*P��n��T*�v��R��"E��)�á�,&hi�Z*���T��L�#���f
t�q��b�L�w�u�?���ɺ����Q��bQ%7ɦِH��x<Vv�^�l6C�P��[���,�~��1��Q,���T�������ѣG�������#�+C|ktp�&gS�Ճ��&�J��0� '���+�?�˰���?��?|� ��F4��_ȵ9[�h�}� |��d~6��v����3vU"2�2��ܺ�=,�~Y̭������  �$��|�bQ��$�J������������[Ae���O�M8ʩ=�w�m�2Z��M}�`0��������E&WA��82� �����w��Ϥq��}<}�T���k��0�NU��ܥ^t6���T}��u�ݮQ�(�&��b���7ЍF#��Qj������v�@��{qq�$����5�N��t�k��G:��������'���'9�`��t:�V��{������=�����=����RB�ll� ��EA~�q+@A.>]�>�z��i�tŝ�>��[�I��~Ea��ȶ|�_q��A!.g�8�:l]��=��2�^h�B��b�F��`Ee]%�5W���-�������:�^�\W�D����hs�b���ʨ%���A�*�X6�ո2� 	���Q�n�z=���V��/�Kܹs�Ba���T2K�Ө��x�����<��h����8<< ¤�?c��I�XjB�bl�j�����AQ�A..��v�QP���R�R6�
����^���;��ӟ��n�B�RYJz�a��\y,ӣy2������=>��3��O�����j��\��=��u�4���ƇQ
3ףV���.{k��&[>��=J�d�!�d�&�t�[�Ƨ2�Z�m��N:i"0qU���q��_(�����0�b�SQQ�`F]L�N���f�b;��$�]v'�m6-���,��U��1D��	HĹ�I.|� �l�l{�R��eb�'O��a:���{
�-4�v��y���e�y%�H���������ﯮ��"�0�^�b˥3�-����jH0dk���e�����4���,���p��\ٺ�ݫ��s�nܸ� ��E��Lq�N������/��?�_|������v�L�T*-���l�|�[��e*aA����`�f>��Cț�z���@{�Tr}�-�}����o}{T�6�����3&�k;��E\@m+�G�烒P�_A�m�&QRݖIl�I:a.W    IDAT�.�SF�'�%�v�f����7W<�S<���)t�P2������888P j4�bf�B�Kz�D�E���b�X�R��ʕ+�u�Z��?�V��^��"��W�ϔL��5��i�m����T�2��ߋ���@q���Q�V�ass7n�P�v[[[������:666P�VU�������f����n��Ç����?��Ox��f���b�	�Mi_A$�>~�ؠ�:��i��[!��]��k��='�!=�1�ϻ m봸��F<�I��u�mG��uO�k�6���޸aX[��ֻx��A�i��uN,����fA�N�Z�M���z׳���5�A�L�R	��������o��v�X,0�q��m4�M��y�����r�����2vvv���*��'O������<}�T9+0@A���`�'Y�T��uޛ6a�ߛ^��xOd��x<���9��9�^���7o�w��ݻw����j��Z���(�`���Iw,W�1�������w�}�{��)��J��|>���|f����Ȗaz��e�������2 v��)L_M�8��+�ö_�Z�E^������V��@xYs(�{N�����bÚ4�\M�?������Y\�F�l�$����]�����w1�{�Fg���mI�9�ǎ&L�-
s�%CP��)cp���=??W���������Ɔ���F���zr���"��&������qvv���}ܿ���C���q���L$0�Lq=�O�O)�]�]�Q�aVw
�Ҳk2��{��尻���w���ݻ�s��ܹ���u�� �h�&�Ȕ��yp�k<==���>���k|���x��9��>J����Q��L��l&M�6��gc#��-.06��2��a.	��8�i��tͿ$�\k�i�$����>�\Q��|lEMխ������u�2a&��憵���>�RA��4�~/��Y�l')��2ʢ2�A��h] 4HV��8��7�"(��~�å�� ��3�����g�ْ�����j��>C��Q��?��Oq��5T*�$+(Ӻ�LV.��h4������]loo�^��R��R�`ooGGG�F���J�+��d��/�s߃Hl ����FB�K^&�]�r~�!~�_��>��Ύ�!�=�Ze�w&S&�|��)NOO���S<z�_�5<x�V��R�x����d>��f�Z_�\Z�(��I��6�0�LO��$]Z�˲�@�Mr�!�u0	
0��II7���$��qȘ�)I�2�. �kR����]6{[C����{��1�Q1��s�0�k�~��a���B�/f�x��(�1Uaz��KM�k��-���ٵ �nx&F8����_���I2��l�~������3<�������q��m�����9#p��&*��L&����t��u��������}��^�ѕ�#���yOLdb�OQy_�m��}�#C��`�����^��>� ��>�^��f��B��>����Rõ	c�iC���ܻw������-
��mx6�m���������m1¦C��r��	}6?�-�M���.&�25�A}��9'��d;�}�ПYl�̯ 0����w�.I�l��~Z	�a:��1�@�v��uP�;P|NdI�Ǩ 9L���fh}8W�PP�APef���Ҷ	�w��<�g���m�"�m��>�>��brV`P �5K@���S��m����������p��ܼy���J��&��l��d� �toݺ���5U����������4���~����/���3?�f�ޑ}���%K͟�f3�8W�T������]lmmacc�f7n��{ｇ��]�C+C)����ҫv8���GGG888��g�pvv���C%K�ǨV����h�ms�ƈ���T֒Xm@Nj�ma����{����U����Q�WP��oE)*�`�i��a��(�,j�\\F�u���d�����8��(шQ&��[25�>]��7�N�S�ۤ����m�~�(`�S�K���T4��t}�/���5��R����{.�C��@���x<�Ç�������[�n�����>�@5���dsߗ�hԐR�p��u��eܼy'''*������Ϟ=C������q~~�:��痂t�}���R#��E���ds���
:���1��2nܸ���]���;�}�6����������֔c�d2�h4ző��ft����>�7�|���:��:�F���[WN~_��Z�l:��\k]�j�A��EP�M�k��� �0�׽��&���Y��]����7$���`��=+�������s��~�����=S��q�~P��m��a������la�u���}V[i/	/Hߓm��('��@�:�,�o8� ԉN&<y��V���H����z������.j��h���
,JPI�;��Q�VQ�V����"o���>��?���=���?V�n:�.%���*Yn
d�)��?�7	d%�f�
ē��ƍx�wp���P�J%
՘G�p��u���???���>|��?������Ct�]L&�Ed2�E�Rn����7$���kv�*-Ki����Ȧ3������#us�\����Q%do��y���L_ i:tɃ��g�l�I��Y�}��$������\+��b0��q���O7�_˾�M-0a= }J�����T���a:J}�m��;�{@��[6��'��?���.�`b6����_}���ΰ����W�b{{�fS��Xƿ�N���z
h�=�P(�\.��<��իWq��u`kk[[[899A���d2A��S.���]��ґ���`���P((]�t���C6�E�P@�PP,t�XD�^����_���ׯckk�z]��|����F *�,��!�N�����St:��m�ѣG��ﰿ����K�J��
İ���/�i@M�_v���gҚ���&k7[i��]���R}/�B��6��4���Q��$0�mu�7��Ll���=+.���5v2>�8�~/����(k�%~�j��pkj�
�`�}�ݵ���c�T��|� �u��*SX�5���w8==E�XD�����:�_������x�w����F��@&���p (�����d�V�^���.��6��>��):g��N�g���
 KP�/��ԽRL=�����]%���C�Z��ښ
k�T*J21�LTH�<(d2h�=���9������<z����J�qzz���S�,5����K�0mv������p���{�����]ij>`6�F��5Ϥ��������#}�N�{,}�_WE��x���$Wrj�g�A�p_�`
���9	$f/���D��v�7y"���	0m���,v�n�gl��2_�nb��� �aբl|.�1����Z|���v:!���ɓ'x���y������;w��XC�\R/��t:�h4ZJ1���2���&���!��9F��J���P���x��d�� �N�n	p/..��dT�0���%��i�U*��{��Io���d����j	Ni����|���x�������N��z�Ţ: H9�,�ۘ?���S͉��l��#t>A����9��$�|������Q�R��G��C@�kA���:��da�"�2�q?�+���h�M.qYH���שk���|��4JaI�p��L�QI2�>�,��+.�`�o_���cj�q�������Yߓ��9��9�鴒�z=coo�V��Ǹs�nܸ�d|�r���9���/�_�xiF/�r���FɄV���x<~�:L\j`��V��%��Lf�=$@�.Y�~�fZ~-e�F�+��t:E�����1>|����_�5=z��ϟ�47:G
%� ����n�gҫ�m������O_oq9VM�BTg�Z.��t��֬0���$����I������I�k�`�.�����}f>� �%�"���3��g��2HI�x�L��e��}��t�e*�j���
u�F�.��9dӅ����sRt1.�6��*I�T����:�}B�1�T|�^>���R)���*��`�N��n���t�n��v��n����m˛N����RJAͪdv9n	Zs���J���v ���z���(��d�� s�,|�T*,��dF�JY�-��h4�h4B���������<x� _|��߿���$S,���#W�^4����a���
��l����+�ݥM��ܰ��(�c���bԣ��o
�I�� :c�@�ܛ(=�1���G.׌ c �������P���6�IFqNpqK)a_ߕ�e;y'%H���5�|On>a�%=^�ȸy�����0ZYW�X�7�5JTp���`cK]���5�.���3J9�WڂM&<x� �vGGGx��vvv����Z��Z����M��ud�Y��EpKvU����I��#�͆��z�� �������	�[�b����U�E��S�c�%ܿ���888�x<V�gtE�U���!�VO�r�s�
��j_�
�Lg_m���Q(�9����7EK�?�L��8��/�
:��d*a?�oS�τ�cw}^=�$l��)�1���,�-�;M�N.@�#�;�ðJ�	��N�F_�n��O��'�:��/7f��$�z�s\=N�j���I:�Ї)���E�X�k�����0bb��:qxx�^����h��h`mm�F7n��իW������e���+�,�ו�U��J�!`k1ن��%�%��iT�U�2�q=;;S��'''x���?���#�����n���Di���*����vuc��Aص<�9�l���:|4�Q5�a��d�*|Y�8QǾ��2Ӭ��GI0�q�i��������/����h��3Fn\K�(������8l@�������$�_nP��t
������O�F�E"�d�k�N6� '�	�JH�gd��(G�� 6+����I]*-������c
4�j5<|�;;;�v�nܸ�w�}����D.�9H���=�rJ�iP��$�1Y��g�[P�@��`0�Ç��_������8<<T���u�K3y�ڞ�-8�]1��l���e��
Z/l%k[E˖XŃ4i��7����oR��:�E�?I�DI�����s��s�͇98$!���Y&��pi����('}}r��A�{6�ܷTt@���b�����걅&V�%9�m>.�҃�6� ����g��I��������U��{`��8Rݜd1�#M��*���nc0��jaoo��q��M���ۊ��!�̭4e��LN��	�}68���53Jؼ��v��t���[|���v�899�h4R��Z���_�fiuD&W���"Imө7�m�I Aۡ4���R��TKM�^�w��[��+��ߴ���g������	�	����\�� Pi�6[���ʄ(��D��[A���.�$�N�>2���$Ր`��5m�oQ��qOw&O�0�6ʘsrc�"Ǵ>���l}:b}���1|�lE���k"����K��~x���ҡ޼y�n�+WP��Q.�_i#cJ_Z�r����jA�hR+/C-.f�����qq�ꃃ<x� �=��Ǐqpp�v��4�*0�X,b�X(0��)Y-�`b
Y���q��,���eP�$(����AH? �6���&w	#�&�3
�Z��X��C�����M�a���Q�}1c�I��ܷ�˥A�e����l�/�I?*ȍ
L��AQ�L��~Q%
A��M3m����l�|�6S|��LQ��Q~������0y�ں蓌�tUp䵦�i���M���t���S�F#�޽{�V��v��ͦj��,n�������e��$+*��� ����@i�iƿ�v����8==U!Ϟ=C��R,0���jeҚi=�.��C�&m����TM�RH�p$�ꠃ�m_����~��Q���ꐍ����M�2�+A^ۗa%�z�>AI�l��7a�j{Varl�#,{����v۠�L=jT�5�עm�ۺ[�hc}ɣ��MMEA�p_����b�l,b;���6� �G]��s�7����Y��δ��K����)�I�%�r]o���u|_�d	[���&z�����b����>��!����J���?�^�+�P( ��/1��rY}�X,��/2�:�:��0�L0�N����̿��x<F���h4�p8T�ǿ��z�t:�h�Z899A��R���f��639��� ッ6h��Z6�ʦ9���dg�yP���6"�A�K��j��!f:l��Ǿ��6�$�a����E0绷���o�u*i�Dӵo�i8Nn}}�]̸H����5}�g�3Cׂe��|H}E�.C��`�r؃�l���\#���lE�4Vl����mR�6��l�ǔeKn�&N��J�0��3`�6m ��Tߐu6H��-5��u��S�G����5F�2]߃8-Fex�t:���>�?�\Q+5� P(P(P*�P(��6f ������b��B��^w:���4��1&X��o{qq��u`�z^6�6x�9��G��5��Ɛ�;��{qq��!�<|� #5��똬;﷔�L&�Wҭt�FT�ذko�=ۗlr�o���q��|��0�hXG��	���w׽��� �)I�(���5͓��L�A�Dߗճ����A�ئ�����ak�	z�Q3�]�$jg�����f�A̱�5����]�]6�m15���l`L�<YZ'���� ߛ.7d�"�tmk�1F��\5=w���i.��@����Ai�|/�;���`��\��;�{����M��2mL2�|v6)=l�ϪK�y�6A`�X9�}˖6��@]r�yȃ���
��"��������|=�<�ϱ���1��FF�,� 9O�[�w��Y��>�Na�{�士Z��+�B������� �+)ip�C
ٞqP%�4.m��>�?a�6��3h|��I�G��*GՖ�&�ip�zJW#Eh�cCVba[/+ ����SF
��ĻJ#6=��雥l�&'u�I���K%���U`�(�� =!���R�9����#����ӴY�ȱ�7>�FA]�>�&�řO�#h3��A޶�������y���
��� �Rn`��: ���Y/��
M�l�~��=D�c����Ev]Z�J��$i�?C�\F�\V�v8�*���
��1��.���1��!Egwm�t&���򲿢����o��a��.��i�{�Vp�g0U�|H���Ʀ�IzpG�Q����BO���M�`�N�>v1oң0����J�Ib�
#���,_�r)Kʫ����].�Q�TP*�Ԇ�MYj<%@�-� ����������@5)����W�F�0!�_�=��9�Q`��&#�m.K0"B]���V�>'�z���b�����T�C$�t[�E�ȿ1~9�(A ��!�P(�Z�*W�L&��g:�Ƀh�XD.��t:����z���x�V����s�ML-5�^������V�^A���C?�pS�M���m8X\��u�#���A�h.p�u	��l�a��}r���ui��<��Z�0�~ҵ1e�a�b��0Ѹ�����]���/�&1��+� h�N��<�R���j4���V���j������]�jn��_�v��t�;�T*�X,b4a4)�+�����F�����Ņ�Lե8�a���D}؅9J��H�n��2EPG�nɆGeh��$��k��u綹lZ���V��t����(��7��jKr�J����uT9F�f���g��R)���r�T*(��(�����r��jK:��p��h�n��n��X]�������CIVi��n�$�����r�F����q���� i�:�k&�����[��z�R��i؇���X\�����v@	bK.�dir�^tU	dㆩ���kj~�m:(�~��W ��󊡕���%��|^o:�F&�RƐI��5u�&Vq�X�\.#��.i���;7�N��v��@n��E��{�:b~1W%Xn�.���t&�Ak��#���^Q�A�:�z�z?[\u�gk�anm�uqq��d�*2܃�,e�f�ZM�ۍF#��e����X,"�N����].�Q*�����>�[�X��(
JQ.��d
�nW���ڈ�    IDAT�r��t�@t�����mR��e.�9��y]͑oc�T�������0X/�������8Hx|��Ĝ� @�rN��{>�sI,>>��wP�6�(aI�:Qݧ �vۢ�S��?��X,P�V����f��z��R�� 9���䮮���~U��K00[,5������4P�����	������m��m�C����?�c2�(���dnM�ao�W���,ccR�|~�E&6����άF�L����j�)�̶^�*G>�WF.�J%T�U�H���TA6o�Z�q��x���pJ(%�������Œ��a#�R	�ZM�Ꝟ����6M��Y:����E��Zob�����!N������"s���� �a��	:EI���[��w}l�\��D&]����&����wtO����5��e�ir�������4F��J�P�T������{ׯ_G�����b����Β��,���^\ 3,5���h�+_ꁹ��H,��z=��}�j5lll������'''��z���KѿzY���pF	�Hbs
��O�U3%1��l]@�')2N���ێɯ���M�J��?q�P@�RA�^�������P�M&2�6!���NH�0�X)ᡓ�o�L��!zO&�%V�w3��ra�L&ꚺ�.:�2�F�Q�!�5~��6�t���v ����QI�0��\�f�kW�CC&�B�1	�\�4��e�\�g�״���)>'����0�+_)��M�=���\|�vؐe:��,h�g��:铙�f�����ׯ���۸}�6666TCu��	��I���JJ�b	z���������fs<��4�/2R�,4���R*�~��n��V��������������F���0�L6���ʑ-9�Um�1t�u�vhw��AQ�AU��1HAɑ6�X�{W@��Ԯ����V�)Y�%�.)?���K�J�1p�����G-��r�Q:ĹF��>n�+V�T��尶���B�v���J�@v���d�f������t
1�?�I��kD�U�|�X��^�g��U�l���'YU
z�a�KsQHb�=uD)��ޣa������Þ�l%�8���[������"2M 3h��mY��d������v�nݺ��ׯcss�RIm���������IV���E7x��T:�:����ʀ�sD�F4y�|^5ᰣ���B1a�|^9/�E+��t�da��g��-��Ut5��5��eM����d�L��46���u����®C6yx����~677�����d `I��Ûn��*��*��c5feń��@S�3��R�.�m��偘kF�\F�V���:NNN����N���0��t�J|������:I�$�Τ+@I���e�}@n�������j�uU�^�.f!H�����(�oX['����tM,���n�&�W�����������r�a�XZ�Q���Ƶkװ���Z��tzd��K+_�����Eb���'SK�u�2�b�@��C����ʊb_	��cr.{�`KMgܰ�jq�/�����f��j��j(
����t:�&�}�4-^>�a��1�[�
����h���>��Jݧ�/��u�X���F>�Ї�u�H9����"��&vww����r��w2dCj_�+�(���1yW��G����סd��o&�7�ɨ
��Z4�MT*d�Y�������N��D��u������AU=���@7ȱ�%�{nQ�����uApI� �|����v|�>s�UB�v\f잫��V�k�����F_����A��rM6<6-�-v6�3����T���kbu�A�F�H��|��\��&vvv�����W�bss�B�|^9Ю����8f������bL���f3e3D�����(P�r����/oz���.������[\6�
���P.�+EƘ� �����Y���;��n$6[:v3, z}��Q�w�˔����(*Ǚ�u��/���V9���tE`����:677Q��P*� ���,R������DJl$�%�sL�b>O�&G7�3���,Ɠ�a�����4%L��)��v���ʦ��.ׅ(�S\[� ��m��JB2��+�ѷ��\��7a��W��ڲ�/�Rwy�������|�fccR��#��&��:XvMt_����	J��p-J�3IV'��ccc����v�vvv�h4s�͌l�����^&ӥ\{�K� ��B��s�;...0K͖ʣ�������ZG�[	<��4���TsZ6���ٙ�|���N������"��LT�'�ze�x��A��W�>塅�P�9���0��r%�k��v�'�~���,�omm��l�Z�*�[�TP,Q(Ը��t���x��x�t��,+�;<Yi�\��a�� �X�ce��57�)���4j��.L���aeee)b���L�[��@��Xc��"���q�'�;��{�*�Q4öü��%������o9Ϧ�Lj��m��e��{�|J�QO�Q|��,D��5�E51پ��6/N�׸��}V�x�|U�ױ�����loockkKYqS�a:ؐ���k��l�b@�ƫ7�Ȧ1i�dyRA�z��^|�{�o2�������8<<T�h�T
�bQu��{��Nz������0�:���)���\a/���zj�u����j��[YYQ]����h�:Ǽ��W���X�&�R	������ŕ+W��R�DVR8�d��d�	 M����P�9r.��@:�臉T*���
ҩ4V2+Hg�
,���� ,�f��d;F�����"6������M��d��r��QI��KB��{��ܠ�� v�u�|�a�O`�k���X�ہτ�r�M��(:������7S�_��:}�oر�k��VWWQ�ױ�����m�l�`�������41�x�cB	t�L����$C����G�U�]��>����/��hIS+.���f��J�L��	-�
�F#�h���X� �ð��Ӄ�w�F#�z=T*\�v��>vwwU��|>ǳg�p��}<}�tIs�[8�f7LRZ��F����JW�\Y���@�k&s+m�$��Gc�
2�N�X��YJ��r.q��!�>�|~�T*�c@K*�������C|Mi[6�N�_����t:eE��ݛ%��{���0�� �a�MI�1��Q�N����
W�H�� ��d27}`��M�m`!��&�:��˾ƱXI�z����u}&WWc��1ܚr��nbԢ�DJ}K��ZW�\�͛7q��5��e�7��\&���s�Mu:���O�5\���N 5�L��Y��>7����͖�+u�z���Z�*����x�n��:��������X$�!1, u���}�8��I���|�����g?ï�kܾ}���T*�Fx����/���899�T�{_���A>�q�r]����|>�J��"j�X��ښJ�� VB��V ��8�es#�)���>��G��6�q���%�Τ�4��9R���"#{�9(a�}��jj���ɉs��m�
#�U3���A%]M�R��}�돂S|�H����U(�A��D��������7������P�.�7��}�#6�W;d�^������qŷ���%��x��Q���mv4�������ܶ��?�TJm�����z�*vvvp���N&K�~��E2���ɜRc����F�3���JSy�B�:�}2W�c�0��^\\`8*9q:���b�����I�l�F�\�~gggx��9�ݮ2�/��XI��R)��?Q7W�rc�c7�� �	�F#�J%ܽ{�W�_��W�{�.�\���by���������K��z�k\�y���Z����VWWQ,U�ǀ����`I:C� �.���n�|~�]��_���^Ҽ>^Yy��P�d?�x�<H_��H]�����U�r��~��b��l6�V�����W^�tl�F���U]	Z�Â�$5�q%NQ��>i���J�s�&9�kyf�ӌ��C��m`��l6�������lv�ꇾ{�7�M2�aN3q��A]�.$�eW�{ncMu�)H���̴@��7|�����	-5nRe���I֖��ڵk���@�RQ2�]K-�|R� ��Te3���$;,��d���P�V��d���q~~�t:�d��[oN#�%���z�F(�
$�C���G���1�NQ(���qqq�~�����tJٛ��5ƴ-p��CX&3�"�ȸ��<��P�Tp��u��W�����?��O����B���[&�A���իWqxx�G�)0��|�*e}𽟦�vY�߇,*?+��|>�`0���9VVV��[M�H!�<L9き`� �'dvg�ْ�`0(��1�+�}}����e}~�u&𦄂ת�� ����c(J����-�zLq�=�m����a�>L�jX���ܷ�i�B�=����Vn�V�¬C �E���<&}�J�ڮ1�uX�.��M�s����&%$h���x}4��4��F���w"p��ET*T*U6ex�d&�á�pa��=YV�1=�!�i�����d�$���畅R>�G:�V���Q/���Qn��\�,"��K&��|�cbY�P@�^�d2Q@{0(&N�� �$�\�9lZ��x����L��+W�������O~��>�w�����&VWW1��V�V�X�b�h�q���9���*[v�@���...��ɤn�+���$����U���'ld��<��]�w��7Y0�
�<��:�9~ҩ�r4��a~q>S�KYC*�R�����4�&�(�k+��bpî#�E���<�k��B���\��m��H�Y��Y��t>�t��aq��;��������ºN���6���������V`�&�T*h4h4�f�����K��Ro*.7�|>���*&��ү����Nn����5J��˙���0by�tBg7:7Q�p�}	d'z:��jnuI*Q(�l6������#�Ct:�ؚ�xص9y�ޒ��vU=L`��b��C�^��۷��_����/����l����9���Rp�d�%s�}�ߗMVm���䵰JP)�<���
<XJ�;�:�*����wd�.�������%ͻ�`����\�XVg�y���/��87+��������9��ϗ��_�2�B�(��O�ѿG��u�w�{�k_��kg[��ȼ ���rYQ����en��?2EI]�eޣ�t�&o]�gf�����d2�V�*��^��^��R��P(,�,G����R&��5�R	n��t�t
�����"����`$��מN�/,�s��#eeF�|�\C�C�5��t>8??W�E,��
~d�h�?qvvfd:�����i}XM_g�0�~��~�\7o��{ｇ�>�|�j�R+?�,SwK��`0���1qrr�d'Ef_S\j�+(��U���荕*J�%s+)=H��(��h4h6�h4�0��U�cO�ݓ�A�$,+����{�=�& "d������_�<K�5�d�)5����JD��IQ�
|�H� �����8�6a�]S0Qk�7�o�;��[}�0{�ۜD���h$�c��7��IF�Ndԅ�\N|���Ea��db������햕�M]��ښ��єP��@�J��.:��&$};�KpM\�i�2-�f6�)}+��Je��"s%�$��]�����]Yy��J����sR$K�.r�8�U��������q��A��>��<\�1��_�������G�Ν;h�/C㑲x"3I��'Op��=ܻwϞ=Sc@Dy�ALOTi���j�L��ip�*K����ulnnbkk�z]�i�%�E�א�����/`%��]�9%[�g/��b�@:�^�ʵ�f��`�K��ϒ@V��R6����CG�F��އ�R��ʱe�a����������Խn@�J��	9
S����ǹ'I`���a	���]�<�,��N���0�vB�����[�o=W]����eXB�g
(1m��l�RI�j��ժbn)' �9T�R�^e�O~>	^����	H3���=(��!斁�$�&��S6��R��� %@�Q*�RvEX���'�L�8e��%�]g�lM�vU>s���v�4���� �z����o���o��o��{�amm��Aa2V���|^5�M�S���?�g�}�?����t:K��9g�َ���و�63�6P@>�G�����6vwwQ�հ������.�Py  S*����Y5����+�E�l�$�]Yy�P��@f5(��x�?�R�C@,Y]	�y������Т/b��|�OX����}X�8��A�!jt������U|�^RItA���$X��b�6Q�aJ � 7,0c��+���u���HV��[�I�4'�4	�t]�mq%y�x�%X�\F�^WMe��� W�iʒ#7H���&�F�R$m��VQ^�4�^xܲӚ�OJ��%�a�d2j���_�+Y_2��������-_Ӧ��X.O��F�m��@��c�p�����>����|��X__G6�U�܋�eM�{�n�q��=|������/������LJ�etU����.�Ѵ>�i�1Y�ɠ6ir쒽m4ȭ�^����Ҋ��%�����E�a��q� ���ޏ���q���{�6=+�$�á\;�~�zY�I�R�#�-�hG����AA�e�ˮ�\{�Aq�Ϥ���c2h�⃤V�x��e2�L擓����J�>&�"K7>X^&�u�m��FMG	;���W]��8�{|�;%���<�2�����ann�j���X__W�zs��V�8�kˤ0�i�{��dɠ���6u�r�-�(����,��Woh��h6�E6�]��)	�_��s�Elmm!�����hɛ��S�<tR}�@�|@�7eW�����xr���h��r���k����?������������rq2E��W>�d���9NOO��7������K`2��\.+��׫�qW���\kJ4��ڤ	A�٦�*>�sQ�3��Uɽ�l�F*65J��9�q����i��º�����l�l���4��֖����<���6Yb9~�vZ���
��� ��M=I��,�Eloo+/���å47�!��<l�����e���=4.��*��!��~N�%�%�\l��P���p\��%��נ~ ��nnn~������ W��]'߁��0�ABr��mzL��+�+�|w���I�f�k��14�IRs��`'0�I�F�R��6�f���	����`0PL7=n�&�7��sʍ�`��Q�TJ5�I�6��,��u����J�����w��Ħ'6�Q�!-��y���q�gʀ?�^�U�Vd��I�ⲃ��nr���o�����t@͆��x�B���7o⣏>R�	�Q��z�G�f�*Ȁ���o�ſ�˿�w���߿����j5
�Wl�k��`�_��Q�sA�[H�}�%0�W�PPll&�A�\F��������~��9�1 FVL�|@�V<$���F��&L2��H5�nnn�V��J	��j�q�YrLrP��X�b��be���&��[=�e~1�t6}EO+�VWW�ܑa�M���K�h����a��c.���2��x�֍�px���OW���1�zϸ�:��������%e�(����V�����M�Ӭ߳0F�>�IhsmIj.�tRAL�i�����tb�Ǯ�L%���\�ZM5�ї�L7J������
��᳍�3����l�\.�r���t�
 ���Ⱦ|�%��q����{*��!�N�\./�l&��� ��E C�@5��Q�f�@�]�Ԧ��6m�:�l�$Hȿ�Y� �*[�-5�������v�~��㣏>��۷Q�ו�T��SV`�r�| ptt����
��������x��&�	J����\_�������'�����ļ%wq���y�������r�T*�r�bo���ҁ��#��,�L:��
���'�
��8N�JŒrmX[[C>�WzV�s���)�:b�.��=̤��Ha���J(���gҙs{�R���o�����`mm�^����t:8??_����M�ѥǍ�N���[�hW��u� ��N'IV�mR&��	���3�6��VMJ
�e\�F� ��	ܺ�� �)r��J�>���������:�FY<}m[��^zӚlcPA��@�ZU�[�U7%2�����Y�ڌ��Z    IDATJ?Y&�I &�(�� puu�tJ]٣�|��ԏ�_� �!J/]��u�̒�����T5������#߫V����D���l�b�����D5��-����J� �K0�5N��������rp����ﾋ_���{�.��}���`uuu	����V��o���������Ž{�0�L�H=&�����fu�#��,9��#A�Ϻj"l�	���mnnbgg�fS���� ��,��&� p�&T��J��t��`��C�����^�#�����2�ZvVpX���r�v�� *��:�-�b�`+�u�Ro��*�%�>ǃɉE���7�Vq��Jf_�9D�-�Gُ|�>�nԗ\J*� �?,�����K��r���ޡ3��J�H�g��(�m,�������Pi,A'� ���%�m&@"�gF:��3~mL�Ve�7���9��%G��@n���Hm6�1!�N��K�0	p%���=Y�浪����h4B��ǰ7T�F�J�n��}L&�b��K�*���sU�F�T,!��)PK�,���@�G�r��t���S�-O`3����$=�0�*�:A��	ӥ��]�n��͛7������p��-T*�z������rȭ�0�Nq||�����/�����?�������j�z�V��VS�&7i%�bӃ�"e�A6`��$cwwW��J���{�8�U��tP��jN�O2�|�BA�w>��I) Y_οB��R��b����x�z>G�PX���t�^���b)Vxee���+�\�� �+�myX�Ċ ��j)`�j.�p�D۸�������o|"��z�'%�J�^}��F��L,�kZ(}O!o#c���ӵ�l�'h�@n��q�=LIⲀn�&삥�u��2�N�4��l�^�+�+�lX`>�cv1[�n&�2%7R���,2�7z�~�ܔ��rC�VE,��w�1���y�s��i���W�\����Ţ��z=դ#7rDY�Փ�����L4#�&����b2c�N�RI�J�'��?�!@&UI�&��2����Mi�	��]���2E��^��>�}�]\�v����֔.��ܕ�%m�L'899�W_}���������d	ct��d2X__WU�U���S?�xݦfa�y:��A�4����vqvv�t��L�c�(O��*�O�W*T�Ulmm)p��d1�M������tߐ���@"c�k�*Պ��3���j�;��R��ݮz�<�������h4��h4Rc&�Nc����t6Ej%�t慴@��� ,5��R�n+r� �7n:����:677�n�q||��i�pFe�.��q�ࠠ�eG��%|�0����a�G�� \����x8	v3,x	���>��;3��QR@����{om��Lh���c�t���!�v(M�������*���×���b��t,���D?\��	�d��bɘ���x�z��`�N��(�
�֪KVd܌'�	Ɠ��+K��7�,�)��v��.p�CLj���S�.�j��z����u�Q3u��C�=bmmM�jȦ�b��ii��N���	���%�5����l���_fjJ���2n޼�����e�r�%b�'�i��)�?��������?��Ox��r_��)��������vwwQ�T�2)5���T��C
�`�3��v��&8>��.���qvv�v����S�Z�%k��y(K�dMy���0v�2 ���t�$���u����#�y@*�J�V�h6���jX,��z��������t��O�����h��fB��^�+�wuuU�b��{�-5ܙt�L�����	�w�X�(_k�)�@�߯�j���@���`0@��V�2�\'�l�VA��I ����|� ��{�_\��g�f���L��j�K��%	��P�r���� M��=�x���gW)'�	$�]���Y�|�LL�m��,���ժa�jUm���v��-�&��"��A�z�H�20K�2�uww�jUuj�)&�N�X,>)����y^�T~�X,>&�k6�
p����c�7O6��8����32��� C2v�܋�"��jޛN��t:�Fh��J�K@����;w�`ww���K�I�Z��C�z=��s�3�V����꒬A���Qǯ�F/渘��L���>��r<��#�G�����������>��=B��U�"�N�Z�b{{�o����.�^�� �	��
�_��0�A6�U�-�K�D�g8��n�qpp���=<z����v��?�/��l�"����d�� 0��1�{0r.J�0F��>C6�5�Mu�s�t:�v��p��#��+׏r���l�ۗ��)�/�i��nc>�/UXx`�쪔��R/��֛ly@�}��L5S�n����5-��-UFt�I�䫷N����Q=~m 7�>x� 7��܆#|$~���QM݅F�g�1.�@�c&u0�lz���!�-s���Q�7Ma6���|�˘(A'�(�S����d�8a����bk}4?��ɍ<�N��l�Ν;�z�*�ͦҷ.u��/�֏7ˉ��R��t�r�2lݥ�R���lll`gg� �Ӌ��O��|�\.�+��'?���?����ӧ��F�YYY�x���r����d����)���������
����r�$�x��c:�*�bb�| a���eg7ˣ�fS���T
�v�v{	�5ܼy���/���[[[�^�� (s2y� ��J�a�|z#����&@i�F FfN���P�<�N����o������?�{{{�Fh4XYYA��C�\�O~���W��{ｇf����	�����&��t@&���C_�%�1��ptt��*x�u�T����	n�� P�T�IP�%<�<8� D��l6[��s�f�Y��elnnbccC�`��ir�v���{\.��l"��~��v?Y,�b�����t.���l6��x���f�	���ϱ���~�?����d2�d=dm�ٸ�P�-�;��2��a2�����۝a��ʏ�d��Ɔ������a8.EK���`������.�B]�4�3D)�ePq���sߪi���M^�[���L�p��� l�Qd���%O�A�6L"6�m�k�><n� lU�o3��s	�QtN>:\�$25������N&��̰���+W��\./y��0�ߓ,)YM����n�dqX�m�Z�v�
oooccc�z��R�����j6��}r���O]���ի�X�������z��m47�L>n�Zh�Z��z�5B�ٳ�O T.����������	e,�JIB�TB�TRrJ7���T���.�~.����n߾�����>��֖b�	X��?N��L�do��J�3�{|=�*K����yʆ ڲ�o����ۿ�?��?�����t�t_xO���p��������֙4J֏�B�Ԛ�l�^���VV!��9��>NOO�n�_)㛾��%0��p�T�����C0Ԗr.r���d%)5�T*X__Wv_�n�VK�94\�~+++����O��z�R�����\�������N���F��p^*�~3��?8;;C��Q�>�G�Ri)���V��,�$xh�T�e@��6������H���:=Y�7  )��V��oQ}X��4ְCA�D�jg�g�	�'1Ug|]s7�X9I��u�J|ӠXJkD�G�.��e�9l�+�1_p��;]c#Y2_�VR.�d-9!$ ��t�,ӳd/˃@�����,��f�E)Z��,KZ����\.������q�7>��g��i4�&��N���o������Ǫ!�r�|>�%���vV��R;*}z�W�ScJ�J}ڪ�r9�)$j6����%����i����
��B�3IK�(�1��11�d�x}'''������_��o���Ǐ1�N��͔,�g2�y�Ke�.f���m W����� ��ks2!�\]]UZ�f��������C>cy�k��\��t֙lf�Z��Pg���8>y���:<T*Ua����ъi_�Z��r����\��q��;w�,0<x���d�L��&���GGG���K�R��B$���1���^�����(r��&�J��Z��N��;�)*Uo ����dEmDWX[�0�0�`��7�D�2��k�7����jx]�}߁4h��0�@A%_�׵p��������E{&�!�Й��t�_GzOҨ�Z�*�K�+��$��-��M*[:�8�e���l���Fj{{;]�T>�r�ʧI>���m��>|��^�o����u�ݏprr�J��BAi?�1���A6|���7`��JfI&����5��Y����7�j`rS�/�׮�J���(G�M��{�v���>~�����o��ӧOU����J6z<�bv��N���� �K\��\&�����6N�`֥d�e£d�M��,:�[2����F���h4���s�cJ�d��rj]yXm4H��h�Z�t:H�R�10��}Z����Z�����Ƨ��޾��;�������duu����9<<���	F���@S{�J�$6�QZ��Hk?���3`r���W�U4� �-�qI^���]�ۏ��4���	Q}l].D���5$i��>cz�>y�qNFq�O���IꊤsY}�>8[��֯�&�$|���x��-#yeӐ��V�zІJO}"�[ͮ.u�+p��b4�Ԧj���۷o����ݾ}�S �}rvv������<~����JZ�V����\.�f��$ZXQs(7^Y�D#���pC�����%P���������5u��eO�#���9h�V�nsn g=� ���&�x��ggg�����Ǐ{{tt��h��}�>u��W����������T�P�K֓����@Ͱ.E��� el���z8::���:���%��x`����t7(���^���b�d�F�dm�C��@�Z���u�j�Owww��X,Ʈ������~������U����X,�]�R����p� �8�^���a�TZ��d�YuЭ�f��8 `f�%&��P�s����Fe�=&�Oؽ'���\'4o��	eO׃�L}O6P�/26`��qOm�X?��A�Ȼ�Z}P����@OJ���>a�N�Il���8��-��񲓟�S:3&''�L�A*��jnU/P�7�h4P��?�֪�4�l�X����⵹��������os����z��ptt�n����a,3���n����f�Rz��^>/�&Ɏn&�	�ݻ�ح�h��ׯcmmM5F�Qn�X��I�V&Ɂh�ז��`0���{����Jx�<�929��,K2���j4:�	D���@�������&$�M���.uUI�@QL2���2�9�{H���w87�Frr���1�{�=k���Zh48<<�?����]�\.+0O )5�d4;������&�	n޼�t:�>���j%���xx�g�wb�E�%[�Rjqqq���}���O��矕�SjC��ɰ��S���AI,^�O^z̲ԪJ�3�����l6����o8@?�B_�b��n޼��u������_M����ĝ�h�sqq�f��j��Nd�6��+�	fic&=�BU0>��#yo�E$h^ؽy��^��
߼�	�N,�"D����	?-�1p�j#8]�z�?�"X4�zފ�
��+�`mQ��y^Q�V��vzo���V,-�=n�2Q�FV�Ѡ2xA2]��U���m=���iT*�����jacc�L�����o��_?|�7���� ���������N8�y��)��:�_��@�d�'�	��&Q.�1�P(P(TA=!% duO`���]]�V��r���>��o�F�X�i�댬��H��.G�3��G�$H�U���|/2��rϞ=���.NNN���.�����z899Q��^�������ׯτM�5��F��/�!����I��j6���������b�nxm���㧟~�ӧOqrr�f����Ag�x����@~:��P(����m�;�,�zY��M��[i�U(���&���~�����������Z�vo4ms���g2�D&��a�Ju��  ��F����_�z��	P�@'p��~j��_5��KĲ��SA��H�ƢŌ�s<I�nY;]0~�6;���N�$�̩M��5�����Z��ӌ�]��w��2�nY�V�`u��J���f��f��d�$`����U+++�_���Ϟ=���>��clmm=L�Rw�p+/�l����J��E���G���l�O>�����$��j���G�ZU�Yp2��v���TjF�I���0�U3�(���{{{��矱����?�׮]S��|���P(�&�+�
��& �!�b��D"���L�N�j(���v����ƌn�R���n:�����.�nϟ?G�V���!���q��M�s�gl6�E<G��R�yqq�N��L&�[�na}}�T
���rGGG*Ɋ��n�B�PD��VA8����Ym48>>����:�r�ˊ�`!!:�aC)�s)��'e�2
��w2��N[[[X[[{�)�V��ᇻ�\�^:��f���2*���R^��HS�HD��gY���$Gwv W������W�~zzSR]��	N��T�y''���f�ˇr2�79V2'@夕�kI�$�6���j������g��Ϋ�5���������N�v�M�bG�Q�ZF�"�e0S>��h��$=�ܔh(O[�?�7o�|���q�W�������_��}������szz�7�F�7�r�|�|^��f��J����3T�U�R)lnn�RPH���Oe
Y��Sޟ�+����z�V�(�˨V�J����H&�J���ulll ��^�+M��Ņ�i�R)���!�L��l��N��>-�j�NNN��Q�t��t:3��vkM�"НL&j0���+++j����b��l6�tʕJE�ꕕT*lmm�&Yggg*#�ɠZ�buuU�:3���t<~1�6��v�1�n�={`��	[�[dke������t:j��z=��`4!�N�K.��?kkk_^�v�]k�}������{���{�dr��ӧ�F�ؖzu�� 
��q�5������$��<NOO�����J�k��� �Eӷ�&`9�y�VѲnd�<�_��"1�� f{V���d`jKg:p6��V��
��aB�#��V7��k�����y��y��� ���ym!��঳2���ݜt��D"��x<�H8��x6��̛�X�R)[��"�H���L&�0�ɼ���N���������7�?���)R��a�E��2��	V%[K`B�+]%���|aD,흸)w:�J%T�U��#�X,���-lnn*�Ӄ�% �H$��К�&��]'''�����jJ�!�2$8�C[v,����1�c:���n��ӧ8::R���i:�F&�A�����1*��JE#8>;;SE���NNNP�וv<����"�N�^���l*���N�|V��MB$�%(a��$�I�X,��di���ik7�/%�&n߾��ׯ��_�������?���xX*��R�{ �������E���Ec
�/uȼN��E���#�M�R�V��{���"�|��J����<ΉQ4iN |YL�U��N�/~�7����3��C�e��$�5n�XL��d���$�����z~O@��	��P�]s�d���7edY�	Eg��dҘ|]2]�̱=����d���u������������򱶶�e���|ccc�����P%�e�Y����~�VS���S����@`F���fqqq��sJ�ɤ�f�z=�F#������.J���(��!���L��h4B��QZRZ�����'��v�ʹ�
غu��{=ڒl.Y�N���h��!>�Az�2����<G2t��ӧ�0�u�V��im�D����^��dr�*���tE~}��r9 @�TB(�'�|���Շ�L�˷i����?���p7�������Pf!]:���h4�B3.	,��U�1�Q�eAo�_�ҥï�&���E@�)�s�v���hg�@��ͫ�v��.����DV�f�^{n ���2�ޚ�K�`��j�y�ĉM;@궙�Ń�>�q^�jӗ�dTȊ���ħV��b����Շ�P���ٟ�U� n߾��ɓ'_N&��J����}��c��^YY����NNNP���M��&W    IDAT�[	X"����l�����a��� %@�������v{̑U�>��>R���-}��d�t�|׵��dR�k	 i�%�i�{�CT*��k��M�Lq��%��k�a���q�y�d2J�Bi�\k�^�ҙ[>�Ѩ*B�������X,��k����>~���X,��P
)1�w�1�}�Z/��D"%�bA��:_����ڪ�༁����� ����i�Y�a#�$��}.��'%/�|��=���zp��d�i6M?��y�"e�V9&Q�o�c'�o�z�ܹaHO[�tѧ��;���@[�"��A6������[�������������|�
��ylnn�R��8�r9e�&�"�¡0��<��Pm��*Lz�J9��ܥ�����	��@�b;\�Ч�u-1��l�ۭU�N���%���Έ������!cu�6�����c�u�*��Ź"�H�N�Mp�!)��Ţ1�#/CRxy,h!��5L��߾������������n�olS�?c�&��y��R��h��XZyA��T?��FjxM��i�v�h��;��	�y�>n�2���fѭR���_nMo-��w2[�7a~��ǉ�q�g ���vz�w-�.Z��faz���M�R������T �l�P��p�EL�o3�.mĎ���޼y�^���������J����XYYA�\V>�l�G"U�pH �#��`�����^��,����5��ʟ���:��ג�,f���t�sb^���L�����>z��;��I�|c��(G �e5� 8%�ܲ�3�ā@ ��Ti��&��)n޼����/����^k���=zt�X,�����N�V�a��I�#1�L
�f�A�:!ז�ѵ�>�8h����mnZU-��e�@7�Nҋ��kw�l��}],��y���&>�v�;͌�ukk�ϝW|o�x����d��urPЏ����3�z>;7���)n����rH&�#��W������?~wkk�^���~���D�cUw������:e�W�q�Np0(�6n�<�Ls�A�S1�_+��֖���8c8���i���bH/�e�N����p9����<� W�J�C�<�/?0���u1�Lp������|��Xk���/>}���x"�3�N�j�ԽGޓd烅�d2Q�Gv�`g"��p8T��ݵ���.� �l�����tw�Z������鐻פ۫8�Eo|Wy��"w�XZSM��D�݆�嘘N�ځ��=��|z)��6TӇ�Zʔ+��4�a*�$A,{�J�~����V3J�q���_���X,��`0�S�հ���\.���U5���tT����,&:��p!�D��x0T,��2�K2�R��3�V7f�v���ɂ�m���nօ�����y!��Xڽ���O
�\����^	��2JYZ�ѳxee�����r_~��ޕ���f��N���嶩��cW��w&�Q�w���nG���|A(�4���ȶ���_�J��!+��y��yfl����ؘv��@����&�2!��,-�ߦ�o�Jp���l)L&%���I��p3����o��:5�e8����s��]�]c��J���F��ޭR�Ș_�r�#�b4���-��կ޿�~ ����Q.�h���P�fRB@�K-!���!h��Z��lرM&������RN>��^ǋ�n`�j؍��JKl�Ͳ��eH
�u8�B[�b�P�ScKP+ύdri��L&��'�`}}�a"���]Zgkkk�?~7��.�L��Q����NGY�ɔ7ʤ��!z��eh�x�����_$Q6{�����z�L�>Mc]���nPq^�ϼ~�&s-�3Vf7�7�a��[�t���3o��2�`��jReIF�*��T_�����0��^'��:5�e8̋���D,��F�N�Q,Q,�J��h4���S�XLY/�̟�[��z1 �;����O#�l'''8??We�T
������*�l<+�U����d�[�<olŒ��pqb�6X�kҪ+dr�_�6q^	��v�	АŇ��V��g\/�x�H�'�_�R��� }qcc���677[(޹b������?�����������%�	x<��^O[�}dG���Q\,<�`�l7\d�&휋L���7{a���+������q�{��������hJ89�_�&�&QX�	�b�eWy:I��L�6S7 j�yM�ͩ}z���<�ub��4a$d+=�H(=�L���!��uU P��H�a4����D"q?��fmmm��h���`0�x<���JRͤ�����q�<��u��I�+��&��Mҏ(�y���[���鰎�=j��.��,.]hYE8y��p���H�w\��Hkkk��Ep����jd2��\.��� ������J�uD��)���=۩]��~>�p�S���>0�z\6 {&p;�c�_;��Wɛ�8���9��<;�[�ҏM�*��Iԣ[Ulw��n� ��e�Zf�J� ���^������q����o�����׮]�9??W��lV�n��R��R����#�zJH0$5����$���tP�'�]�����4��unA>X�����
�J�+�[0� x9���P,���|�AC*�������vh�E�V�5暡�� }�	p�3J-���������$�m�3�$�4Onz�X^���ꏟ���W�x�Փ���U|�y"�M���U�ɿ��J�Qz����P0�X4�X4�6ɘ�Z-�j5C���d�]��������*��"��1���J��@U��?����H^�!�*\�^9}n.^֬�=�]a\��JOf�s��{
;���TP��A�~L&��eQ
�.���L_ ���SC�L&C��:���x�D��r9`2��Faq��v������zb 
��س*$u��n�X�^ύ1v��M�z�y���h��>��&�-��}S��2�������\��y^�8��=����U��į���d2A��A��@��T)d�f>�`:�"(�5����F20�L��v)YM��л~ӊF����������Z���`Y4���Q��͖�{K��c-�%����Gv-C/Y��^[o2�e�aU8��V��а�rJ2�2��bvGc�'/���f� ��<B�Ѓ`0x�]_k�T*��=�L���k��t a!N[5��7'��0��Ꝥ&�N�z^
K�(�y���|\�kx��p�l��p%Y	��0��ⱫF�J�=���d�Ư��78_��s�)��?jS���:�0]�|<�5�WL���+�`�ykk�_������ڃ`0x7�>H�R3 E�y�Z-4*��?Ҏ�1�2r�-Y�0vܲXN�_�ul�V��tK.Y�ݿ��K��H�[J�Y)�x<F�W��,����<�����������FC�Xl&ю)�tA��%c� ��t31!��c�3�5�ū|�����bJظ}./��$.[��'��:_�<|�ܫ�tI�~�wZ�n��V�DnڠE�V��-�w�u�%��N�)����L�+u���1��h�Dr0|�;�<>��Ӈ��O�t?�F�JZ@3z==�ZgW-����&�8nj=�t���捓6��/�Z�Β�sbb����$K�d��@�u��pd&�L�N�g\����F��b��t:�f�R��{�֢����x��p8�#��ʂ� Z�z��� �<�_����>i���o~���nM�@M%Jn�6�� �M�M�u���{���%���y��i��_zt����q�s�ݪB�)S��5'O���r�쾛��И���O2Sd��
�- @ ��p��aiD&�X,"�N߿}��;�(��8�� ��^�t�DB#&Rq�L&���3��d�%Pb���7���������p��ӑ��S��c?�E�>d�@�#��X����5D��\�0�lD�xIo[�p8��t��:���lr]���f��d��C��G<�`0�����^������ӟ�
�����Oh=,��J�Y��O���c�xL���1	�V�׍g��Q���y�����	������[4�p�l��Ȝ� n ��b��3�N�l��y� ��j'�7�ѵ�Y�$θ�x�MS��c�r㰺a��HZ����X�m��B8F"�PV2�D:�~�'���dRY{��u�2%�	j ��[��d�`pFCH�C.����!Z��b��A���Z�p����9�wL�Q�ǫ��J�Kl�S�L��A��w*����=���l�VKIV:���G���p8T?'�p8T��D"�^��\.l�Z�F���K�vd�(����O�=�J��x�3#���0�e�����~ �7�2��޿(�/�K�}P�J���'!;��`�i{�л}7��ŗӍ��r쾧����U���AQ0T)dd��!����~�^oF�����E����ޗG>�G��B8VPrs�F�D��%'��$Zm���)��M\9LE=/�+�8�35ux6��,���H���
2������'��t=`� �����@����얄�a$�I��XX$�xY	����tex_<���nWu8�m��.<>R�l���,��������<�ג>�~�?�S��[���`�ݽ�)tB�*��I����^�\#��C�D%+i�ńz��2�{=�~.;��[[C�S��N��J���f�J��H$  ��P�N�2�]z�����`�Ax���B��z��p8���R��G�^O�nH��j(F�pu�7�x<�b���7n�/���9��Df  7zӴ���*Lz>��$	$�Id�Y$�IܺuH$�Z,�����x\��J{{{x���Y��u��02���&B�Ќ5%r�ӊ=ץA��#���"x_g���}�ǎ&@��R׮_�)T���B'"I���٫��6qm�R�m���\�����^�/�m��޶�������M��iv�<��	�l�@��p_��L%!NI5�7��DԆNP�MD>���jÏ�c�O�э��-n���U�~_1�U��WR� }p���� _&�QL��@��m�j�W6?^S�����`0�I�2cq��MB[�u�4�/����5ܾ}�n�����_����MunX<���Y�@�����	R����pqq���t�\2pR$m��v����X�*x-1��}y����N�7 v����ؙ��V~r� ���� �.9��Y�e_4)"����:�T�\�.�S`�۾��%�:\~���\/Z�y��2.TX��V�2/���׫��k�<�O�e+��	�kz=�|V���<��-�_�s���s�W�+[��d�dR���65��8qӕ�9�տ����ƍ�u�VVVT1�F�j�P�Vm�7��6��2��ΰ���R��4�,XL#Mo�^ug˼nz����8��,�_��_����ϰ���|>�\.��-A?��]�I��F$���)��4����|A���G: �Rw+	�_����y|������������P0��{�,${+	��Ig�^��
��͋آz\7���Ǻ���(P�����E��<a?�������H}���֋&u��cZ�]U�u�L��b�kF������(YD���5}y��q����@��zʭ�f�<�����e����`������>��c��_�%�]�� 4Yw�5���Q�T����l6�~�gggh6�J*#���v��21,�����5|��G��O�������M^����]��^Ŕ��N)%����J�6��$�(��^<[��G4JO[YxHٕ��(aJ��[�7�8�&,��@���CY$wQ����o�5�u���ۂX�C�*bO?�n��%��@�N��e��:iP޴E�����10YT�������@`��N��o,�	 �7miS���=�����q$Ú��1�T��,�����H��	p��)��6B�2�666p��mlnn"��$��]�s�6oF)�E�At�]�&v�]GP���k@�u�w9��Q
$�I����X(�X("�ͪ�>[]C��]d����@X:��9��W댢ԃ�9�H��V�d�X^�����6?��$~���������q�N�c���.aj��Ў���9�D�B�+Q��zQ���ȴ��S�b(���0 `����Zi~�LнH0�*87����`5��2��l��4�r��,��$Д����c�A2�\g��``�`�#�A���{W��c��ZIZ@����f���t
%���p�z]���ׯ�ڵkX[[�t�x��Ԧ~iT��y�D"(�3�^K'''3�^;I���t��������7O�w4E>��͛7��`}m���v�h T���5))�&��e�|���8�o��B�D#�3'r �EO�ߟq�x_''';O�<��R�(�Zt����a_�#)���{Դ���]*��Y���if�M�c�959Ǧv}~ݛ���u�����܄T���,�&S4�	^�,=�l^]�i�bQ?Y��ͩ�u:�&�\7���Y�������j����݆�R��1��Q�V�L��Tr��UZB�c�1?۬|-�g��A-�xx	HYpC&cH��`0P���n�L�|���XYYA$A��E�ٜ�n��7w�[4E*����&>��cT*����Z����:��k�Ĕ�-�ۏ"ߩ�b�t:�k׮�����裏���ɠt:5�E��;D�Q�Ca�Ƴ��dn�fⱗ.R�K�v<������@�����ʢ�r"N񞬳/����d2Qul�!Lq�	i��3�/� �cI$�2MΉׯ-=��i4}n�����I�����:�PVL�W�x���/��o��N[�_�ȣyg�~�p/`g����m�P'�kS��d�5�9�<�vj^ϥ����~�J}3�Μt֜����I#� :���\];�X�^��ZΒu�6]&� Z<G*��5�dp� �����d'u���ښj��>l�n�יT�D�y�s;�0�L�-M2�D.�C<�	R�c��K�Gp��ID�+p=�¡�aL��`0@���x2F��ye���Ȯh��/?8$�>=���x0`:yy���h4B8V��F[0�!c���M�=�4��`�	�0���*W�l/|�AIvŀ����s-�3i�\_yЃ�4��U5�L�����+�2�N��U\P�]/j��h�,h�l��(e+��;,7`isdW�H�R���/=K�N���`��--�䠌����H��J/��^2��N����N����m�z��� )�"�͢P(�X,"��sn��۱nט�ķ��e�s+����V����l6���� $����N&\\\�\�,x쏎�P�Vg��hw.=[i#��1���>N7=�������+�B�ٜ�z=L��=g8�k���t0��]��-v�Oϓ���~6I��;����6/���{y�v3-��y-R�\���W�k��9��k��/Û��&eރow����ݰLA'M�	�v;�v:��c��$p�m7��Q���}&ߧ�Tn�L3�B��b*�7�J�x�E*M���8VVVP�p~~���C"��!��Ͱ���Zi���.��L`��gL=���n��ӊI���
��jh48??W����M
�daB�,}�+��j{��h2��T*�T*)�*�ˌA[���V��U ��/NNN��ڵk��5vtt�szz�E��P������&Tx?�Z�ÅN�0�}Ս�qj��3�f�&��������n�����`V��ڝ/ѼN6k&�'|Q��	�u�~���Ml1���Ci�z~���A��bq��y1�Xs�)X}W�������p8TVTԐ��$0Vc�]�Y��D��B��QS��P��(9���K�����~��l�V�R	?��#R�&�	677���FA0��K������� ��K�Ъ{#�������>Ъ[a�q���������\.�N��2�,�L΀U���vϟ?W���L�<��~����˴�S<W�!�A��5&���R��6����`0��;p'�� v�A��t9Y�K����s;���Xu���\�M��
���M���<{�UZ�\V]h�x��;LN@��=^i�    IDAT�w	����$.��>L��$�ٱ�^��Ll��i����S��e��Nŀ�)�x%J�d�^f�O�͗��bK��X��$
���U��G$�����_�����M�����	�%��d��G-�7t��j����չH��8==���>�� ��*������&���p��lmmauuU� 8E�\N��R)�r9����T*�V����Y�z��F��3/E���δ�"�+VWW����t:=�y {�1pqq���=����ǏQ�Vu��ք����U1'/l�(��͢����u�2���'�V���q��E�۝������Y��Y:���,=���`��ya
��'W=D�ց4m�ۑq~�L����_/j���=/�~nN��!,S�W���jŘ����zM�����K��2+B/��N~�V���c����d�@8�1�L&iY��`� ���`�ɓ'_�{}Ō&	L�SD"$	�t)��u��vQ.��N�����D"�X4���<z������r�D"3m�\.��>�l&�K��%�sG�/���ٙ:�v�_�׍�/�]n�vl��Ѳ��]ӢZ�������������O�W�	L)�(�J������?�8VP7�cOɇ> �\�r ��.3~%H��OV�pߋ�I�^�)"��D��}0��l*-4�ȡY9S@�+eU��<�@v�v���#٭f_^7��]$��5���n�gVƊ�^&Au�Ņ���{�e}q7��EX]}Q�&��q�LM�&�6#ӡ5��c�@�H��a��<׉�����&�Mˤ*%��e���a�N�nwf�m2��<wj@��h4��q����@`g2�(��Fђ��7e?���7U�X&��d2A4v	���*NNN��͚6�rY�O8��ʊ��"��H�R����/~���a
��}t�]��[u�qN��L��d��t2^�^� �A3�ד�E2,�n�E|�����O�W�W�}�6�ɤ=<^��F�VS�fS�jY�H�=�-��M��%��%z��~O�@t: ��Q*��e}}��-(+�������V���d�x\�qح��4�#_������-A������˝��xyܚ{B~I���<6fN칩Å�`���<����2;�^ρ�L�~�bp���"��<`�ϋ���!��&-!����`/�����[XX\���4�3�75ǖ�YP�N��@2Ul{��"p��z���V��F��L�\./..0���&�
���Lٖ�-���/V�_2�2P�(u:<~��P+++X[[C*�Rvcr�H&��v�rm���P矖URRa���RW�+"���l+�V	re1o����&>���q��m\�~7n�P��W+���~��P(�Ϋ�FⶹX��"u<;�O�%�(��uU.�����O>�d���|�.wL:����h�����kp8��h`0(ͻp�^��� �z]Y�I�7��Hb��m:?�DbY�RM�?\ ��uD獔7�l�an�Z}=Zu��H���0���z/���q���z�������3'I��Ea5��;ځ</��W�o�C@��9�˖�'Y�P(4Ӷ#k$c1e{�ޜH�R(
����O?��spp�E�RQ� �`�-��<�2y,�H(�-_7�H̴^�`�{<��*=e�Y�%;�D��@6�Ň~�
2^N W^�v �jMY\�`���ڵ����2�%����,$tɄ@cBr�AU<���"�kBOV��$	��cT�U4��;���_�����ѰV�a0 �H(9��F��z��@ �t:�d2���
�� P�Y0��:s?X777%���K4�U%�y�(����z�γ���R��y����`M��x��kp�L���ЙՁs�&m�e�J��_�y������K�����U{LƏJ��
Tȡ2.~>�����0��Ǳ���d2����Z�ϻ��N�\F��W�@2G����3��<~��.�O$Qry]���K�ș.'���`a��m����L����Jb���m�R��c �O�Kؽ�d<�x2����v��mkm�=�s�7vצf�:������c��)��M�p1X�^����[[[;�l��dq�����?����ٙ��q���h�ZJ�Cɂ� /� <�:���d^��k؀i�������5a�M@�[�<>0����'�ν����Y;���"�� ��	���3��	�.
�L��&���"�@{qq��S^�pݦS)Q����IZ+ϥ�.��������/���;{{{wP.��{����r��V[Ҏ�`X=ju�����ʩ|:bl[��QA�DPE�Њ���8y�\���@v��,�a�z^��MӔ���-���o/..f��kߍ����x$�f3��)�Ї��{�\��TJ�������ӧ�Ecw�>}��G}�΀ܓ���N���p�]�Tf
p�,7�W'���Z�,n���A^zr�[Ѳ�~lwm��0��a��U&��n{��4�y�I��n���9�|Xu�⃻V�*��"��2�^-3�A~>���*,b�c=� ����G�`W�9�s���V���uR�iU�IP�"����O�~��G=|n�\����b���T�����$��>ɠK���#�*9���&A��Z��#3�S2�C2�V�<���J,�sL0���|O�u+2;�	p%x׽|y�N&4�Mc����t:���PA2�煬c�^W̿d��[�|q�3���n�ɓ'X__߉Ƣ���l6?o�Z�'''j؏E$]$��j�R�Z�������Р]��	�:�y�ʷc7���f׵,�k�Y�CNi�WE�ٝ�����N�G⤥ \;�b�՗����l&`�	���Z7Iv��;�U}yI����=�v�����*��j�#WJ+	~d+����T(B��C����F��������N�N��?�c���������>��4��,��j��h�N��4˲5���8Y���_؉Q��m�ɫ��5 � �/�E���X(+��.�!3+/Y	B�Ϥ�$;l�Kf��1�^�r8<<D�RA�՚ig��Zo��H$� Z��B�VC�ZU�J�e���w3:@��u���!�J�y����۷o��E����������O����PIpxݐ��l��H�0������p0�5�r���i�lf��sK�s
�sO���M�^�/'�ڋݘ���	��g�}R׵^�#�L��9Kcp���(�lYQ�n�#v'��y�N���B��ZT ?O���|��.�ºݮ�D�)�d����߹�1�T*H����x��b���������������ө��կ��)�$�t�f�͗�Xn�dv�6>Z�u:KK��B��H$��������[�V����/�SQ%�IY �\�zep��L�����d2Q�����8<<�I's*���,�IzQ���F���qvv���Md�Y5\��D�6�H(0K�&���i������������ʽ����^�~��^s�v��v������j5D�Qu|��02��*<d�F��d{����`��u��I�i0����p�U��~�Y�?�3l'�p�C���L�\6��B���4�%�EO���]�Ԣ���*��ʯ��b������9�7��yRҜ>����Ҧq�(M���Ώ�f��{��mT*������A�7tɬ�-�j��^�w����wvv�	������Ri��� �^�x|��V�y���M3zP��2���(��,��)J���c����^�c?��VWW��d�J�`ҭ��{R?,A���o�ṄS�J�iH�M�~���m}��5+y��h4B���y��������ǯ�0������`0@��F��C�P���:j�Z��ҊF�Qt�]�z=�k,��y]I�(;��0����d2��P(�V��������ɓ;����T*j}1���+�F�K[=%Nj�ym1����RlY� �^��E�����)=�
�ͫ-]���ɓ���Nh&$�<Ci:�`�G�kV�-��~�T�E�����Խ�	�'ЏI}?u�V'pQ��w\�b��,�+&L��ʲ�0L��]�/�����ב��H$�H���8�I�dy�^0`;kkk�����nll�� ������߿��?���L�(q�%�g��)�bMN�3�,�L�P( �L����z�FCS�k����ϟ#�"� �L���ߑ�z��n�/[�|��d����A��٭	Z�����x2~EK�[�9i�:<�d�����88<@�TB��G<����C�����Q��a��y���(��A�A!x�p�,&e�D(B*�bgggg���o1�N�<z���/~�n����ۇ����={����3$�I�r9%=�9�k�zd=[Z���3�F��f��_�k�Dh��4��t
�q#aܮ�y�)?�d��"7�a�r*���r�w�S4�_��d��i��Z\X�`�zڔ��hbC��@�"�S�9�{[����Nq�~�V�~��]Q��L^\�����O���n��h��n���B!L1U�F�V��C����1���v�պ���w��>x+A�?��].��J����C��}�r9
��iD���!C�pˍ3�7�l6�b���x�N����\\\���C��;��.����DP��q��Md��Wb{	�� %VA�f���ߥ��|�MVZ���?�>$�d���B������h4�m�ɘ�$�8U13���e)d*�&W~N�x)]��b�>.�����dr'�{���ݷ	�l����;==�~��9�� �_��x<� ��a;ݿ��,�J��b�����I�#� ����� �~ @�{�W5;�L���oI8�	.V�U�l�L͘��~M��y�Ye{�|^��&˸]�~VbV��>��WaV�bn7D'�lz����:܋���-�r9�~�B�N� �ʠ��+�̀��@����px�X,�;99�{�ڵ�
䞞���nooo��o�A�VC6�U�m$�����'�N�/7�P���Gc�'�W�������r��j�v����@�VS�v�T�������n�����7n�P(̴�nG�����VU>G���Q�v.� ��K"����7X$�mƜ���t�|��5��E�^O��Ѩ�X�-�d2�~��4�$��@<f�l�d���o`;����~��go�z;>>ޮT*��?~�~����U%�`�H�i2j��Ϙ�ӽ^O�x,���eA?-'�ΕxqZ�>O����~�;�������\;�?��pir��0�o�2��{��M�.�`
\M[�V6eNѝnz_�4�yt:������f��ud2�b�C  �)���V%�j�pzz�@ ������zk@��������o���j�im*Qi:�^��T�o�� ��Ɓ�5RO�M;�H ��8�f��^���������
���@�\���+�	�����W���Vgp���u��u��۬�L���jݺ\E�s!�Ĭ֥��z��z��d2�x<�N��j����s���#+_j�9��%�q�[��q$	lnn��n�o�A0ܞL&���曻���/�����ѣ����{\c�*��iea��J��r-QK�s����l61U��x<F�wY�3 B���5^�:�z�H�Em������vd�V�Y�Y}Fi��c??��.MN�,���.UA�d�qAXh��4vZd/�)���*c��)�@ �v��z��v��ҷ�Ѩ�<��3�I�#�bVN93Js:�n��{���w����h�{pp��j��|��7��O?�V�!�Ncss�bQ��d�$���ˍU2N��"�%���Z�ZE�\F�^W��z�҅J@DPI��.A�[�^'�)�0 m�$��%5:��yY�v,�S�m�#/���@����G��c4��eu�L�S�j5���P(`ee�LF���.���R�1���d��Ű�����]�����h4��������/������ѣ�R�towww�ɓ'��(�H�ӘN��V�
�������!(�TJ�H	���1���B�E��L��dug����5�b�^GD��^����\y����N��6��t�q�H/y96K23y#/m�7���ss��
��$B����8]�ݬ�>�);�3e������<7
�+n
l�I�J&��g���'�e�KV��B�Z�l�6�7����矷�������v�TB�TB"�@�P@�P@6�U�uz�m�X,������:�F&�A @��B�ZE�VC��~%:���X�����2���o���א|o�l��r�����ҢIP^\W����_��|��݄�<���U���� �D��b����g�)o�9� ;�B�R	_�5:��N$ٙN�{ppp��͛�}������j������o��
��R)�t�h4T���RK��/�h��d�嚘L&��|��2S�;][n^�^���Z�Zׯ�^%qۻ9& ���O�'�UBi�m��e6MZ��JoYƠ�<�K�3[ŗ:]<&��<q�vI4���T��T@�lĒ�"KD��f��X\�p3f۔���E�k�r��k�@���ظW.�ﮮ��Q ������z��������#��P(`uu�d�r�̶�� {�J��N�/��ݞ�`T$A6�U��^�d��|�d0:�%�.'��������79e.���T��u+&��n��vk�ױL���Q�=l�ۨ_\JOVVV�nv?����4��"R��ͦ��Yy ��R���p��5D"������F���������~�Zu�'''��F�l6�����'''�+�j������D�'	DcQ�;�b�畲:��F#Uh��k�?{���J/�D���n��U��t����x�t�]�qX$~��2�w�+�irL�^Ji�\�$���V���m�e��f�^�~��]��d��p~~�k׮)0��D,->2)�="[\�/����f�^��ٳg��۝N�����/��/������o���������Q*��F����|>���)���j'K&�ѡ�T
�x�2f7�F�a�x�|�l�V���8;;S��<�DWʢ�k�	k�>"�l���$#mu}Iߩ}���uݭkbW�0Y&k��}VY��/oݺ�|>��ׯ�Z����{{{�v�6���G*���-�*VS����b�
�A%���{j�oܸq������_���W��*���4��;<<��ޞ:���N�hw�������$�^�\,(i��s�uC�U��Ua�F�8At�"� 6����^xzrw;�[;�� ����9�Ƈ���y�`�xMS�e��ңZ� ?b��p�|�.�,�E
�E%�P�S���@�T�U���bkk�lV�4���̈́6crXCOj�Z
s��L&(�J�FۉD�w�}�ݗ�d�?��h���?�����www�J��G����X,�X,"�� �N�hP��n���p�Z����:�(���)C��<::���.?~�j����t���_��S�?�����fa�e�r����UAw�E-?(B��B�RQ����:VVV���� n�P@>� �0��tTW%�� �H��L+���Ǳ���h4���3�\.������������_("�H����_�ki�����h4���l���coo�Xׯ_���:�� �:�������:��\G�,��sޫxX�W�UT*���WdV^��M��y�z��^�zN���Zvrz� ���μ��U���&�Dx_���Uo�0��}�TlnzT?������"6�n�����.ʹB��x[ٔt�]T*���(r2� �J)�Gf���8�(���N;��`��������2��\�0̿�ۿm�J�ߕ��탃��ud2lll �H �J)]��i �������f����p8�d2�H$�n��Z��Z�6#O���bg^�C�ԼN��_��?���"�S������*v� ����NG���Ce/F6��8� ��dK��v�l�z?��NOOw���w����o����/���W}��o����h���~ppp�V��4�Me�V,���N������U�����:�S�����`|8�jj����qqq�
+R�0Y%my�
]������{���׳�x�EA����|�*�>+�`g۪&_���<�^�Ƌ��96-�    IDAT�t�7�eP�N��ɂk�V�ׂ�?����M����n�R�2�K�`&�t&=����;I��ʍi2���gmmm'���;O�>�2�u��u߁����N����Z���Ƥ\.Q.�����0�N���f;�d�	���L˘L,S���Jt0��2=�k<+ˢ����et:U@�$\����}�:�l���"�)����h6�8::B"������4VVVP��pzz�Z��k׮!�L�D@�%�I��E��������D�|�T
�v���899���	�������ᝣ��;���p�X,��,VWWC�T������,��;�~��N�3n��h6���j����@ �spp���=�̒����=a�כ�������r39�k��
��L&��!sN�\wNp:�NE���.Rw��[ga�pIZV��l�^?�m��U�^�k�Go��D��,��M���7N�D�M��ע���`�*C?n�Vǁ�LN؏F#��ub8^n�7�H������<un���_Z���V��A*��a�J��2��N>�߉��w���?}���/�0�=>>���z��J�;�v{�V\h��*&��PRG<O0�^~ɪ�b15�E3y2hdm���R�����`�R����]���*oZ��*�qW	��Ҡ��p����m�� {���"�]j�j�p||�t:�t:�T*��7o��	�B'�x~~�9������d�5��c��f�M�R��������o0�vR��N�ZE�P@��F0��?��?�O$A��4�L&Ϟ=��N��B��F��B��Pl-�\�����a4�M4�'=����r ��Z�z����O��v�J��h4TQ�{��ک%<τ�~�
��_���".CN��e�޷��E+�&<���d�q���u�m�.��XeS�	����[��{�i?�=�����m��`�F��&����+�d�ߟI��{H[�@ 0A�.7�D"����8??G:�F�P�I�R;�X�������p8(7%�7��rC���j�&Ϟ=�"��j5T�U\\\���_:$�H$3��Rj� z��ө�.H����l8b8*��cI�`��W����ϟ?W)Zr�ˏn�Uh�t�^7���a��E&��b��,0��H��Q(������MP,����d2�\.�R��J�0fdB����{J��kt}}�P+++�N�������vww������u
��t:��B��yxx�N��
W�)���d2J�T(�����T�̮��2U���~���ǁ�x<�|�	���X�^��R�����J%��}%5�c����
Q'&���/�uY����x�]ބ^_Tof�'q�X�"~Ю"����J�� ^50��E��b�'s�=�K˪V��N���[d�Oo��u�>�������M�� 
���p8��dp���+��-O��>HzgR�(�84������@ �L&�d2��t�N��~��x<c8�?�+�A_Z:P�|qq��ku,���e]���:%-k��3-{���'�Z*���f2����F�/��@��u떺fB��*�Xd@�� ;2����b2�(0�L&՚&�K��K����`2|!�L"�L*P���i6���m�� ��,�f�!a7��]�q_|��`�� '''h�ZJ�����go5%f�ݿ�\�\�i�?�~�/��xu��r��4f: ���y@�p�:T変��`����Ns[ݨ^��
�������p�:�FPGstF�&��1��"L�X�n
�`�C��&F H������c�j5t�]ժ$S%e�X����H1Cd�h���������g4)P��f��0ťwm"�P�d��v:���Tx4Um�H$��d��d��Ζ-��ܓ�0G~Z瘬�y�oN���ڠ����j5��a���!�!�����O�<�d2���
6�m�ƍ���3���KG�lF�Q�}�}1
���`0P��Ԓ��yl����6��0���}Wޗ���X�X�xL_�c��
%N�9'���A��X,�
PYDO�SU�������9NOO����B��6��{up�y����Lq��^�E�+?�y�ح[��"�&�
�ev�M%jK��aX}8����d����Tv��ۉ��1��,����*^?��������V9��Gx:�����%�� �<���ZM1�l�mR���O!A�2�~�.I�1`�{�X`�B���B+L�ڴlk4s������p�iV�~�v[m��|�H�TRI����s)k��a8�L]2\�b�FC p��r]:�3�ֳ�aɁ�N�~���Q�ZY������b/�w�Nԏ�,������F)�A,����_��>� �n�������qtt�F���D	�Y�qh�k��`���F�h�5(���]O�� ��$��L�t���
�� Q���r@�k��V����,�e�,x��BF��{������\I�� �i��t�1!K��+B�jO�����S��-�Z�L}z��Dv��^XQ���*`M�4��^|����΃؝�,�L���d1��h�S����w��u�,v�{�6ʢ��EҔ������dA��H��&��J�V��^��F��r��2���	A#/ّH4�(�3�!���������h���WWnfܰd�0�7;~g�)���x<�
@�s;�"zYv�]�Z-�IN�G�j���Ȱq��d2�g̑�Ug�mJ�t`�i
������ia+?���dnL����
��u�����俇B!��}#�>@&����&��2���{lll�����P,���@�8 Յ ���A����YJm.;'ҫ�zs2���L@�w֋Q�@�.	�:"ДZZl��>�n�K�B^;�aPC_��Q*�prr���P/�)n���^m��z!zL�kEz��{v�[�γ���ʪ�u��Y}_'����JZai�p�nś�8�X;�U!7�V��d�"��duS���_����j�_T��k�%ϓ	���2�>����m�F#4�MD�Q$	d�Y�r9�6��Bᙴ!�ݸ�qxK����G<W�l�:��R�'h��|�$5}|]~f��>�r�Nl��s�'cƁ��^�B��6��c<�R�����RI����2t]v��S�.�k�['��6��y���Y�vr37�B���h4pzz�\.�b��B����M�j5|��w�����V2�D6�U�����n�Z��T�:�S�v/�2|.N��k,�!�\ǣ�H�����i�+�K�l ח\�R_K���%��V�U����JEi�e欺���%)�3������u�^�]zി��l����Iw~���+���3�`�je�4d�h����~z]h^h��po��JO�w��oR?fa'[ѭ��,֬�]������p�T*�6���eR���Cn���y���G��W @�t��%�#?�2#���H�V����rc�FJ˗���e�Uj�i�&Y$�_<�,
VVV  �R	ϟ?���1���m����tޖ�i�E4O�̢�IK�/o["�is����h4B�VC�TB"�@:����F����"���?D>�W �fR�#�G���D0}��	p���L�˵+G%`�D"�3�[:��ie��"�,3;1�NG��X�:'C�l6Q�V1�����t:������ppp���#\\\��!�X��z�ң:]��y;��:��[�}�{��<��{��fg�赛�N0�n��Ӆ�%��m��Kƺ	;d�H��|N�+�J�j��|��P�׳S��s{M��r}S��@�����s����X,"�N#��\n��ڝ�ZRnLVS�����lJVI&�Iֈ �������Kj��� "����&��_�XLm���JF�`Y�o��l"�cssS���x��)~��g+f˭��ḩ��^_�v�!������͉��k�u�v�i��R��T*���M���b4���O�<A:�F.�S] Z}p�v���,h�����(��zQk/�F�s�K�:#00E�=U\����/C����6�N�n�qvv�z��\��(�*�
���qrr�Z�fF3O�dw��]��N�c�� z��Y��ؠ���ZVHּ׏	&[FJ��`z�6�]ण�=h�Y�lF�U�iS�����z��m[9�~M�!�y��a+6W��-���-�b����%5�t7�������m� f / )# CJ��j�%�%�C��'C�D�1^Ig#P�-]����\	(S��bX]]�G}�T*�X�Ǐ㧟~B�јa����E
:7�NG�&ű[�N���{������e���8��!�R��	GT�������O?accCE�R)�%+��V�Y�\�n�4�+�~+8��$c,���d2�m纓:ay"p%���g�	,�#��j��j�f|����;<<D�\Vk�E����e'p��4����G��VӰ��U��NI?��~��N��!�e\3���m��T`RQ���1����:<�V����eި�P�l=ʠ}���E��x�$��4���x��Ǔ�q0`4)ۮW�@�P@�>A�$���V������<F����'���Dښ�9�-[���G/�&� +A7�/5�H$������.~��<��z]�_�R;���%XDj���jv״�{������y|+ݺgn(��X>�R� a8"�!�J]��`ww�L7n�@<G:�VC�V�]:�0�ﯯ)��%����]zXK�Z�z�g�Xr�����ޟ̯bz_�1$���&��V����óg�pvv��`�~�n��˵��5��-N��~�������r�X@�9������u���¼�oJ����w������y@�:a&��~�1�a,���n8v��i�6�����];���ͩx1�(�J~�?��e�� ��+����D�b�xLyU�͡�OnR@�@	��i$Q��r�$��n��3Yi���!`���39�|S����nW��K	�u�/�B	h��-�j�~������ǣG�prr��)+N�qV��E[n&�ܠ���d��+�5�t���^֯��I��J��d���5M���P(	_���Ngggx��9� VVV�I��31� R�&�揿+\>()�~�\����t:��8������4�t|��r:�V��\��v{&}�6i�f���8>>F�TB��Q��\_�t �:Qn ���Օ[g�
��]��1I�X�N��~ha��e�9���z =<�����iOL���$	�M������H;�#/F�V��n��f�/"7��x���VS�:�v��y��4��d*�B P!���!�U��)��d��>���&M$�h��2�j$-���R#K-#۝L��6� Z�v	�[��j����p+++�uzzz���3|�������qvv�(}X����n�2,N�[�-J���Ip�Hprb���ONE�fR�[uZ�
p�������h4��X,"��b:��\.#�L" �N�5������Z�kH�$��)���R�ܥ���
e�C^�,^)%�(a�t:h4���:��^�T������g>u�E�8'=�"�=��pcq�d{}v]�y�����2?��~�{Nׇɹ�ߢ�vIyV�I����M��iˠޯ���3�	��77=�]\�]j̼7('m���ƭ��R��U�N��j8���T�p�\.�s<����(
�Y"�0]���W/7wi}F?L��m�K J���	����ڬ	,����f�3��ץ��Z��p�n��F�����%P�,����~�-���k4�M����*A�չr�68E}�xZ:]�v�Cy�[!g����%��K����t7qv�f	J�:�^�n��eI��l*���1����j}�b1U������:�.R:�?R$���|9�F �'�Ɉ`��Q��tt�]�!�o�^G�\����������u�L�ٽ�}��`���^�tM�1��57��_d��/ܳ(�嵠�*���}�IeY��*��M��<O��<@�Ԍ�Cm��ޤ������l��� �@�����. ����ƍ
,���>����V�;5�R{KIZq�ZF�r3��pSM$Jg+Y�H�e�}:�ގ��,R �}haʍ�P( �� ���Ϟ=����qtt��@�t����]��_m;'ً���<�;�k�����v<N ֮��Ɯ9��,P��+="[�L�Gs=Q{:�y������3�-r S�r��ZU�ҫ��O�� ����+�\3�]�2.��m��S.�|�\\\(��R��ֿ�y[T�`�>!���'m�I��S��7�p�q��ps��,��Y�����2	I���uQX6�v�0ٜ�X�Xx�۶t�	�J퀂��臨��)Yn���r�r�����7�����fu2~u�� �L_v#E6u0(P-5���A�/[��\����� B�o�htf��.%��`����V:?T*����������G�RQ9��0VE�WM��d���A/��kϻ���x-�칼l�Vߓ���������d<�x�2�D��b��P)O����#�t��(BX��K$Qv7��uH��tr�=�G3
��@���p��O�e�`�R���������Y�=���#e,�����#խ��:h
TM�#n$��!��漅�)���w������w��,���&o���3��+���:�xu���S�s��oO^yc�(5������*Y��n��͛X__G�PP�x<F��g��v亲+��<G�Iq�䪲l@0��������~1��� ��4���\%R��!Ɍ̌y����p����IRB�A�EfFܸ��}�^{��o�.�B�&���V$r�Y]�N��H1=hf��A��É�9�1���``���V`�pXf����� 	X��uy�ⅼx�Bj���7��2��+�* ����ĭ�y�@�r���UWJ����ه69��p8�f���E$Rl��{?3���+�5�/�vǾ�f/�`~(��/W: %R��\ʌ&�K�0Q{�~���bq�hW�l�;~q��-��>f][9'7�sS�~��J�Xo��69p�]���R,;����;|�N�L�*��6���@���W1)d�I9o����t�Ȥ�B�	:��á��-�d2
�Q�|l�G$ r�|�C����e�ndI�R�N�տ�8^Lg�F1
�1�����G��F#�V�rrr"'''R�ו4� Ѹ,Sp;|Veq�� �>JԆ!�a����o�0��fUj7���l6��h��<���J$��D�|T8�
lˇ��a����Nl!I����2�}�����l>[��f_���n��X�/^ȳgϤV���sC�*���YgJ�Xo���(l�%���tr�%�[��Q'-����wu�6	��CNgw���։a�|�.�&��&�[s�*���L� |88ONN��2��d�Y��r�L&�uL&�מ�b�/.��b�|u���!��l�a��|>�J�����=?<a-��h��<;����(M`�^�˯���	t��M'6���m�u�Wum1�����	��];�Xg���c��z�l6��n�����K|L��Y���E�=�G�~�{�t_]nDÄ@�Y�3�q�dRɈ��}���r$i��K�3��ۺXg#�q�15���vl4����͹�kۦ�W��&c�&�ȫ����ܚޝ �[����2����R��+Ҿ
�1/�/烫j�y[ vS�����X�2='�/`3���0R*�DD$OH4U�S�> f� 6����q5�Ho|��EIr��惙F\\\(�e��d���I�ߗn������4�N�K�F>ĝ��7WȜ��^�S^��-x_%��ݟ^]�n׽�G�S7���	0��FC����u��ّ��m)��J��%Z��`�
�F��_�7�_��7t�e{ŨZ0���m�ߗ�|.�dR�ӆ����H�ْ�ڹ�������#i6�����>ac�κ1=v��B/��沱I�{��t����g_5&�ˠ�}?�3�*ba�킝fZ��ӈR]�I�-?�����ѻ��v66,^��^�p6�    IDAT���`i$��`�A�2X~�Nl�=��e�֪�0�����H�۽t��}$r����d���E��h4R�+;a@: ���C��?��n���ЀC?�N+� �v`7����V�I��RVa �:���^�d�k�)������M�Z��G���޺ �+�t�~��^zc��Pg� ,�;�Ne4I�דr�,�BQҙ��u�ƨ���l@���e Pvc�\�������t�,�����T�ݮ�z=��N&����y�d2�̬�jrvv&�jU�?.�jUZ���^���]nn%N���K�^�Z]�5�1��ff��ijrc�@�&{hV!ߥ����0�Ez%�i2��»}g7�@?���}�y#/c|����U6gm�٤1�* �������]'�������Mj�m7�*e;����]��X�ժt�]��\\\HeX�l6{�	K$QLg��W��0�2p#~�#�L����>�/ot��X+t���~��n���˗���si�Z��e�@ �d��K{L/k����&�n��I����O������
pk��(?1��7=7&X��Mh��TZ��4)�R.��P(,U:���cq��.u�g� �gsY���,��W]Xs��?�	&���H$"�BA�YȖ�ݮ������<�\��ϥ�h�p8\ҭ3H�M�L{�����k���J{�	 y5(:}��0/���;�<��*���Y'�������9M8���!�V�Mk\�$bæyeR�R�n`Ť�)�9��f�*�@�J��&���nbnW-���f����D�����l��R��|c��jD�d2�a���td0,}.������x^�����lb��;��(�N�S��z2���n+9�NOO���&9��r�Ml���X�y�J�~,wl�g7	2�b/�U��$��VOl�z��)X\������y���R.��\*_N@K�]ͣ�y�:�"���!X� ��O�<�H�AL_���b�`2�T��jU5����K�ە�p�ɼ֏-��*��W�eJ�X���l��/9���6�T[�u������Z�u?}T��%7-���5-r�B3�V�6A�K��gu~��vn�]���3������&�ɒ��y��0��w;����t:�t:R�V�ٳgR(d{{[�ŢܼyS��d�Y�f��L&� ��x,���R��0���?�ͤ��+��KˡD"q)M�/���m�vww���Hhx����ɉ��~4����ҮS��פ�U=7)q�ф�f�o"@�V�6��������^���D���hH�VS r�B� ;;;��_��tI��*�l�R���#�݁�����!J*��x<���өJk��<|�P�ժK��P��������8=_]^d[AQ���\r�I��u��6x�}��Zn��+���[��p~��Uް��1�)l�f/d/��ux��rmA�U.r/��I�/7�.���Fq򩴽��dpo�i��^n�jK5�L���,i�r��t�]��j���#R�T�Աt:�@)ʝ���-��8���F�Q�D#�%0,��.�9�~��<}�T���`�M���{�&e�5N�͒_0�����n�D��x�Q�W�ڸU4އ�*n�/�v0����������ei���n�%��H2�TV{��د���̐J�T��>z����g��Ҵ��}��j�����|~~.O�>�n�+�vK��u�D�p>����s�y�۵�M�<��t��Y�EN���$�b���޵7��8h��{^' �WV�\vb��T�Xvݕ\���^���9yA��Q�t|NA�m�>l�s��n�tM�d^ޖz��>���p�w�������#���^���x<�z�.�FC���|�R����Z�ʍ7dwwW
����i	Jj�F�h�����h4Rf�8��Ɍ?�������c������T�U���k�7kX����A�����*>���M�i���(�M24~2�9�׉��$��5X�ߍ�c��Y�դ�l����E�6{"��D Z�F^k�Q-�F��m���㱌�ci��*�=��^2��K��u(Ze������u�،���i��%r�� ֋<���P��+��r�sX�)N�]/W����Ѧ��4��h#�4UƮ�"v
򦃈o�[6ᗦ������� ^��|] kZ�nɄ����a��k�'Q�J��L]�(߱�.	9u!����ͪ�z��t:��/_J��R%�'O�H�RQ�Р�����X,J>�WC&:����}u����-��D�������� �����)�$u�]˛Hf���M ;/��&��M�67��j�+����M��� F�){vv&�LFr���r9I$K� �:t��TJI}��������z2�`������I�VS`R5����-���ί�F�:��9��:��Dβ'���NN?[��cob���T�ޖ^Դ�7�y6���aF����f��6����et{7�H7�����d�^��S��;��"�����+��Y�N��� J|]z`Ѓ���l4m��r*_��N���z���W��+�r|�^E"u�5�Mi6�r||,�BA5�e2I$K�� ���H���E	�2�-�^v�C��w�ӑ�t�`�D���lz�M��}���*@�\���I���8�|�Q52��,��u�h4S
��h4*�x\ML�ӒL&���fK�Pz�<b</Iz�_G�&?`?sՊe[�J��\'�3����w��8���� Ӫ[+�>�I���6n�E!����b �s�����~�7�3nY�I���fۊ�_Rs��_��	6^�@LԴ���ٗ�A�2����{n��W��6KAnҎU��|?�Z�i��y8�p��p�$��90r	�E(�b�������C��J$n�2SF��-SB���ٲn^�n�7���g�ە~�/�jU1;�x\2����^v4I(R�x�U��f�\b�g-e�k�p4�p�a�'��ƉIq�Ӧ o�q���x�Zn`�M����ͦ�k����/���n���wz�:r:����z��X,d8�d2�V������d2I�RK!�TG�á�Gc�Gj�0�����P8�����76�^Wn`Ë�s���,�!���gLL��z���D�Hr�|�B���u��VM]e��* �K���l��6�y}��dV�3��|vÆa��3kN����w��5�%��u�+��bv��S��k=��`bӚ4��.r��M��XZ.k�G��X�HD2�DcQ5�Y�:�P�)��ɗ��:�5��W-ʥ��`��Xh��τB!i4Ơ�C>�`Px��aI�Ro�x^O�L��,�41A^l�����2�M��� �U��N����)��mF�����f�Nk>�X��V��!A}�Z�7�R�{��_���f3�
3h温����6� �$����7ub�2{������9i��M?�Al]����0�J�W:�&�ٸ@��LJٌ��t�ƶ��+�����q�1��z�^�ދ��f�2�M��;-B��sS]���e�ɭ|d�z�����qj�qZ�^�@����ˎe.]95�njSӒmw�M6�μ��x�����%~��� �����ٰ2N�`�$�l��tɆ9���L8m�(�|��t�]T�6l�~m۪��㕘:�I�I�&�g����=᳝��7��M�u@�ʚ��s�x�~]~�[�����t$N���?;��g����[����_���Y�D�yM	��
���n��I�j�G�je�ou;�j w���d�l֙��T����{W��&nfh#���Uՙ]S'�SyD�T��t m��/..��/�I�&��ũr�Vf�=���?�^l�1�Qx�a`6*
����q�^��&ƌbf��LAt�� ���M�ZO�L	�*Cl�z���s{3/p����GV�TY�v�O��5J�eP&iUn�굖m츜��m[վS?K ��D"�ͅ��lu��D��U5��D���H�<4M���t|�t�/kw�Mul���/m�M�7&�O��3�u��D&�F��z����>؃�x��]kk��Dy ���� ���5��Q2�rg���)~��Qh�@0���
��{03�ۿ�m7)�W qSj�V= Lٱ���?����=�aG��T��uzO����H8��m�S�k��D ~ߒ�w������Ė������Y��1}��F�&�~@��>wz���f�2脌��n��R4�.'��<,���D��'8�����7Ӵ5��8/���k�=���u��գwc����7m�`ॹ�
D��t�L1�J��JƧO��`�� b���x��ze[�Qs��?�k`��	�rC�y������>?M/��t `�4xĉ1�-�:��u��9l�Ҩ΂�@���:AQ/;����/��,[vז)0�����-�l�~[������ZuB���_��/�֓�ϳ���*���gK�x<�Fō%V<ʘ����x��q��r��f%�Hc���1�z��^>����d���^��ĵ*�u��&:6d�� n��Wx��c�3�[������(gò�̕�$�]5CәU���T�W #�`��t:��,t�S���su8*?H�p(,��k]�d2��d"�v[:����R��ӉEe0� �����K:�&?]�6Φ'���Nxu���{��vj�4YǙ�U�67���i�_�t�W�'�}�^�����$�pk�]�@��C܏�M�f��8i(�T�k��m����u�4|o�0����1��l`��K���.��"ve�aCH����Z-9??�|��
�<s_ߋ�t���3�x�;�a�M�����u����N��lحM{n�1pb���'���tpuXN3�tb��$��%�g�N�
�$�LJ6��b�(�T����o��$�I�F�2��p����f���C���d�5�#٘�d��A��Zz������U$3~׻�ϵե�k�T*t[w~�
?���T4~����&�p�n�S���xpگ�Ƽ���c�#Z�ٖ�M��;�]�;��ֿ��I+�ǒ�+��V���l�'����: p����`rn0�3���ف?�DB_>Wp��~gB�+�87��^���Xƣˊa�ە^�'�fS�ݮ�n�,��#�ݵ�A������%�=����ņD|[x�\'Z����G�*��M1c��X&pU�N��R ���b�:w�rG=O��x�%�)����AI&�K�l6S����0_~��b����%`:��p8�n�+��@�s�ݸɊ�Z��nS�ϵ)�l�-Z�߶�щ��gk[b7�i�{ԩ�
�T�
�n��4=�,�u9�w�6H�0s��]���~��VM�l:��xU��T�l�����Z�y�:��T���6�u:�M��܆�8�~�>�N�2��ï�1�Br�&bv<�l6��g�B!5U������DԠ��h$��T��`Q�IſE�Q�f�
����l����n���hH�ѐN�#�VK�,��ƃC��J�I�5�ѴƼ�~���U@��>�s�x�Y�����5�6A�֤x%9�r��I�����U�3�:��`���ĆfF�m��ᰚ��(�J���%�N���p8T���I�\��R)Ŏ�q 
I"�P�"�qo�����d"�^ONOO���T^Snb@ F�>�L��W�i{�a�ܘH�R�:̭M��7���N��S"k�������~h{�[�d���t-�f6[����R?��t�@�@:��2D��p�Цq�.s�秿�Med�
��|�O\ү�kM��;Y�osn"��b�[~��)�H�X�R�$�RI2����j! #F#�:�τB��W����� &��f2���P@8�J8�H8"��\(�VK�����u��j�h4���L$91�NĆ�>߯��aC<���z�}�Ze\g���\�����}1���16 ���YϴP��%�I���H$TiF�~`�@n8V��K��
�cZV��W��h4Z*;���g��s����>YR
���� ��ȖG���C����2�A@�		��r�mb��:��H���5��ƴ��]��[��6�9�s�d��w�����ƺ����=8��K�́ߴ�߭�Oc�Ӕ�MT>tS�U@����ܶS6M��ٲd~�&8��X��~��r��[���Y�D"���%���R�T�P((����bgLcV�eq���A�L&�����v2�H��Q��!b���Auvd2)�R.���lJ�Z���S��F���3&��`��U���r����7��G���a2� \�ɍj_~���}XW/i�=�2=X�d2��	��{�41��X,J�PP�Ll<Q�u<]�Ѩ� ��:{�ׂ�CƏ����c��bt��
��f���h(�;���b�s7������1���C�A�����f*� lA�����6�Nr��m
�	,���;��Z/��q�����H^e��Es2�wKllK�:[�f����aٔ[�M�Mg���6A*�Zd�߇�^���f�A*�R�<��,WO�����ޞ���H2�T$���GL�
�ԙ�z<���s�3�8[b����c�[�N�ekkK����svv&����l6e0���]0�!�/гqU�
pk��t��1թ�������n�������>�U:7���N9��#�M&��N��&ef��x/0��lV��B����u0��(���b���A��X��F���m\� lQ^8���������U�T�b�(����j���jI��Q_^ ��p(�NG���~gjۚ��_�!n��Ϛ�5�  <m����ToBs���C�:�'�A�6��i?8�P�k���rrX�;��+�u��N��]cܘc��w6��vbBm�m�7��mӔv��X�|���p��p�-J.��|>���y�"�>�%�dRvwwe_����R)���N�KC| ���=#:ӋX3T��d2�R��_�2����4�M	�J:�J��֖bv�����B�0%�F8�w<K�ߗ~��4�~����X��2�X_z%�^�_�}���o9���d��n�o*#��>���|=�Hd	�F�Q ��X�J�T���֖lmm��Ei�W��Q��D"���>�88����ql���1��<��p��Ey	ݴ�bQ�����H�Z���s�v�����ǟH$"�Vk)`z��Wes�8 M]f�v9^��W���].�.��n�L`F�i^�8p��p�R/�2�&}��2Y�py�Đ�\ܘ]/��t�N�pqK�7���5�y�����}��M�ĭo���%;��f���u�&��h��uO��b�nܒ4"��y��ݕr�,�HD�a���R.�s	�Z�k ��b���q���`0�{�r],�m!�H(��K�w����p8�V�%�\NR��D"�f��DTO����d2�F�rzz�@,�.&�����6�:���~��_����&�n�=���N�.d��(W}��{���NC�\"�{Nml�^b�Ø�
�욽��b�P($�RI����X,J.�S�TDT92�����`0x�� w�L�^�l���iF�� ����r��f:�3 �'�I9>>V��K���x\���>���v�
�y�#�"$&�+��}�mY��&Ь��[�nS^קә<��`��Ynj 3M2���T��e76�+���i�01b����J�[�G/��M�V��ƺ�P/����m<�W�맄k3���Xӄ<�u��qs�>nS 9F��qn+���r9����n���#��p2@< {���׃��9�:3����^�D45�52%��I:�VRH����~�dRj�5���q�îC����c:{lu��?M�6>�n�i�����+ap�4��R��H��ܦ��t��u�0��؆��nx��1�d���-���ٲ���s���<���,�~�#����S˃!p= "�G���L&	I����UGn(�'O�H��Q,!�d�.�+@�eS�4�8���v� ��#���}9??w����қ4pp�u���F�^N&��cf��(N�VN�����&6�I��$��mlz��9�p�跚�wl#aӍ�m>��W="���¦tk����6���]�zu�h��    IDAT��dA'��cc6����#��U{���e0(Ml6�U�;��ę P�D�Ǵ�e_uO��5=Y9�׏���!������l��`$�肕�d2R�V�Z�J��QןL&� �>��͵�V�J�����v��Ǽo^��M!n/?F?�íl�Ǡ�&�)�ǆupZЦ �ۺ��&,x�r���|>�\.';;;���-�BA�٬�b���	6�t:UY62^.�iM�R�T�X,���F&��~�܌� �����1��	R��F"I�R���s�����\.���������X` qM������A�t�@�\.K�X���m�c�D"��t�����L���������XL1���F#i6��h4��lJ8V>���*�5�É���ө2DO$�N�%��*�J0��h���8���^�$�IEnGܒ@\;0 hܫx<�3����N�������)� {����P�INX0j�pTyL��:0�S��v8����8���x]�함��-~�X'�থ��B�9O��w�f5�8�Y�1��i�q�\�vMr���b1P�Ѩ�����*v(g��B���Y���X�XǺ�F. E<s&` ��k��pN�9£�A���	�`��%I��cJ��**����:q��r9u�v:�7�7&������A�w�F�&�&��G�;5�^�D�iJ���ۃ1i�J�n,�M2�`�4{NǦ<΁;��0��!�3�h4*�bQY�@K�R?�RQ�q*���C#�7�o"Kp(��� cb�Y6�4��3q�� 4~�TZn޼��c�?�^���k{{[e�NGs� �l��mSf� l���T�oooO�Ţb9:����������|�R�����d�٥@d<K�ݖf��@��ޞ��e&{��� �d4���af��P(H�PPq��������d2�������rzz� :��X;��\5``����@�	�aࠁټn �%$4��3��gS��[��!BB�J�.9rZ; ∑���đ5ֳ�L�ַ�m�,b������6ڒ^�\~+���ֆv�o�S��R�&K���M״I����N�ewwW�+��>p%�$���m�a�`�c��ѫ0X�w��[ �c�i�D"�D�p?�����b1�bC������ӧ���e�X(bu���{{�D��:b���[��Nl��I���rc�7
pW�n��U�ܶރ6�*/M����m ;h� �����N�R���'GGGR�\���Ѩڬ�p����>#����d2Y�XvL����� �"���:&�3���(�ڈF��J^~w�3z���a��5õZm�}�Y���@/]*�����ꙠI#��*W��x���4�Mi�Zʎ'�N�&;'�[�TT n�^�v��lmt�J$1��PHj�h��FJ^���%�LF%gggR,���L����s��K&��X,�Z��˗/�V���&�C�wX�����ޞT*ň��e��">\M��������5���	���z������$ ��׉/�~�//_��j�*��d���8\Տy�*��LdUY���ՍIv�_��e����ٌ�u�Y�̈́Ϝ\.'�rYI���"@*G�[�2 �=�ɩA��'�Y<9-H8V��}}�&����qu|�2�Ƶ`�@2���@@2�����駟[�vhr1!�d{�d�/&���o���u{xlbߪ�����m�� �:bW]~�-:�['M�`��yQ�����rrtt$������+�bQ��ф�T��C���+~v8*V��,|�"`��c�4c$#��~](�p`Apԟ%�88�/���eooOr��v�x\�Ţ�-�=F����m�l\L�}�-3�\N�������r��-���UZhh� R�٬��e5��2X^|�h4R]ȰP�`:�L�\.���Ă�?�2�~4��b�%�;�e:�.Ieب�P(H&����si4�n�@�w�N���?*J\?�i/�&\3�8qooݺ%~��������zM�sc꼒[�OO����6�����F2�D"r!r!K������?�,�T��@���~&g�$�W!as{���k����^6r~���	�kh�t�n�@>oB������a�ޗ�<Oct��U$��ƽ�!I;/s�!`�g��H�u�})ύg�>����p��g!��6�<(	��~�A�p� ���*	`��ך�[��$����6�_	�}���ܬ\����)��X��Ը���3����|.�bQ�ڵk�|
�Ԡ�Zxv6tH���c�� 6^`�P�B`�g@s�20��x<V�`;��c��f pG���ӗ�a>�W?�h �|>�������a ��W8e�^�8$�Ν;r��mI��KL�o0ϐ� ����Z`���f��fp��2�3�$ɍx�(���%d\���T��J.�S\�X'��D�٬��c9;;���3�KVu^L��V|��r��m)
�9�Y�j��SSy�ͪ* t��Œ�[3�hEu��>��/J��Wl�ِ��S��z��N�}����8\/-��o75�x�GSC�S��W,W/�3Τ��%L�@㌆1�[�Y��"$_<�K��B\��z�aw��y����ͱ�0ǋ��
J,[ި���%0�'�3�HF��s�H�l���x����Z-U��f�͚r/��ߡ&n}#o��O�O�[\';-�&�)ӼɅ.��bnu9̲ �	3 ����T*�J�d<K��R%j�e.3�~	A`�Y]��(��]
��C����`�e���##�����I���}8*6  Yw�T����%-2��L~�6�Y�@�M^XLk�tf�`g�[O�ں��������:�Z}�6?K$- �(�[`��yh�888�r�,�DB����6U~ް.�T*R,��M%&?#�h�%�l���5ha�vaN���+��[Wr0���-�Չ{�\��@
�cxmA�)��;��N�kr�x�	�������&� vX���	�I&��_\zg���p�\pp!���済}��@Ҫ�t7�oL<A���I��Qqg�� �̤'�8�!�K$rpp���Q�����=��jj:(��6=J6ɜ)�y� ���똇_u��i���\�J$xq������JvȄ����ڵkrxx(�RI���Z-999�n���	��C.�s�O���w�3C��wsC�D�'��De�h��f9�3p���x ��)�?��d�R�� y~~��N�)aq;���`���tȲԁ�+|�.3-x�}��c�u�&��[� ��tx����J%p�������3[g��n��h:1�����~����ɤ�5ip� ���&B��l�p�T|5�X/�	ϟ��>=ϖ�˨^$��wZe�<�9�G�bQ9�`����&dS��Zy$�����߅B��jH@�bB"�X������n����C�b)��1�����I�_/��d�l9���e<��u={�L��j��d+ˋ/�������jT����$8' w�9ɿ�`��K��8ęM��DdwwWn߾-���j"���ͦ�F#��rJG�������<���"�@0�2{HX�����Y���F��]�(���M���r9��8�� ��ry��<==}�^1f�n4ַ2�:.N��� �*��H���d�'7U�t;6 P��&P�c�3*�ٜ��s��qX�/��?X7FJ��W@p�Ϧ>�ީYI��Uu���'c��[Wg�MqĦL���l���{����q�� ���C��e{�W�Xq�5嶎��Px���ϸ��̎l���1
׈q� �l{��ū�~-�B���3�X�1��u2���|.�^O�A`��鴺�^��80�8��MF�A�=��ޑ~�����˗�F%��+���8�����?�-��>��^�ٯb�h]E�ޯ>Ô�RJ[���	��7| �Z�z�٬���4g��LF�ƍrpp �BAB����}i�Z��v�v��w�x0<e
� ����ѨL���.�L��HNNN�����6�T�<"�!H.5=��M�����tH���OH������ 9p;�Х1��������*� ��dG	�0t�����3�#��$B�$� ͥ`}��z���0�[h�x}r�`b��nG�����~�+�Y<�W�N̬�Dy��M�����D���s6ڛ�С	'�L���?;��} ��k�$���i�����N�I~G��l����ڋ�>�T4%\h�*�JR(�C4���&r��r���r-$ِ3���� 8B���Hti���r\��2�N���3Γ�h��" y��dR���J��;�����S:��$�P(�͛7U�I�^�l6��nܸ!��L~��'��g��(q������:q�mЃۚ~[r�+��ڌA�y`��unҦ �š?�ϗ��b��n�������dwwWvwwUC�}�Z-Ř�`(oD�ˌ�p8��x�tX�bQ�岄�a���R�ץ��H�VS#9��s��,�˲���X;��E��t:�����Be��go]]�]��u��}�T�Z�&�z}i,���A��s Ժ=�̜�j��0
�fLt2��T27}��h3�5�&�w��Aj3���TNNN�s{릧��l6�^�'�jUNNN���\�����q���sN��΂q��$P/����/�q�&P����gf�q�8`u	�~`Y��M��,oj�ԉ����i����x�r���$?����[�U���{�OT�
���J%U]�܅s�Ą��E"��������8����P�x��¡ �!h�%�Ù�3u\�������v,[��f���~A^X(d_�����Çr||,�dRr��lmmI�ە���%{4�ʎ�%�g➍�Ԧp�S��vmo+F����	��l�*�y�m�R���p�<ֽ�F�%+-���C�$��y#�a��[F�Ω^���
�3h!ED��:�7L���_
���E\� h�٬j����}� ����l$)�7��es4=q�MNc2��	�z�|>�J}N��9����T*��4�����V��j�xt+��σ���<y�D�����`L�.N8p`,�������3�&� KD�����t&����+��g��֛+��~�+9읋&��`�T���y^w�~��*?C ֩��y��uӞsJ�l��ʦF��Q֦�Mu�� �+ Nq��*l�鴒�%�ɥQ�6�ˤ;��a�\\\�xrI����^t꾷,g��l6�?���F������&����}��z������6�_�D�Y��&�Z�۸��M�W.�}�v��Cy�����u��ڒb����G����?7�����]5y��B�t�n\��*�����kn�/�c��;��%mH���F
�B /"j�.~���-M���	*�d`�w���evs6�I�^�j��&Y�r�+�������E$������bqo8�q��^O����cUV[xtt$7o޼d��kR=�J��^���IO,8�&.fo l����s�r3����h���x������F�L�Ϯ��ucmu)��иiCu��	L������O�������/_�g�%v����ŗ/^ʟ��g�T*��ȉ\#;N�y�!�n_"�L&�1by�	��z@�ȶaܥ��6.�'�I���R	�b��~��� 3��hTi3��4��%��U@�&�h��4Ml������M,�����X榩�o���Ʃ��4����?����$��z���s��D"�DcQ%�`�.��P(t_D�N&�A��j�����ץR龈H�V��l6�b:�������L��tz���LYw��F
��"�ܣt:�l.u�Zv���1���*�Z�J8�T*%�JE���4��7�M6O�*���ǭzbb���^�$
z��S�͵ݦa��ކO�&dn�[�0��J����n2`�a������t���.�b�� �q�2j*`Y���*��j5�v���o��oe:���_omm��":CC�`�뭭��N�꧟~��l6�����C��bgg�P(tL�`0��/_�d2���m��o~#;;;R�Td{{[�w��V����*E��c��ݲ`n� ܻݮ%��u�N]̺��>���F�{d2�H�ەj�*������&0fh���q	�+X��Y��e2�g���ć���5���n�+�?��Q����n��C�����ih�g����-�����K�PPC�/Y%(�Y\,��XF��A�b����5��~DYU�ˁ>�Z���I{~"i	�BR(����rxx�ʧ��zB��k�Ǧ:�$�Q�Wyй�}��~3��^5Voj���fr�j]~ �k"�k@{�Ǭ��WP8	�&?���y������r!O��u`O�rW��F��F�����ݷ�?�r������f��f�3���G�ѽf��F_�!;��)�$��^o���k$�l�����8�׮]�N�#Ϟ=�Z��F g�Y)������0�����s��um3�m��^��ݜ�2�Sw�͔�u��%�A��@��`b2����i	���3z<t��E5�M$���C�t�)-!�	@ӊ�9s��+�8`�
�o��䷇����޻>�`)�����q<�����`��ŋ/...���T�Im��$�N+�1�V����4�e{6�fp��³I$���fY?`����%&`�`w�T�k�������_�"O�<Q���H$�4U����\�2z5��P�דO�)>�n ���VV����l6���/�ft�f����f�V���s��`�������l��*���Bf�ףwٟ�!;6�d1��tv�PX����vl����ɉ����G}$����MɈn�� Dg=M%�� �6��T�4%J�8�,�ަd�Y.�Ĕ\��O��{�$R�d2���~�YJ�v��R��VXuE�Qw��#a��δ�"�u*��D�Q�̮�*
�E�~������}�D��B�b�x�ٳgrvv&�jU%�h6��&|lS�Ԓ<��iG�1'�I>����]5���J�T�t:-���2��ŋK�u���0�ĉ�5U����7�t��ِ^&۶��	�Ӊi6M���	:$�fh�������;��DG=�N�������T��x\r���.���)�0�L����\�~]����B��M.���������[�RY���/���ݻw����N����2�L�5y%}R3	z3~���0+�&L;�v�ǔ(�H 5э����ө4y����������K�7`Xp� �r�����4�٩L��<3g�s��4�HP=���90�u��P��W@Z���Zq�<�¡�0�^es~o�[Wg�y߳N�=.�)���X^�|��{.�[��?��x����نm�&&�U�V�n��n�4�&1}��H��s��˦��N�����֌cb��}��r"�d�m���Q*���C���Vk��m�$K G@� Ī���E(��-�J=H&�(�J��.���9>>�f8~�N�?��r���si�Z�yE����Bه�hz�1�s`�`����\./=�l6+�`P�á4�ME^�$:���}�&�ӭ������5�u
Z6e?�|6���=��亽�T\R{�2%-t_f2���F�8_7�f�/7�  ��a��6�M�t:����w���T*���L�l6��7�_������Ϟ=��|>��^���/^�������D>��C�v�
�8��,"�2C��E��R �Bk7
x�8}p r���"3��fS^�|)���rzz�@�ȥG����ଵ��t.��*,z3���ǘ${br��o�f����`^fu$~o�e��tV�%X/<��.7{�gq�w�<"Q�O��Yh�3��j8����4�v�ʦ��͛��T=�Q�X�kOgoݦ���H��	���Iʇ�S���֍,�����A��Q�~H/?e�����)�k!�����F%�X�RIR���&�!*�裃`�?[�[�oP�Jg���$��I.���J����b�^%��_j��"����|:�Ͽ�B����0��;WX�'�c�o�p���q)�JK�h���q�e
�}�S�mrhy������m�U�6��z]�[F���L֊/W    IDAT��������@��U��!��н�0,X��Ћ�}�$��`x�Y�ѐf�)'''""���N�������on޼�����}y��W������r��U8���l���/��\���$�N��ё��"�
�gV>�l:��)Gf_���6`N�p8�n��<����g	����~_i��y3�d��$	�L<_�Y�B�L$%
�5@ǉXA���^a�e��52���q�x��'��>a�zXc�\�S.Q㞳�]F2�-�����zЛ���@����i�)�-��zb��@�Xpvv&>�B� �rYr��Zc{�oD94}�*�$�r��9��6����41έm��Z6�+�nq�_��5�\���w����^ӿ!A�Z����.�F]s����W�T��\� �&�I�q J>��`0x?�|�N��5��~�f��o���P(|�l6?�V�R�V�T*�����J%ei�D���Y�<K�q���#��\��Τ�l�L�tZ�Ţ�ř�]ܚ(�
�ms�*x7lwv`n�kܫ��KM&�j�qNf�^���o��7��9���lLP����f%��)���3��zY9�J*�Re}l�v��<mg��|��gr����R�}��y��O?��A������U��?���<�\B��loo�{�����T�ͦ�W�k̢q���[1���f3�x����vY���� [,	�fVU���~M}삡k9yD&@_>�WN<�g8��k=g,S��P)�����y�v[:���>b�XG$ ���\ټ����랤�<Q�W���������"�J���`��3':�Iy�K3��:���HB��j��X+HP ��yqq�4��m�D��f:Kn���U��g�dWN�M�8{��v��T�������>ӏ��<��{���u�l����'�NK&��l6�J�ا&���@�0�՚D� �� �-�o��f�����N�~������ŋ/��Ͽ
�B�?~�Xf������*M�|�ź!����A��}5�SD��!�����������mbR�_k�M��~�/�*��cOa�^l�Is��^Y�U�R_5���BE��,[qi�}a��́�n���BA>��S9::z��f�|����RNOO��N����������^�Z��t*׎�I:����m��j�! v}���ӟ'� ���l"|��!1q����2]��[y��s�+����'GGGR(��&��đH$T�ź���6s0H�ӑ�p(�~_�tFs#l���s����T���z]�k͍^ �pD�@R q�/n�<�!���dR��ښ������Mw&'�o�+��+/\V���ǥP(H�P�T*����B��#h��ְ�&N�˺䀫$�����ɍæ���P�+ n�u~ӫ�:�=N�A [X@B{���-�rY���L���$��vz��R�1�J _��������f%�H<��b_�O������=��ڵk_����>|(>���=�b""*�tZ�&'�"؇�E���n�U��*!�ԆS���^��w�X���:��<������,�2զA�߇Ǭ"o�Ā�4� ����e<K�ەH$"��DIF����m��z���巿��ܼy�A�T��ڵk�U���ٹ/"���ξn4_M&��[���Si�D#ʾ&�`�m��A[7#gFV�Q1�q:��``���y)]ˇ-�w��rR�T���@������Pr��@g�_x���s��h������c�ەZ����3����� �8�)�+@C�ד��Su��r��{�G�br�氏$�05z��G��w|���}l9��kէ��g�On:�cF��c��<^	/�T*�&
b*���	��0�קҹ�݀#'�NL00�g�3�uvܴǜ��l5�] �s5�����:a��iJ����Q�6�)����E���֖���|i� 9G<�*I&���X(Pˉ2�,�O�R����o+��{n�s�΃gϞ}�F�Z,�������|�R����J%ł������XO�� �T*�|>�N�#���2���l6+�~_���A�˞r��1xS/�D��xl?�"/�e�'ë|�m�_]�M�K��u+]]uc���� �2#�l;�y]>��	�'��� >`�p\�_�{NNN���T�����>�>��A�Px��-����<z���r���`0���z"��P��*��$	j1����4�u��*��\NiV�5u���v4��t�gf��`�A? ��q8K�R���+ׯ_W>�h���k�
_�xc�rI�������T�U9==U�,�t3w��H$��@�.h�:��ɶ<�PH����,��`2��X,d0(�1Xc�!�I|?HU�sh��k����X`j�d�/3�����7���B�ɤ��[��/�-����AN�S���tɃ�1������Y��U�4E7��m��ۋ��,��nxN�|��pN�7[?O6{��Gg��L�=�[(T��>�I�~8�^�h$*���$�>��`��|>�Í7��3�_GGGNOO�����JD>���,�z]��д�����@�$	��rJ[�"�;���M(��2/��Xm�8 y__a����`em�%^��oV�I�����!�+�0��|^����8D��=�4ԇ�o{{[vvv����lJ8��?�X�_���T*}y����>�ܹs����ɗ�`�^���O?�$�^O����\.K:�V�4q8V�������}��(��XC��H�`(��Ǚ6�IP����x<.;;;r��59::���})��2���h���dD䲑m4��?Cߐ=������S�����X:��Ҏ���K^x�]���b��P0�����8L٫�,�b�P>����VE�3`�0��W�Nqf�"^�݁``���4$�؃ �	�|1W��O ��Ž�1�pA@�:k0���s`ⱖ�]�4���+K`�M�D ��D0{��ev��9�IL&��<t��`�`����o�]gm*t�\�e�Ԉ��b�9�$�ƉbC:�V��)$h�|ʿ_[�|�s�D#*���{;���O~����NNN����_M&�ϟ>}*�ZM�2d�Y�*��v=!�~bR
��
��R�^2��n�+�FC%ٺ_���ȭ��*���R����~7�����Sg>���7�����9w�����X,J6�U��-���:�q���`XB�V�v�-�DBnݺ%{{{���/��U�T<y���D"�U���VZ�|^������$1�Kg�8������I*�R%s���Vጞ�亯!��u��tZ����ƍ�����d��e1]vO��o������&�����ȏ?�(O�>�G���ɉ�"�av�U�d2�^�'�v[\|$	�����  ��6�)�-�^�y��$���Ϟ�Zw��DCPp���RxY�9��#�ͣ����L��FQ=> ��%���	��Pvip��\� �s�J�����`����T�{|_$2l����U#�`��������t:Uk��H:�Q�o����i찟R��a��|>�u��g��5@�� 7��Ʌ]l^���X��_"`�T*=z��7����?}�TB����y5����*��?G���&�m� 7+V��멵��.�O"�w�y�U���X`�Q�&�4���ݠN�ԉ��{C9�����ɽ�e�Y�:����T��.�J+:Jy�C�) 
]��XL�]�&�JEB��4��z�}�H$��{��_Zй~���?��O_F�������?.�BA*����i���q����Y�<Xc��nK*�R.N�V��2�H�'�5����� �Gs;dA�\H@���뺹@  ���b�NG������H�ZU��Д�4��4� ,�ƞ�������=�Q�&$}4�4B�f�!���Ϭ�E��d")�dB1)xq��\.+��
�"�H�2� 0�H$�\.����
�d��v���~�/�z]�ժ4ա�
�d>�+ 93�Q��x�j���m��d2)�����G�ݻw�T*������H��S �I����Z�&�?��O�*Y	 2��Y� k^�������+�LF...���\�?�F������ź�z�y}��A�'���$��*=7K�8a&[1���:h֛�0��U��~4�í[�~q�W�?��g���6Q%�[l%yD<W��qoX���/$^�0�g׆��d��n�UXc��(NU��i
�zM��#�g���*&A�۰�kr+�9M�Y73_��5��p�{�bFu6��T:�;f@��,��ё�R)y�������h4*;;;�K������t~���=�����o���v�-ggg�冯`�PP�u49nF�ңO����R.���hH��R ��_�,� V���z9�5�:{�J�$��*M+�k$�B��� 1������h�a�FCiMwww�C�f`$��ϥV��a��J���M iQ�fX���4�{�GS3dfMu���Fs[,S>��TJ���TJ����V(�m ;L4��v�rzz*/^�Pl*�%p��ED��h(�8�Ld0H�ד~���WX��`AF��l�|˥���C����;�����?�t:�F��&$
x?v!�g��e'��t*�jU��ӧ����˳gϔ��4��)a��Ž��E")�˲��#7nܐ۷o���r�9??����/���cy�䉺�  ؞�f� u��[̩���}"����-��U���lAgjt剄H��ɤ1�N�%���*N}���b���ۿ��7�p���?�,�ZM%J�\N�����>������@p`�9� �D�m�SS��]����;����0'��0��ʬ6�����/���z雬��n��k�*���ˬ7E�Q5���5;��p��s����%�K�V���^NNN�����egg��_2��kgg��p8���ONN$��͛7��dǽ^O�J�גn��af� fɁi"�6�+���k�A	�1�:���`��D#��zPf� ���`��-��n��W]�Ћ\�Sn�ġ����������#X\�/ ,�I��pL�_��pbs�h4*�ZM���JE�٬bc!���D"��fewwW�����k[8�����3�/��xD��ٙ�z=Ő�|�RR��Rs"�� ���c��U��%�����������ۿ��?�X���Ur�F:8I	t�����-�T�Ҳ�w��ɉ�>�x�>��c'
�j�`P�����͛r�����O�ƍ�$�ճ����6��Ty�ˤ9Y�y%)&��=�� �g
\u���,C�����yZ�ەN�I��d2���J^�o��������F�ޏ?�(�BAvvv�W5w<)1{���!����j����D�٬zV���M�[�6����*�m]�2�*�3 ���R�S�0Z�4�nv=�^E����_��Z��2�HJ8^����A4�0s�r�`0���N=z$�nݒ�?�X*�J��pvww�?|���P(�ϝN�ޓ'O$����֖�l��Y$��ܢT���� ��t:-���K��[b�֛�t|&w���T&���~x�&�O��u�����R��dR~,��{���zh�ӳDD�� ���5�F���j�ҫ�;��2�eP�׋�0�r8>�,[��}��목�'2(�}�����|���p�Ё��{�m>�o>�_� ���=��f�I�����H>��3�������J��^�Ҝ�"H�����E��www�T*I�T��Q~��Gy����e޻x�^ ����$����,���o��?��w�J�X\j��&e��x,>|c���o�ɦ�@�#�!aCR�	���vMh�L&�J�yK$��mO¼�W�R��_��_�
�{�HX����ɳ�������	���KD��u�|ۯ8���^�΍p�3�����pk����u�&u��o�&�o�Sb��jQ�ꔏM-"��{,*4���q	��Φ�J$K�w�$ ��eٺ^��_��؅�q{{���t������w�>������S�Խ~�/���""K��V(�1���-ָ	�� �L����ϛK��Ee[)0r6��?3r,K�p����a�(��ѐ��dT�r4)Y�~�`3����}�N����x{��P� �O��xt8\ ����.x��c�� ��t:�V����l&�\N�ᰒ�`�I��Vp�o8�á�C^G�Z�&����n�S��\����[���$	�~�������|��GR�TԳ�'�yI����\��f�.A���dkkKJ���"W��%���%�H$�����=��O� �rY�,�_.��\.���F�!�z]���\�֭���(���ޢ�b�19�[�k dRh2�D"��������+�N�N��Wٻ7�T�6�M�tZ2�:�Q�a��h³٬4�M�p�	��\��F��Pok� ���:��fp� ���%y�7E�ii~���[��D5�V�Ѥ��hs [6�ϖ��11����\����ٳg�h4�Ν;�L&��}����k:��ۑP(�|[G��
�J��evV�<{���� ���5�$G	D��Q�a�kA�R�N\���R>x�u0�����ƛA>3��͆~��n�l6S�E�l��������J�����j����\.';;;���-�hT������˗/�
���� ~�l X���o�P���5����(�f3��Q�T�X,J8�x"�F�����--��2���t8<]����Y`3)� 8�9���N������Ju�� �I�c�C�-�_�	,5)�B!y��<�\��J�8�a��P($;;;r��m�����K6�]��F�9�����I�R�B� �z�J��&�&�3����dR���F#ՠj:�9ư2��L&5�F�sppp��v�ܹs��_���o��=�@R�Jj2���b�F3'L� �M&��h4d4)�$ ~��C���l� n?g����������NY�����W�\x�0��^ ״@��;ꓗ�F .�����Y8�Wv�}+�v�-�~_�٬ܺuKnݺ�_�+�J}~?�?�駟d:�*-@�~0�!FgQٖ	(���1�w� ʶ_�L�Tx�	�{�♣�����5�Q�����	<n�j<W@NhD�u�oV��I&�R�T��>���CY,R��d8�ӧOU�\�X�7nȝ;w���PR��y���b1y�왺&n�ĚG�W*�RefXO�Z�%4':C�F�X,��֖��eŖ��n8J�ݖ�h$�VK�ժ�x�B5��E��A�D9ZZө�C� zhh�(`z$����N�5�^ ������H9�O.�u�7F����;{&w��K���%�y�JZ�����*)K4�;�ĩ[�n�o�[��o~#�oߖX,�d��R��|.�VK��xN��B����&+����{�{�0�_ CB�B��X�c����	�����J{�������t:��D"�~��g)��rpp�<�%���\ױ�R<b���d���Wr��ztj��W�g�����n�ˋE6]��Ifn ���ez��M]��ll�t�M�L�
$َ��o���@�ٶ�D^�6�hK$��tDD��?�����b��_i���l6�|���?/�{��L5��Ws8�l:[�\q�riXDT�7�;,��^��b�����'T(M1{�k�t�|2���W��f�X��H$ (½@�{��dd��%�B^���b�t����ڒ��C5�?�����nݒ�>�Hnݺ%���J�
�74]񁌆���}�s����(��g0��ŋR��u��@a
�6@��{��K�ՒgϞ)����s�["�PSʐ`�dH^�F����1U��:\^����ϛ�u>�M��^��5����_0��{��|��b^��|�����O?��a�5~oooOn߾-w�ޕ��#�f����c���xjx�&�I%�kl��j�Q?�le&6/��}#A����2�2���%�m4a�|�k���r�|����߿N�R�`G	����l.	,9'��-W8¡��zi��ep�\:l���a�	[bӏf}c[���1�    IDATbM,���2[�47э�����&�6ٮ�å2�@Ah���\�k�K̰Y,��f��H$��[�n���֠S(����׉D��t:�H8"�hLI<��,.	/{	��@�L�6�=��fZٶ�5l^��mʟ�fQ p�w�(cJ��L�0~��Kh��X4&��e9 `S��b1)�J�C���|>�|>/;;;r��M���$��+fVZ|����t:2�$�J����ܽ{Wn߾-׮]S�˶ZpA��,���(]�%�䠌�c��Js�
i� F^k�0�a {�pd�Y1s�;fpe@�����I���N��g�%�8�7.�r�H$��'�����L&#�\N��\\\(�v�ٔ^��$��:��ّ��9<<T]��=�� ����x\��5�)"e�2�~�^\\(93�<hCg	Y��؇��D�D-")�ȯ����#�\Nɭg��C�/�E��p(|�wھS�7R��|�q\?���$��}[/79��L�7��-�;\�#6�T}Ӻu��
&��'@�YDn�.<lѽ�``~��]dЁ@@�˚ͦD�Q988}��'���S.���pX����8��d�,���������@����z��8��(�	�[[��%�=�裏����E.��w�h|��r
��F�%�9�P��ԧ������c����4��%�I��#"Q�M�R��Q��nW���\�D"
b �&P.��ڒ�ׯ���ץP(����q�\���}y�왼|�R�ݮ���ȧ�~*�}��*���.p�X�/=e���P�fC�7�j��/\;ۑ�'8�\���]��%����7�N+�z1_�t���ƺ` �7(��Z�iy���Ib�~���9Ͽ�l=��e���8!��w������iIv�w䣏>�n�+�z]=z$�v[%x�hT����Ν;��'���ޞD"� ���M��pm�N�ɅbM�����߭,ms�p��a|� L!I�������ٷ��>��ǿ���5�X��d2�|���^�x!�fS�����1Y\�I$���~Y��g�B$�H4����{2���䟟��m5�o�eR��"b/m��/͑[@11�6f�~��*���ߙ�,<e
�`,S�J���:��c�M{㺲��]�<�΃$[V'�N:���m���9?���Џ�� � �Н ��mY-��T�y�Y��ZG��νu���n�% X�Ȫ������k��6@�OR�σ��Ec<����C:�D���z���ȣG�Ԉ��x,2q��o�w�����`�Me,A���ZP>P ����d{{[���u����dc�Z5|�ۊ!z9���]���`�.[t�t�������l4}�IkuuU���nW��B!�Fjz r6�U#��keM2f�G�Q�"��d�Y5���I��P޽�x�^I�R���&�xB��ܳ`P���-�H�IӇ�����T��������	�6i�fEe���(���rt���U����4�k	%�폩��2+��tk#Sb��\�l�ㅹ�0��91�9�ͤ�i�%��tZ666d}}]r��T�U��H���ewwW2��b%M>z?{^���5�˂��xvvn�6L��Yg	�K\s�
\}��Z�i�w0��p���0��|�C?k�޽��o�ۇ�|^�ͦD�Q���2���8��N�� YE���XT&xX�SY����JK�}��j��䮎%
V۩�Tbs����a�ɚ�惛��M����)a㰉>�6 �P8$�z�_2�̿�Y������n�A�V��V	�C"3y�R�A�i��H�p8��;1p�ln��?c��h 0��g&����ر@������z0�3�\:#<��> !��D ��p8��j�ח��=g��C90�ä�x<��`�J���j�j�F��F��~�f�j�.��x���@�u�\vדv/�q�hi�ZR(��n�g��4��C�������^�WI.LC^hd�30�2'3� ,�6�TٵN�\�z]I0 ���{�3�ht� ��=9��O-��l6+����l6�^������q�������}?*�F�`;��m�ޖ彎��b�?3��5O."gX����S��@ ����+�q��T�����6{8�R3$Ltq����M��N��������N]����M}��4�7��y#���u*ep�i��6x�����%�`0(^�W5�T����^�����NNN�� 	���d�%!v��L���jZ�1�̒�Y�ӡ��էP��8�r���k�G`���q{��z�<��ƺ�~���އK���7����#��X�ͦ�9��C&�e;�W$��2V 7�HH$��` �|^.���r��\.����e:�J*��{��&1|F\/XF>�tOW��6qXq�9 ���t*�FC]#�#3�`����;��  �2���0�G���9 h$>�C~�9B��J�x0O��۞�����DJ���{r�KٱXL�񸬬�H*��t:��'�G�6��HX]����9Y�n��}��(�m��a)���V�;'�mV�?'g�������?��졍=�q�+D�/�`Pi�}>��A��'_�����Úc�I�$!.�̦o6��:�g�SJ�q�8>C��u*7��4�ݔ�vi��..�]��E��v7�
�ZeSvZd�L�%$f�d�����l�K�n�[���t����%�H0��s	 �~�-r���14�0��CDD����q����;2�6S�z�J�`���t�]%]@ C)��jd`@."W����jL���o Wf~�`�Ὂ��F�j�d<K��R>� F�k��R@�����$�#$hVk�Zrzz*�RY&��TkU9>>~��W`ƹ	�$m��.�r�}� �<���h4pH��� 	�֍�z�DC���<<Ɍ׼)���ק�=��`M ���~qq!O�>�/^�����áZ��tZvvvT� �����>�d2)[[[R�V���BJ���l�d$� x~,Cҽ�����*��>��Ǳ�	�����$s��窎���l*����o�/3�88�K�J�����{���5<AU=u�=^��oy��]�+)�l�F�&�l.//U���4o�������	N�w���ӑ���´1iE�M��pi��:�MF܅�C�=}�"3n"W�6�LF�ߗ/���p0�<�%n�)��{N(���@7C�G_^^J�T�|>/�����TP��� r`�=�X+
���R�t�u�eԹ{<׼����
��Y�NGJ��T�U�u{
� �u�]%W�}�L&2�L��ÛH$��j����HJ��D�QU�O��
��<R_5u���Vp/H$꾷Z-�`�Y�Fa�prF��X�U̖s�����������
=.9�C��f0�����?G��ᒩI.er�` ��t�X,���z_T<�f�KFyeeE>��#���f��~#����	p�������+���J`�y��%�W'�=��\���u��MS3�}�N��dm�� r�i8J�ՒP($�Z��_��_~���5�@��>�K�VM��5�+����8�焟�$��&&vI������cp����ҁ���{قht��*�Y5�p#��ĉ�P�e�6ʨ�^�)�R������a 8 ��iN�(���Q���Y�j��"��k�j5��󲻻+�lV��38���� �����, ���0 xbV�N������h��&ʙ(�W�U)�R�T���(���3 ��9�����2�L�^��˗/�ɓ'��d����a�5C_��t�F��|>I$��%�+��e�Y��[�6M�B�>{�r#�&��/0�jΤ7驁�`P}.���?#ޟ-�`3 mU
d��%݃Y�_�����N{���a~yy)�VKMþ�w�lll(�ʟ�� '`��b;�v�-�Xl�a���c�Ղ����*���a�}��[����"}JK6�W���P�z=�3�7��W����`�s��{����ت�w{�5��l:����sl;Y�-�K��Z�t���UV2����/��:�v��~' �D7;�:�
N�Og1�4M�y�V�N5.4\� ·�+���ᆣ�l����}�>�@ �f?[Hx8����O�^�����F��nK�\�J�"�VK��l��2����@?p� �?�DB���@B�엮-d�)�2MB�u�`o���4�MU������أ�,��*�r||,�GiN;�����ݰ��Ca	����5w�]�L&jֻ��������s��a!��,^�|�%�~�՘O�{�i�8���D�F�zC�$ �XL"���;�F}d��ݷ�ҟ�l6S>����#y�f$4.�K���N�r8�Gl���F�!�jUM���k��ďE��ǎ[�y���tp��ybz=�s�ʒL�z�Z�X���4��O_�L���x�v�P�

₈��3���.��	#3���=�kN ���VI��p�E ��?���u�X�
�^g8â�S���1��pY��9�|d�������(�<�@�!���x<>F�1k�C��n?��?���ާ���M3lc�L9���~�`* ��"�f�`��~ B � <�n�[|^�*ꟑA�θ��	Me>�O�.��ʀ�-��z,�Г1�ԇ&��Cl"��"�f�����K��t�7�%�JI*���}5�}��j55"��Pc�`�
�[fjQE������;� >�
<�ˏ�w�����&P&I�n8��҅F�5�zR���Uv�
���;��P(�����m��ܔX,�$�t����V�%���""�j�duuU2��d�Y���ܰdD,e@Bl7ʊ%��Y�ϰ|�$E�ڡ��E�<�H����^�5�/�ɍ�CTާ/���{猈���&ON�|�L'sx�{E0"}6���,����S�+r����s�3�k�E��:@sٛ�`�	ȵ����~L܎Q�KQ���^1�<��b��[h`¡�N��������k0T��z75:O�B�P�n��X�0�:�Nn��r�vn�Ih6��Gb["]f�� ��������čj��,�u��I>��Ұ�ws%@�K�
���S����?P����%��J&�q�KE)����9>>V�	8��c��g��f��n����ج� �A��Ɖ���&U�Z1`ź�Xa.��R��mS��&�h��tG�9����j��0}Mr2��';"���o���T677euuUvvv��?�L&��(,�П'�<��ic�ݡoe��d��"�l�/p� py�3�&�R-=�gv��>@�}���fS�׫z]<Ϝ�7�A���"�/pH��i"�c����g��qw�,V����E�M _�uo���tҥ�Dj`b�t��k�nk)�g��JD|H�,z��� ��A������f���WA9,$
(��P�C]�c\�M�3��t��A7����24>7,��70���K`��=A�|��ӊ .�~���!ʏQg~���V�f�X��I �>����b�-�����\�L&����n�f�v��F¡�4�#�%�����i�
�L���^��`Yр�{�~�G�2�Z��}]V��dduuU��g'��k���Y�a�I�����l�ضN���A"��P�ŢT�U�v�����F�=������ˎՠ��kG���)�1��rx)��H(]���#���(����^�|��7����k��_ƣ��'�'wLI-�u�DW}��^�Kw�������:}#+]�Ck7�`
^����mg��7}��XS�����j蝺z�{�"v6�f �fݬ�}߾���ӻL��>�ժ��m�s�ŀ��-�A�̘��6�fq�w���z�o���L0�3�vr���%���1�e��3fLY���40�Y�)�����P�����e�
�暾��s�@+�D�n�D�v8 p�3@/|�����K���? 25ň��Y��t��,�uTwx"�N]J���ښlnn��ʊ��e�*WEh##n�0_t����|�{��(���H@�ͦ�j5����dwwW�8n��.��G�H;F�Y�rR=����\��&�1��:�d��=�����3��~���3�����;�� 9ti%��1�Er����u��M�U�k+�SO�a�e��o�.�{S��,^����Ee ���v`�*� �v��gC�1o�W��{�rK����_}���X�Eu��q�\28�A��|f�����+ �<'"`	!C0\����@���t*3�)3�\��T��W�����! I`u�=`��1��-;V�ez�x��y,5��p8�N�����/�zm�m��$O[3�ﱱ='#z��A��?Hpo"���8����`�����I �
�DI"��nW1��^��O�t��>� o��&���l�����C�qeG�I�x?}�� g�����Ϟ������Y�O���2[3����;��'�;.�Y3�n�����G��ٙ������1TLC���5�&H�1a0��������p�ګ����5W}EL�ZE��yݬ���1N% V,z���'�@�M4����Ak�I-&�{��aQ)��Ij��X_d�m
2z0d��,�	��JMfO�p����H$r�P(�����{�h6�L�B���q����d���	@�etL�`��O�,���.2�������޴��|x��+��<�����r���v�{�ca�k����v[�H��Ⱥ���4L��a7�~�RD"eu���~���ly@�t:�Z�&�F%�JI(�t:-�LF�L%vֻs�27���;�uA�,+5h��|��y�^���<31���Hbṩ3�H�S Z���L�p��l���g��W�g���ϗ����l�h��q2��, �9)ųc6�/��C8�s����+�wy8���X��VÄf2��t`r"�Bh�����s�,j�����z����F�/<ӱG�q�\���p^��S�ʘ��&|a�a����N[5�1������N%
�Fӳ��t�;z@5��e��L�Vr��+�����dl��#z9#G6ͬ��<��p8�/"����f�f���	8Y㨏��ሱ��..J�\2�]��@�l��b��~���D"�L��e�ɼ����N��n��^�K�Ւ�l�ƪB"`��̢�����Db�17ǥ�i����!+++������R��xz�����E�F��6�N���4�`����f�h8j�Zs k���H$��7�2��{�u�.p�X�Kp���Ϭ��N���9�:H�ѽ�����M�f:��C�l�ƌ/'KV1\��HX���W���K��\�&ML�w!E��N��VD�%���w�;�`�J�ە�l&����+�ʿe2���A"�WL����&G�,���Lr脀���ڻ�zab��h�\�4ɽm"�V �οﺥ�e}pMe���?�t&bW&`���p=^��j��� ��^�'�KV�r��z�0 7������>71�e3�����V�Y�����8t�jI/��Q��L��%��l�L�͝�:�
Fb8J$�d2)�Hd�R�6X�'��\�x���3�Z-��z�}666���H�ߗ��MI�RTg2�B\���á�j5I$���!�dR���k��5E���E2���2 \+F��fv�
���^�\^G��3�ziPg|�)xH:�áQ���&'mx/X���`]��e�D"��̐�pLd oW=��	i��� �& n���|۳a�sfȵbo���ϒ�������H8>�F�x_Ȕ�x<��k�c#�bPe`��nAF�M�7�@-J��!7�$�N�ś���N@�v�<nfj��Y~:�lU��b�|'@��Zu��;�Y/撫���rK�ߛk�ab:�J �T*%.�K:�������dT*�:���n��t��"��C󌮇e�6h�p_,�X����Ѐ?`�t[ n� y�I�4�HzB�3}�������&P�k.��`0�,��� ,Y/�kU�e�,5wܟj�*�jUR��bm�~�%O H���`0�p8�@+��L� ��H$"�Fc�#^� �H��
��=�    IDATI8�X��feeeE�٬�f3�V�s:ZR ��2��6��	�� �1�-��tb�[�T�z�.Jr���������23T����:o��+[[[���'�o߾�w{���?٣V7�7\$��v[j���Z-I��jmq�97�b&2OT<0����'F�Vd�hYƄ1�8�NU#!���^^�H>8��8�f�)�X�\.�뭭�4�=???8>>�_(�E!�q����F��֝���ڴ�����d��i��u4;�e�:��o-Q���{�5�X1Ǧ�2i�� pZ���^�ߗ3=,`�b����quȂii6�j2��p8,�XLf������{�h6���j�*�hTY�x<��"���L-�4�\&�i?�u�^/l���o��Q�%'k ��p��Y2�+��������񾖪 �2C��{
N �&�>'������ ��(�6�$b0�� �=�j��R�H�^��d"���'�hT�����J�����u@�6���'�'�ׂg)��(���`�l����f3��js댓��d2�.�^|���yJ����\�߁�1  ��@�Ri�ѐr�,�VK}^�/2�&pa-ƃ"tp�͌���ؐ��G����Ύ$�I��4�Tqr����4���r�T̬�몬�{��ǩ=-3O^7}:aѮ����Z�5McV�^�ݮ�]^^J<�`0��V�o�Zq2�
�a��+^�U5�V�I&�9�F�?xI�x<�������[�v��L&�,��N'�9	"{�31�!7 SkW�HE'=L��V�e�����XϛZ������Z�df�Q4��tc�������:0yW*�F;�<�9;8��(�5 �GP�@y	%��t*�z]�ݻw�\.�[6��A�z�>)���l6#����KO�� �3�oS B������YY}���D�[m)Y��=�C�U,���Z�y�=�&�Y��Y*"�!�wR�4�t:�v�J_�O����������nK�P�b�(.�KVWW�G?��d2��j\�������v-.g[1p�V�
�hT98�䃁0���F���.��Vi8J,S��H$�:�����Y5���d>�i��	�/b~�.P)	��j�s� _�Ngn���ښ|����G�ݻw%���=�A5\"����{W�@��#�1���(���2lвU͛d��n�=-�s�a�:�ҫE�$7.Qk�U%�/�k�Z^�H�8qr��*i��@��������N�37�����ӽ����������]��Z5�9fpM�\1f�gob��6��̚�NM��]t�������G�2���|�h4���K��U%���M�9n�[��x�ރ~���Ϫk����ei4����J�<��:��t͠���6O�xA�c�"�&�<���e�j�����̪�,*J_�����\�Ѕ��a]'κ2�K�\��gS���nn�[9#�ae��l6�f�)�\NNNN$��K:��P($�TJ���%��(��j����+I����T��y��'H�ȄB!��b��kRq=8а_�^$  =�N��t��s�8�z��L*�����c����\��i*y�H�b����i�,c�����HD�٬���ɽ{�䣏>���]�z�~01��nW���U����`8��x���`�8�j�
��S��k@�,�cJ`8�@^{�ە�d2���V)!#����m�^�p8���V*�)*�prq�1�����1�� E�Ѩ�4�9a��.֓UU���؍�^��5�Op"��sKipM���o�B�3V+�kb�בS8e�X3�e!t��Ie���2,3�PH���j5i���h4F?��S�V��fs���n��`3Y��>�Ċ��ǧ��TSn��/�>��^7��1�e�-��B�`��zE\W�z�.�bq���cb��e��x�*�����Y�׫�;�������K&�+]��ɉ���H�ZU6:(ׯ��J4�;w���v�='� Xe��]p��D��U>�yEcJ�Fu;5���������X׼fX{jJL	�����G��p=��b1Y[[���)�.(�B}��d2)[�[���+|��lllH4}�z��b�۹0���M{V`�m���3�&�`+˴w��-"Y��'�
�>�1�����gƚqv���\f���j5	�B?hI��_�����W*%����+G������x��0XΣ'+���j�z_4-։��2?g����t^K�k(�E���s��] 0�to"-��<��v�����R��`0�Zd�n�a0�6�NsW�������~�� Y��ϟ�������Q�d�<� �M<����X���m婫�L������XL5p��|��2}L,[�!ؠ,�>�TQ0�Ds	@J�ӑZ��� �����V�����V���)@Jq8���T*e��l6|yy)�jM��������%W�kO�N���P
���\.I&�""������P\.����J<���iJ�f�n�n���6V̪�w(�%�M��޳�?��IO,S%InL	�B��� l��Vq�)� W���!3x���f��ݻ�r�T�	��?���%�LJ&������ܔx<>7 ����ά�hH�^W�QV����M�������x�@c#o!V�gd6<����L�d9a�ę���p(�JE����G����?����Ιb�xpvv��J��qq���)��v��	 �U��W{�#�&X58~�@תw���w�kpMF�|��:���fK?��JLV�(vY���:��`�u�V4� ��f2����@��^����x<.�VKr���b������)���_��}L�B���+�>�췩k���Mo4��t�XGBYg�g	���;��� a=%��`�� �Z�J�\�|`���1����"0��f���s�� /�ЮT*2�L�X,�ѹ`?��4[M����i��rvv&���
P�b159����
�lllH8�;l�����rqq!�N�X�g�
eF��½c��x|�2�:� ���[Q�6���"��b��\F���~��Q�$�L�y�2�`7�E%;;�W�����0 �D"!w?�+�լb�t�hH���܃�bLq���@5%�J%��38�@*����bb:����nc��߷;�����b`I�ӑD"1����S5 �=�vkhdk6��L����������A�7���~�������J%�F���U����7(s��	�"���W���C|}W��ԕk�*ǵ\��>�y��in�"ۉE���ǟAJ���v5�ԛ�?di����ϯ���BAZ��x=^I&�����J� �(#����F���ˋ/�q~�2�v���b�����˹vtt�F�7kUْ�]���	��J����GB��� �۸��Q�Ֆ��%9�`�{�^O���r9�#�iZ�fS�����v%�˩��8޻�jI�\�N���o���˭��g���E3x S�v����K�T��` �bQ�nW�ժt:�9�6h����v�R,%�J�N~���|^�ժ4��7,��X����\4y"q�y}�	�~�/��D&���T(����]��n��o�]`�'�-�x�2������(9����m�����<�b��������f�>�1�H�g��l�p�fǶ{��s# ������a����Lg�I*h:'�ᦐ�f��؝S\̀��5��@@�ݮ�������~����y����Q�^WIw:�Vv|,eC�BB��pI�v��"������̲���Ly�ibt���ʋ>����D�Z���m7�Ճ��\�5���tu���c�bz�Eٱ]���.~��^���1����rrr"{{{���*kkkR��T��m�8У$���UiE�������裏~0��Z������ONOO�������S� ��A
����㯞����b@a��7��]�7%^��$��9bM#)@����me97	�~�����{���x��ރA%�t�]�G���ƣ��z@g�;�Y��l6��j�{£|q�� �F��F��a���\�^������X�v�Ո_x����Mm`^e&2�W��5?ɎA�>� ��� h�0Q��.V�����<؝���	<#f>M��8ԣѨ�s���,k�q�zu��x,�FCr����ש;�eݝ�T��}�5�ש�9�d."x������p0���qS��}�Y��u����rI>��/^H �����׷n��A����?8::�zz*��D"��:/��ʤ .�乡�	;�`� ~f�б� lu�ّ��IΜ��E�jQ��>���v��p���ȺF�x\��Y9;�&�포��L߳�Y��;�n4��� ���^\\ȋ/�޽{���*�LF2�����(�-%@�@� �HH�^�Z�vP*�<~�������}�)�J�F㗝Ng�Z�J(�H$27�[w6`���� R��E�EnO�2��&8	0#���_N�L�
<�@  ׉�	X�jU�_�v��qz�;@�O�x]�%����4�O��\��m� |xZy.��Un6�F�B4p��T������$�I����@b�	���W����9���l*��k���x"n�[�n����i���l6U2���,�>�c�	ܚ�'#�VK��������֖�����/[�W����	��s��س�'<4�\.���<{�LNNNԈ_�C�FPW�U���L&�6���dM�@��r�$�]���s�ns��@�lZzb�>�<�y:�J0�H$"��P���[�d2�@����j�_�ŃgϞ�kE� b1;�p��g�Mv�A#28�{4K�8fy������'t.r]Yj9�8q�r��Z�i�:�M,+|��:;G�E�Y� ���n�M���4$��ut�$���ʊ$�I%_������P֠[<::�h4�?�A�V���R��?�\<����9��#O�C��K�z��v:�����3�~��޵��C�'���e�'�V럧=�-X�`0(��X齚ͦ��m�ES#��zIhtQR��� �`���	��y�X$S�]�#�����vVXj��rq`g�p�N�2��zF��2��x�깸D���L����
m��p-�PH5��L=$�뗪|/�,b���D�!&�#�jN��^-���{HU^�|)Ϟ=�r�,�^oΏ�Dr�=C����b��d"FLL�M�WV�۲��N윬��{����R�H�ZU�;��I�_�x�z<Y]]�J�"/^��p8������[�n�QW������ן�x�Bz���|>UQ�F_�so�g2�� ��.�4r�b���5e��:Yo���N�[��jU�)��A�2����k�a��:��2�uQ9�����K�=NNN��˗��J4�d2)R�T�u�{�� pED�@ ��������Gt����OOO?���N�%�J]Y��ؕ͠W���c�.Jʋ*��3 ��$�IŦr)�� �x���m���^��^�W5G���}k�R  Cg�L3�""�DB�;���5�z��zd�3�<`�e�e�(��C0��q+�������x�L_;v�f3�x&�xx�d zd0�l_���������e�˥�kb9I`)��$BO�tF�n��Ϸ��K�^�B� ������9==�z�>�w���Tb�~����l6��jR����V��d��ܺ.��Y,H����E�M�� �Ԡ�������"[[[��x �;h�Z�O�?����	r?����R���R�쟝�I �T*���!ӝp����.G2v�U�u�̎�����}�S�aN��"��"fW���7'M���ݻ,����:р8���R�M�����9ѱ ��ְ�nK.��g�>��w�J"y"���e4I*�R  �|��Al��j�9��|�����ӿ�ۿ��:����r���bq�R�H0���	�W��t��u����:@�&�!Gii�g2�{�y `�]0�[��e!���?aP�7�1��l*��F,�pfn��$�YG+"�_%W��뱟�d���k ��B��Z�5��ѿ��5uћ��uY�q�m�ͦ�j5�Y����: �C��WY��KXx�Ak����	ց���ZvO8@�l�"��$��˜&�͟��v.���O��˗/%��+)
7��1K{ ��~�CoN23U���%M�w���:��qՙ���Ki4R*�$��(m��,�����KHJ�K�b�(ggg��ܹ�R�|��d��Λ�����/
�>}���_���D"�����R��٫
���%�7�r`���i��SًiZ�SfU��j��*�v�@o��Z�@|y��[�	��ע�]�Ĳh�Kp7QRr:�y&�u�(t�]yy�R=z���x<.�nݒH$�4���kv�����;99�n�����_~�����Gt���/NOO����k�am2�0'е�|p �d�z����Є�YL1+�70@�}p9��g4�fly�0��� XC3��!'нMx��2�Q`����$��H8V�@��@�nXӊ?8t�*�M����kЧ71����[X�z�.�\NF��r���t�æR<�O5�����s�f��X,��3J8V�%��̓�x��!��d�*X$�T*%�dR����+�w���*)��cr��5����J�P��ϟ�ӧOս�u�x�:#�g��'�DB���$��J4�c~��e}��2=�/�&m����` �z]�ժ���^����G�s >y��<~�X����yp~~������ys||�_(�����������c��ۓT*�h����X��D����\1��!z#L����AV�e�< ��[�Zf��l������. 4�7i-�J47}��[f���^�H[�L�M�W�G&~�Z��O���֖�P3xh
ҙD�h3�p��f��ă/���ӟ��gA��>�?::����H�ݮlll(	@J9 '�(������yf�i��/��Up�=G��`��b� .�| �-��V�L��	L,�D"�L�!��G#�^�8����#q�up�r
|N�����xE��יN�oz����X,J��S]� <T��,�1�`��~�J@�LF�����jgqL�K�:�ד�S6�>ߜ��>�K?(L�S���A�i҈��G��������	����l��.�t���M�V�"b�t^���	۵,)bb��L�VX��l6��lJ8~C��� ??�3�D�Q����_���'��[�n=x��姷o��^�7Ϟ=�/�JNOO��={&.�K���e{{[%H�`r����$3Cl���P(t5�V�J��ܔx���4�d:Ix��K��}@�d!k�ަ�V�`�X`
�&�oU�[������Fބl�Joh�yf��᰸\.eɔ�唟��֖�wbv �G��܇�essS���\\\�������~��7�|������o���z���^��w�]�d2���&�p��٩�S��ރXo(�����7,t ����ӏ����� �=d�,5�H���K�:�� �#Sy��LtH&0�>�L��������S��^�Wb��L�S��rrqq!�FCVL=C�쳻kJ�y�^���-*�/J6�ҋ��N0p8s^$�P(���4C��b�PJ��0�Y�/h�ao�}�F�&�u:���*��I����E{k���55������2d/H4���܈RݖM�?�r蜜�c�儒ǨZ��m�Ӂl'�q*!pzn-��9ѡ#��^�^�t:�ֻ�iD_ל���gQ��VM��@@��<z�HDd�֭[�k&7�����ϟ?����ϥ�l��ښloo���D"%��u�/vZѽ�nQU�ʊ������uf	\�.�o����M�^;�w��H�D�q��W׿�%��)8�z����C�����F%�J6�U�A���
̅B!>T�����q�����H`1��C��驸\��~���_��_>������]�y���A�������'�Je��hH"��l6+�`�f�� �l�`b#.�;	,v>���(1�M����o�^�b�(�z]5t���n�PHy��=ᇋ�	����XLVVVd}}]����&�!�B)��!`W    IDAT��v[�i6������L�ѥ)��D��3����&C~}Os	�tn�����DdwwW���d<K�\���s�*��~�F�j.<d ��c`[���R��].�\�����i��ܔ��-�d22�����L������l��kI�:�eg�q�Z�<lZ_$6�������z�.��Lb�����J6��P(4�3˞˺V4�H2�TF���\�;��ޤ�W;�J��=�����edz��l�3L�cꌷKj�H�ݖr�,�LF����A;πq������~I$�n�嫯��׻�����O��־W��Ç������|~��/��R�$�dbN>��
}�O.�%el�������u)��jr���Z�]7��Z�N=q���M�6'�'���^�lvч7Y����M�[�E��8�ZL�,N��޴�m�F�,����F#i6����K�f2�9�V�ǣ�ybL+��(=�D"��b�r��^���驴Z�����_�|��W�x���t�{a#�����z���B������j)��P(�L�].�LgS�5$r�C����|&R?��*E��n�D��`��	0�0�&m#�|>/O�<�l6+kkk��$���8�=���'�`��áJ� Bм�]�n�[��ꘞN��l6�T*�
 G4Uc�[���E�V�jr� OfzRY�a�/�:AN p���z��%�Nˇ~�Fev:��J��N�%*f7��+�	��&$C:��"���C��d�Y��ّ����|rvv&O�<��O���ٙ�7t�|x]Z9m��5�r����d����X����ONN���\r����yq�ݲ��!���Sϖ'>a�V����U���d$�H��V��tSU�G]�(e�L��{����ӳJg��S1�$�.��{N*ED9*$	�W����?�Y�s	��ȇ�!�&�p8�O�ӿ|��ٯVVV~��d�������������bq������` �X|.�¦�b��:�E��{�>Ʒ�1�bg�X�Z����k�Q��0�N��a]���9��v���	=!�^��z�M���V�$����uvϪV,)�L �P($�LFⱸ�����C0n�ۊ5C�>��"2gR�j��Z����9H&��L�����~����ͮ����J��X,�?}�T�ө��i,��!(0[ˆ�8Xqs�J���DHX2�$��gȌ1��l0��g�r�>��^���I>����C�F�2�LdccC|>�
����`�[7� (�v�w�~��/��n����|�B�� ��v+0�!b�M߳:c��FwQ����Y3��O��W�'��ښ|��r��-Y__�߯���`}qb�{L��>��x�x<.�TJɑ�����I>��B����v¤�<\M�29��&�ۓA�}~~._��<z�Ce��vK�VS׎�#��]ӌ�euuUvvvdooOI7�s���w�kHuj���(�4�\*�;���WA����zr;/x'A�Db�6�;<�WHBMͅ�X ���!��p(������F�������p8�?GGG�޹s�;?oNNN:���R�4:<<�_(�����q�h#6#~�UA��7�b��&����ys]	�wa�u�@�	v��V@���b)Qx����+��y�& �l�J�f�~�}������V�%�xL5�u:)�JR.�%��I2��͍M��2��5�0���&n�@�J��jU~����������ʃ���7���_��wt�={vP,q||�I�����r��v%�H��r��2`EP�6�%�o�p�a��*РD���N4�z҂��Sh4yL+���L�MZ��k��<��<y�D.//�Z���S�/���s���W����d����H�RQ����n�qDc�Y�)-(���vU���P�����a�F2�a�_����4�M9==U:�j�*�~_=/�&�l"A�{���r|?�n��d������DW(�����cy����y�t:o4M9�4�2���֙�g�<?��#�^O�岼|�R�?.�������q�g��$��9@���`0(kkkr��mi6�2�L���H�$X�І{� �A�YX$�c�$���L�tѳ�.��'�v��LB<��zj�C:��s �}����8���d�'��A�d2�v��ys����H$�����>����������������_6��}�n��
�duuUy��M�����-~d�Il���v�^�K�T�j��d�����:��|@�ii'��:���m�e>�ݸ�� \;�l�l�ti�)���,E/�E��ځ�B�FC5�������$���3I&�Wڶլ�F#�T*�h4(@�g<W:K" ?�x\�Ѩ��q�v�R�����ǒH$�S��/��_���[�|�D�a*�zge�B�p0��W�������Z�vprr"�~_|>����I0��t� ��z�*�@�ʥJ�Ч���*���j��y��Uʥ�{�HD�٬���֕%��`T�?�^�S.����RJ��$�I�f��D,]��� Zg�d&2��fg��c��X f���!���̱���n���pQ�	J񇇇�n�%K����%�tZ�Ţ�F#9==U	J��nwn��)qo�os�2V�#TeZ��E�ή�z�.�|^����)]��3P^�]��+���K��������|!O��%���ŋJ�!"�����1\Uև��~I&�r�Ν��X,J�۝+��F{�!\%ǯ4�H�B�p�H���5L]�p���v����#�ύs���q?8���]��k<��m및�Ѩ��jR���ɓ'���������?�D"�h4����766n��9>>>�v��s������~������� c\6�O�#fh٫�>�"!���G��������j��L������&;UY[�"&/�Ecp�9����v~�N@�2��
Ԙ��٭��� W?�0�V���̶M�\NB�������Ύ��q�s����H$"���
``�570��ĆDw���*�6�̓@ p����T*��ɓ'�Z[[��M�b�x�n�Q,?��z�BA
��T�U%� �G ��ka�`���)1?7Bx<Ռ�XF�L�ј�[�J���H$�t��~�fK&���q��V*������D���4n���P0$>�O��`e�����x��ye��~�j ��C�v�I���jb�U챒$��]H-...�Z�*m4�^����H� �`@��hA	�K�,�`�|TT0���r)'�(���������Ì��N J�þ)��R�V���f�)�BA�Ţ�B!%/��;���>��d2��$�ٳgrvv��8t�_���-���*���s�n쯬3�HB�K_YY�k�d�h��tb�u�-��*��>��������hH�RQ׌DU��Ι5�pM�e���y1%���R��&����^��=z��T*�����k�9�j����������ɓ'����`Ч�������~� �l-g"ưf�Q�XW��J%)
R����.�>�?�/���i6�ԐxY�k5ié���E����h��1��f�&�6��h$�FC�~���i4�������ϕfpssS�^���u�p`�r9)�J�h4�Ʋ��ҧ��f�^�W�ݮ�E�s<���9�v�������h4�F��P(�pmm�q�)
����`0����������`pP�V���T���*����+�{�j i*[��)�5�䌒2�}�w4���ui4*�1�tʌ�$:��	���W'&�ܝ�h4�g=�d��~8�\.�x;scru�.Պ������{�~<f�Y�>��8b�����md �L$�J�"�fS]���`������gd-"�?�{1T�	^�~k�K�˖���sV�D��sS3x�L��o�Zrqq!�����WgPy�"6ᵲ٬Z�H�...�Xr^S�@@�����ݻr��mI�ӒH$$�JI$��/�B�q#�J��۷%
)��j�����,v'�]�l���k�I��jR[�ݖ��s�][[�h4�8}Z'��gB���F�F�����q��Ţ<{�LQ�d2{{{�F�_��W���&>z|>��L&������d2�?�&H�;��������n�����|��7���K�&g2��-"s�=�&���-��ɵ��9&��E����r����Lc���/���L�t+3�����Cq2L�m^�)Vz>�����g�=�����~�/�jU�� FigmmM���S�j�d<K8�X,�J��A^^^*愁5"� i�f~���v�b��JM��������0
�q�[��N�3��r�E� ���LFy��A�=2�*1�F0� 0�;���i��aт�>��.e��Mo��狏.G�iw��O,�g�un����3��9i��'�A7�nlp�������*Y��x�-򇶳�A����1�jA��Ia()2X�d�˱s��Tf�~�Z��c=�t-�g�Kf��\�5n��[1�V�}�X'v�`[:�Y��ǅ�s�ɇ�n�E�g4���t�Od�Y5|�h��T����/�'�'��������y��dfH#���7�L�\.��ё\\\H�P��h4�n�m���y�'7��z�<�M�����U��v�-��s��Ҝ�X5b?�Ac�XQU�gk�Z��7߈��=�z�� �A	�d2��g�}�/ggg3�LP�1��nW�W��~���Q��=�<�^�����?�k\�t2Uqgv+��
)�����j��
n�\�)o�}��y+�kR����.@8�GXe�N�'L,���fa������n2�H�Ւ�h��[$Q�/��R677essSvww%�L�)S ��������󪄇$6H �����|z�˥J��RI���b��H$r��,}�-4�@����8��:��w�S�OgKq�����lllH6��ϧ\pm�A=��Z���ٙ���I�\Veh;��J��,
�d�ݖB�p��!�Ƣ*�����~" B�@̲�Xy%�F���sS9�ԩ�_��� ��Q^g�s��Lkîa�nX������:f�-��o��b��iIg˭+���4r��"���R"$�!�3z�e°6�Hr��5�l�{�{�l� 8E+���U%��|f�a�6�N%�*�A�VS��deeE>���w�|���r��-$���ހ���|>��n4�nM�H��/�׽���L��v��e�[Ĉ~�j�����T*�4��O �o\�V�V�)� �� �	)��T*%+++s	���r�H&��}c���B��X,v��v%��K��T��a��v�%�L�����k��C���(n�[�A�'$`�[`O��n�ƪIҴ�d"�jU��ϯ�m��*<������i��ۼ��@,;I�|y#��Ӏ���Tv\�s��N�[�����^>��âq�vץ{[5���:�l��hȗ_~)�DB�zЌ�f+�l#���|R(����t�\��c���z� �� �*��� ���Vgx_ ���}e���B�_8�}>��������������b����\Zµ��y%��t:o�,힫s��o�^��+�x\vww�ӡ$��~eeE"������8�'"�z9��@4%��dc
X:P���N{0�x�z��n_-�g�����tssޏe#`ex8 -���$��J�u��<0G���C]xm�	��}4y����x�<��� J8��=������m�Z�����R)W�X,ʏ�c��ٙc����cĳL&����v[��߹sG~�ӟ��,{{{�L&ED������ťw4��\.I&����iw�j:�d{��V�g���(:!����á
�9g ��� :������������݂�@�A5k��n+�����?�)w���NM�pf��#��E��n8��S`5�X3`��D6��d4)�k��j��ٙ����&f�b�+Y��i�$k���%N��c�k:���#N-+��W�D���J\��^4��J�kw� JݡPH��<}�T��~����}�⹋��R�H��Q���!q��\��+�%lZH(`{��Sl-�wjs�^_W\�G)���& 0���68Jp�(�����i@uyX(L̂�Mg'�bT.|?1J�	���P��11��@����e�̌�y�5�l�]�l���A��Z�7^V�d	��Ag]MC�*>8�p�Oo�g:�LԠ4N:���X��v
#��'���X��� 0j����t ����}��x��]	��s�b찁��7yo�=�����ݻr��]n�%���'xq�f5ِ����T*%�nݒz�����5�]G���X�Eg���hED������"��J2��p8����ёT�U�ʥ�~����R?�.�i2��k$��m0���V�Y0�����x ����6%�X/hT �����q��9�g��	^�I�h�N�ZJ�.@���t��:�Vov���N����ՊY3u�/�3��C�s[�
P�5L� q�XL<���u��/��?��#��ڒp8�vd��XLJ��x�^%�g-� ��C��f% "0��߂�
�Ug�X�g���5���Y?�{��O���D\��24��i��jr~~.�|~�L���,� Z1�hb@��Y0c�V�s�� �T*s�������E��Gq�f�;	��15ujs��޴i�4b�L8Cށ��D�7����f`��b��M{f�/�t��a�/_��:�N���۪�[�[8=��<ON�����1쭮U�f<�WL��7�*�ZlnnJ0��*�z �?�3O�Ӫ��H$��r) �Nol:y��.ՁtakkKM��v��F,C�,S�p�#��ͳ���h$�NG�F�ϧ<�!(
j}µ"���ښ���ɷ�~+�|^�� �g+8�k�O�aK2f޹��>�Pԓ���dd�.���76��#��k�b�(�\N�� � ��f�ݲ_o��}_��V �	ɺ��H�e�UZ���i:tpkǦ��4j�2�}�?�*�0�f���(����.�JE�����?��w�J&��ϯ2Ku��D�	�%0��1pd�  S�P�D d�K=A������:��<�ù�~2�H�s��=::�Ǐ��Y�׫t��RIJ���u���ꀱJ�x��s��aYYY���Y__Wc_YcȠ�9�L�|��j�̂��\��	�0�/�P��`��Ę*� ���(��;�n�v2�i�����#�oh&aQ�;h0�e&ׯKL�Ko��Y���Nn��x��Iϫ�R)Y[[S �ru �7��+���}��y��D�NG...���L�����Hq�0l#�J�q��lV�u��y#��!@�;3�qF���}}��
���k��b�='��w�PdefW1e-<��Fc��D�QŨ��m�T*rxx(�BA1�wnߑ��5�'�H�\�k�DC�n�Ʊ��Dt�
�a����SMɢ>Փ���5�{L/�'ܤ�*.�L��G��Z-)
rzz*gggR���$PV��z=�1[+��~4�5�u2@;pkǒ��s[�!�J���f���D~�D����8�1�k4)F�V�)K����'���&��k��p*�Y������]
�=]G4�L�k�a���e"t۲�:��l6SvJ~  ��6뫯�����J�n�ܻwO9R45��=-��$vI
3�ذ;�΃ px�)������b1�d2R�V`FY�5�<]L�3���TL&�v���u�H<q(���24<�~��Sc����1��'�j�!(�L��ޞ�@�����!���n&�3�l5��)�i�\gͪ�N�e�e���.v�0U(L�z0H��VOB��VO�jUr�������9��W���E��J=z$�VK�ܾͦ}[��am�{�z=�Uk�)�� h���+��u�{��o�?h�sV����+}� 9:��+bP4�s���zR,���D�����\��螄#a��ޖ�l&kkk���̀'����N���i<�F��\H�� AC��ץ~���5y�W�d&2���̮^�K�X�B� '''j���n&���{���� �T�3�Djzo�9m�r��H0o�6-*߼��[gGL�N ���p�96�G�z��0��Տ?��lln�u��/e]xΖJ��q��L��8��}X��M�g��`��2D8V�� 9V�JE...������u~R�    IDAT�Si�۲��)��L��\\\��ܚ�u� ���˫��`��f�Q��D"��dT)O����ppi���F�5� 1P��l6��t&��Ԗ���1{��xh < %;�q�Nˌ��᯺���,�آJ1�n���Ձ4y=:�o�^Y2�[x�sXPu@l��2������Z���Etm�^E2����%\TDDu��7�|#GGG�j�怷ɧ�c�\����*�W*��ڒ��-I&��ϻ�jI��W�` ?��s0��bs2 �3îD��/ѩrr"�|^�N����,j�����׮��-$�㱔J%�t��l6e:�ʷ�~+�NG���4[M���S`�tZF��t�]i4j��=,+��U�d�Č�z�p��-��qτ
˪8���2��A�P.�s�Wiޅ��uK�����:�벫x/��V�'�{�7}٩bv�d�e'*6�Ect�YDV���6��PZ�/}s��
���^�T������r�,�JEI`s#3q���L&���8L]�C�G�"+5٥Y\���7�phȤ3���.�x\�?p*�J���3��o��n��Ύ��i�*�b���&w��0�D�r�,�RI�X�ɶ] �h"��3ٯ�z�L��'Т� |6��Lf����%�v��A�D�TR�] *�[�]���%�J��Ɔ���))�*�O1k=s��#�Nu�i�sEf���1����p]�lb�um�n�ƿǟ�G;/ҋ���h�˗/���ڒh4������r99;;�z���=0j�IwakXA��m����>�@�ݮ���*�#Ns����c��r��*	>7���ˉ]�3�<;��I.��z����q��]Zk�Ub Bo;��i�CVWW��4J�R�G�I�ӑ����Hn߾-;;;��feeeE2���R)	�B""�l6�y�M�c`��.�@�39!��Ʌ�%.�x=*Y������K�V���999�\.'�FC�@��i��9^��Z��h�~Ӏݩ���k�Z��7	z���%�)�6u�.;-Ɖ��jZ�(��o��b�&���%h`���=y�D�át:���r�Ν+�b$�(�"���gggrqq!�^O�v���b�^����8h ��9Ǥe��<� ~mmM677%�͊��J��ʩ������SU.���P�>��c��,�o��E`���Pf�|�BO��`��&� �S݄_����^���*+&��ʛ#�]�Z��� Vq`�a}�&:S��J��O�[__���mI�R���rn��t�0�=��V�$���`RgaQ��j�[�G�溌�Jb�8��	>����
䢊2���\�ݮ�Z-��j���*�x\������I�PPN+�d��CӐ ���#�nW�ĥV�)�<4�b������B��z=9::RU�~�/
��G�\�&#�����+p���e������e@�)kN�����V�)���tԸs0��f7�M9??�?�P>��#���SM��&
�������c��'�P�\ћt!�⸉D��
r�e��r��9���Ekx�[�X�
!�~z\�.;��Q�
-�������2�sYI�y
VL�i�{���o�;uZ��۸̸9yH:cbwP�@Ӕ=Xe,V6b&vW��q�l�]�l�f�˭��/^��Z����?��C��ޖX,��4����q�a��9�n0�<� �q�������@�6��kW�n�������x�\.�����ɉɷ�~+�v[��p��z��A Իl�V/�#`a��j�������Rz��bAСΒ6�7u��g����}��`ݘ��@s#�I���K�S3��fox��SĠ�f�Ά��ZO`a����xX.��\��Iw\!��U��,��T\nלo'�&�;��������K8�5���ؓ���`әkL,�Jr~~����奜���1��pe�@bE:�����~i�����c%���bj�79??�z��~��L�ӑ�O�*;�j�*�XLf��ڇ�]`�t}�7D�>�Z��A`��M��랧�H��yV睾� �{���1�L��7Tj���$�����lnn�_��_��~�3�u떤�i��ܔr�,�g��j�T�������՗I� g2hDC�˃88�Z���w��ar�`0P6u����u�T*rzz*������=�&�E`Ӕ|,bڝ �E���0�V��:���p��;�=�u6ܢ	+��i��6�d�&�j�<Let���޼�;є�͕����r%�R.��`]�^�'O������=��ڒ��MI��W�ק��+++��fU	���^�]����̍eeH�80��A/kٞ6a�m���  *�J����ŋ���s9==�b�(�ZMF����~_...�:�u}��(-�1M,��l'�ɕT�\�L&�JUVI���U+]�Wn���Ʌ�M޾��e��|h����j5��+�iw��x�<�>�043ۤ��H��{�2��e���v��кZi���jp�,ɠ�F���c�͖互�P�y��	���"YU*V�~@�f�E����I��A2Y�I����dS&�23��>$��
O������з�F0q�����˗��������	���Ņ���O��ŋ��Aq�V��Fx�0N#�>??A<��^��(T������ի���\_7�����xM&��V���@��C���ռx,a�la� dl`�����[�b��V�����Ç�&�����_�*��FS.+��k���k���A�@?��">����h~rvv&���a�������C���˗��@g�b�	c��6��f�w���D��~^�(lsS9�!��y�Us�5^��g^��R/b���+8-��s��5�Y$a#�Fa!"RE�H�O�S���C���.��ߗ���7���Fn߾��%��ݻwODDB:�}Fu�R�ҁH�,�K�V�R�V�4��>�V*�Bem�\�V�4[�J%l2Ϟ=���N���?ˏ?�A>t�������ؤ��mKb���K999���}�s�N(���0�E .��x��^�?���Ϸ��k �t}Å��{N�������ip�`iA�8 �V��R�$�����k��U�T��-��"���5рr�����5gP�٠��3��R��ŋ�o��hpQ���]�_)�����#k�Zv,��H�>}*���Q���
����|��lN�oS�)�H��l��B;��Ci�Z����� Y��` /_��/^�����S�>}*<�_���r��m)�� '7���0����`�ua��co�C��gf�3�LB�{d8c O�W�^�������u|��}��5�q}_�]IZs�������Jg[d3��;,=�Lc�v�N#en_��Y�o0��5n#:k����d��g%t��>�͛7k�b_}�U0��!��޽{�������C��h�������,31R����P��H���i����_�"?���������°�" @���R:�XǯT�:�`�7�M�w�^p���K���>�j�?-M�N0��|תS�V+ݘ����d2��<��O��r�\�zg�^ �N���t�ΐ�Dj�ښ�GD�T.�Ea8�<�T��Z�`��ԣ�O* I�n�H�>{�L�={&�_�^˔�ZDaM�v��0�,�"͜��T�4��n�`�Idh��a�v�e?4(�j!x���K���zݭ1_o��j�>dT���a�n�Z��
��h4�?���rvv&<�������q����W�i�Rb�d�]����y�l�����%\6��l�ZAs����V*����"X����O���+�n��H��ꄺk�u���cye���"�:<��Xj?���^�͊c`5����:�=f͠-E
���l���W�U(@�Ç�o�����Ф���00�`QX��6X�v{��B��B�F#� p�b�C�w�~���ӟ��y��  �n� 6`]x�)-��E{z��g|.�R�$��}�-�Hh� m6r�tS�V�Q�J��%�����ق̒װ��ftu�Ǭ��|�hP����y��<y�D^�x!kU��Nʫ��1�o?~|���-��L �Y��%�0��Ǥ\��6z�oI,"��xl4���Q����Hb,<;,�g�wp�o HK#��)iO,�dM?�9�0u���g�f�>��ϭj�5(��^9��Vr\H����������������t:�����?d0ȧ�~:��� L�v����MO��tڝ���}�znԠ;�a�9�Ms�F��yyy)���Ao����5=��)ۖ�,���wp��k�T-�gSK���Y��$9��5[��T�`N5c���J��*��d�{ж�^�K��X���z0��������L�;�Ε���V��2 ��j�R�����"u�Oh�pvv&��00R�:99	��U��rTS��5K� �t�Ig`^�=�o�[��|��i(T��:.�f#�MgP���3����ֽrW-��t�p�E�g�����Zad�Z��  �����L$�v@?��_���/ y ��v��N9����f\�}������סAd9�����~� ��P�$c^�1��{M��� ��A�y��>7��9F��<dЉqB��C��z�����"���2�@(f�	v0�8�|�v�����|���q ��_݊{�x<��/_���<~�X^�x\�̏��$Vg�e��G���Vg�`�]���<M=���7�̜���i�HL_�ޡ9,tщ�5��M�S9��\���,�W-[������_m2͆��̛�ؕ�ey��U�p�����O?����P��b�z���d"��PduUY>���0����g`ڎV��4�x�"hm�={<nQ,pxx 4o���p8���� c�B��h�t�lu>|�,���B{c�o@V�)W���eb :L֘2�\�;����1^(����۪r���0`�D4�rzz*��B=z�f�W*��R����r�= @Cg%�ta�p9m��ض�=p�\K��c�"�3��"�(���r��߷���j�<E��x��:�S$ȇ��y֖��w�YM��Lii
wVDV��^�K���+��p& �����CF�:�ˠ�F���x������\^^��Ln`�kF1��F����!a>䦴���~����e�w9w���	���a��5��s3%)Щ��v�9+Uȡ���Uǈ��1���bta�?��C��j�tQ��/��x,/^��gϞI�ߗ��=i4�"Z��T*I�V��r!o޼	�F`c�岼y�&�о�4��p v��`C�=K��\�`q�c��fI��&�7�u��~��ONN�l̴��A$��@Ί�-].k���ik#�?�E뽖�T��u[M��1#��YJbd=_���~�IV�U���^ٯ�4�3�����J�4�EX~o�k������６���i�W��l��bE7������<�s���]�$h����U���&�c)������s{���l&��(�2���rxx�������e � �`Y�� �b-�� I��*��3�6$�cN�p�l���]4�lG,C��ab5�kev͚��m�s�kN"ֹ��M9�+�ʩ.���"[�s;�e���@pL���̋l0�h4
�J�ݑR���ܥ��� ?�,
 jQ��n���<�R���� @�hb���vvv�� �Gt��v�A�ӭl��2�����&���A�iV0���Z�O=�S��e���_��,����[l�����tѦ�(��A8��^S�v$R:N�v��[^��$#w?ӒO.�Qm5K��7y�ue���os���eS`O{��n����o��uU{Ԧ.�y��ަ��)v����<�x-#���~������X�1�჎��@];���?Ѩs� V�$B����F��!g@��-K�b��Z�v��S-�l"P��3e�:�r�e*���U56�w�݈��M����펖�xށ^��b��R��YO�"��2��$ f�S�	��4�V�>b�3��R"�f-o���&����XȚ�"�L�VϹO`��Q�j� Ɋ�S��u [i�����pzVv\��{Hy6�W�ZВ�� M:ou Jyݦ���a��i�Z6�g��fc٩m*�������ۦ�s�)��ǜb�]�	ؽ`)��I��Bs�+�5�}�eL�da-.�
H�������F#�@F˝88���x<u���4�D�[�<�mYU/@�5E	����^���MJ����lW�k�hixc�*<�
 r�h��M6�"zݘ8GX�M�i�^�b��j��l(�؛@��Pq&\q����A���>��vY���lD?3��xW�R ��}���c�R`&׿s[���T�^��:���׺7��y���aW7���ϴ=$�d 9�ݶ�'��He�R-4�%@r�]l�i�=��)�����j7zSߝ���Kȵ>�?$(p~��U Y�a\;� 5|f`�x��t:g�.ʼ����x"��K˅g h��J���&Ư�̀��yR�������U�6�]�\nq��3�Y��1r��$��KQ�H�4�.bC
�^�r\@Z	�W�i��0Xc�x�C�߱  �MR�R���� � �16��@84�Z�
�ub����d>i��ZK��8uE�3n[�2�O1@޼������ �"8���k
ئ؋T*;�y�(XM����}�H:p��$�[�n�-����Fj��1�z��s��<g��f��Y[�m��* .y�x�b�v[���פo���{�s�{�E�X��E�ع �]�oW�ydӮ��6����æ-{?z�Xۼ]f��+��؃�tچa������M#ļc�M_����\Y+��X��(�)+�d�Z-��M7bl��2=MT�L;G��S��[��67u��3v�6���R�{r�wN��X�)]���=��x{���ye��z��\��T���lV@R�Ś�ļqs����m*�S5E��9��H�8�r�f`�tб�����^�R�f3�T*��@�
 ~[�֚W.[��9�Zzhi���.@��1�g��G���}�iEd�9�������k�z1�qo{`��ȭHr��Sl���m~�nY�S]�1XV��U����~�X�:� ���A�}1��U{9��V4�@)�FI��ԇ�)&����؋JE�p
�l��Wo(�r�\,�@��m���s��k(�[{
�|Kj1��:�D��"R�Z�q�lQ@�P-:�r2$�q���� /�ʙ��;�)FfA 0��@���:ݱc�nHV`�2�6���ɹ��mς"kl���ҿ߄��M?7��""��t� Wo�9��g���ޔ�n�e�i�c�n�>H5��ZC����G�葪��*6�T�R��_7�X^�1�Y��턷�"�I�ݴѻ~v7��>�J�����E��ڜc��&E�)�g�y���]n ����O[�0��W���X`,���6 ���L�&�6V���Ldgn_����h�<�ø&�;�����c˱]=�� k9{|��c� .v�Y�ּ�)YN�L�������o��?����_������n���x�C �~x)�XT�;Ib�R���"S�CN$��5|�km+��~��˪4�<R-���ɢx������ȁ��������k�;#����v�4�
zN�Ty�.J��E�w��n9wJ����.4±��ؽ�O���N��1�ls�ec�Aj��g��k��2���R.S���[#l�3�掶t�=|s綧I.JZ��f�!J*� ieЊ/`;1/�7�-�<�7F�pV䉞#��z�eG��Ѳ5O��9�qζ��M��Y��ĵ)-�JR�����Ν;��B0ZNiĶ������4]�S�\�������E�o�kղ/x�CD{J���M�F�C�:Pt��
h���h���u�,.v�3)�˘W�u � �%[����S V�%��\3q	�%ږK{Zz�x�{Xǝ����b}�������y<������M)
x�jtc�����d�Vy��|>vo�ᎵN���x�����Sң�Yԟ4�V~���4[��>��1�i�۹�\v؛�����׍�TsGE��ݘ�����>�y-�Nz���ǻ�V�ӛ�d."���ζ+�?y�'r%QXX���u�    IDAT`�V�E6WBpװI�P�Uc�C/ R��\c嘏eʕ v?̨���)@V@�2���Mx/���C�^�S@B20�a�+k�a��	��z�X�C.�����5��.���ZR���|>����2D/�k��.>�3�FqsNc23d��Z��n���i�;X뻈z�(��/`��mP9����X[����`�k���.ĳ�й��/�F3Vԧ�b�c��c}�u_^���<{@-�<`I����{��-���z`s�H�Y�qek6=�-ۮ�{γ�ao����s�K	^�Ly�k��׊�rz�o�P=��k��@n�|��dN!�֌�l֬�>���,����_�ﵤln��a��n�:�0��U��HG��ʱ�f���_��@Hoҩn~��O�d�j}h-�-���F�载�5�[�q��'zN3������Bg#|'Ҭ`���C�i�+ ���{�19���������_6Z{�>���X�)ƪ���Wkm� �vY�Q���|����1�+h�w�)Lq��Y���},kh��\`�����'A�3Cs���(�bmq'1���M�z,��C��X�m���&�re��>���ۺ+��\O�QBN�RT�|��v�ޡ1�3�R�^Ա
i-!ȱ�ɱ���Cl�8\�ͦ��5�V~1��f��V+�V�R�եZ�z�������͓S������O?��>R��&J?O;̇1��Z-b48-�J+��S*������RѰ>,5�����u�t:�n��Ν;�����t:�k�X��Ņ���G�O��u�4��`|qxW�U�u�t�� ���q�T4��9�o6��u(����'�1�r�,�rE�y�v���q8f�,KY,k.'��R�$����)��5C�:߁e��z��v����0 �����1��Ä7o��w�\�r���1��ju�y��(��S[��`Y��9ҁTN@�ʆX�LA��A��j�*��վ�X.L�7;�f,�Y�2\�VK������@]���� �i2����\^^���yXg��4dXz��3:F����WJ��I87�;���M�q�u��X�t[�]"�w�&��.*cU�1&׻G/5�͢��r�U�Y�Nٗ�e���r��-988�V���q����p8��{pp`\HNOO����0�öiV�L�1hP�L&2�v�̔0hf�`�c�O����.������"�@�KSt����fS�ݮt:�}���E�<�o޼�7o޸�����}��(��`	�������n���p(��@���H� �|>�^�'L�F�����2����j��p��Bf1�@�P4��RhM������z�mo��a���u�Z�d�Z^Җ�'v=�$�g�l6��l�����E�*��t:��@�t�F�bH&-F�aC�k=f̐�T��,��.��^Xo|�ERg�x�\�V���'GGG���/���R�TBp&�?k���R��<z�H���{��r~~��s��ՙ��m���]�[�d("���m
���걷��ήw�/�J}�4��$%�.��X��?�.��K1?P���.���������n���nK��E-8 '���AkG����"+o޼��/_�6��9O&i4��t��`���=�q{cKk�È�� �c�����ı�#���̀����+��{�m4!�� ���	_����1f5����;�n� �|��o4�9���3�~_�w1@F�Q���F5���)On�]�<���k�3��r \�w��w�x�	�f�Z���d�-Fѓ(����w <���6��S(|��0j�]`��5X��DELW�n�?�߰��%<?b�m� .��	0��ݮ�z�����"� %��<z�H��ӧ���#y��y蔉}%v�m�K���?�W������,��)�U��n%��沕�Lf.��>#�"���.qWcr��6�|��7V0�yƲa�ѐ{��ɷ�~+�~��ܽ{7 �f��V���_���E����-��������u�ݖ���p�d�^��8 4`Kz�m�Ã�O����Jd%�͔WH�q��,ry�;����Ǽ���˥�gsY,k.��P��F �8L1�̘q����@C���X@�e�L\��X��Y`�?��5��ytk�W�[�/3^�f�Ā�geY�t!dA�:h��'?ЀӺ&�����֏�[k�\� �A>_;Q����[����m6�An�n�����*�- Ƚ�=��ۓ��^j��,�Ky�ꕌ��^w%�d_E�N��ၢ,fю����]᫜n���>�{��j������?���Z�V��P$B� ��S6E�:zI��ƀI*����;<&;Vɜ�?҅M�X�lͤ����ߗ��c���/�o��[�n�,6R��`����L2Lp�j� �yF���p$�R9��85cW�}Ӈ�u�ĚBX��.��U�ZU���� �A:���)m=�<׈R�$�ZU�R]c�x���P�g �̠�.X\@Ȁ�V�I��
�2t�(�Қn�ƈ�o�:4����fOZ����3���Y��]y\p���r�K{���3��� �/�� E\�9��</� �ϲ�hH��\����d�ҭ}�5��UD�$����s�^�*��X��2�͂TEfZ#���(�z=��zR���/������L w+�!N��Ϊ�&=����%�z�Tqy���X�m��9U�����*����/��/���r2��E���"m�ի�-�z��k�H�Y�[�5�X�d��;��+0�
��E��|>EH�~_�ݮ��� :٥A�9��ӒZ�ˌW��`N����h4�ڀǽ50����]i�}x9��㈠��p���v���:YLk��y��1��iJ���Z����B2��>OH��|apfI��B� �������ަS���=�	��gsY�j�͋1V�C}��f����+�7�k�=0ОO-��QHl�~�f�9��� ���'�N'S�L�tەJEz������~��6�ʠ�
�����eV���>������Z�xN����#x���G�{�d>���ׯ�ٳgrvv4�bι��p�i��M#�TmRn7�8;Ƅ�:��1�~���)D�1	H�Km����[�Q�ZDN������gM��ߥ�:vM9����fJ>�b,o,����X��dJ��ZʫV��t:��`p-���nYiuw�t�E�C ��h�6�L����L.��l������ض5�'� +�1�����U����R>�]ۄ�*i��!�����\,���"R�R�.��>���W�X-�����: u����o���yz����+�3��A��qWA�yW��T��p-kL�z��uXE��R9̏����A>ā)�$K�N�*�q怗�=�b�N�:`ey�gs�ΦA�� �����:��wX��9��y 7Nr3�����,���UL�d�~�VE��������5��6���3��R���Ik�MX�И0�>�M�\�]�]7�����7��K�"i�w���R�1	@NJ"wY�/9����sq����\#��;w����t:�5v����Xzs�U稴�%*푒|��!��{�g�u��0q��v�3 ��\�E⾚k�Rc ,S� ?<�VQ�w����U��u��P*�L�� �*�*� �R�H������M�)������j%��\����Vg�ʥ�,�`��(�.*��,��B�T�Z�&�Z�ݛ<?g\��2<+Ojc����M��g/�5N���]�Rg��Yz}�@t�\�l>[c�Y�2��C�U��O�J���ڧ˥r�r:`�v8�n]�ǿcP�s��h4���˝;w��O?�f����cs��b�خ���P�c�?�B�]>�O�E��.�+Ŕf�W%�7�n�_ul�<s�ZzM��6#N-�j5988�۷o���t:��)�檻�Y�Pc���>u�z��&V�UHI�N\[eI"P���#�K��P���`�X�P^�Kʠ4��j����Q�:I��h��Y_ E��kĥ�ʘ]�E �RYʕ�5/����O��*��@�;���'ӫCݜ���]�~a9c��T�=C`�\HyY�X�����.]s]��������笖���n���YZoꁺ����*�}?���Y��b,�/�D#@@� ���v�""t��
~������kY<�����29���f]��F��[�L����j��ё����<{�lm�{�Tq�l��ƻ{������S_�Z�=EڏǺ���3w\���H3����}��ncZT�Qd`��I)ف��ԓ2g�(�����������P�����t�l�:�i�������/��]X��)�X��: R�J+�� �Չ�{�[,�N�eI tюfo9Pх1��P��	�g2�ć�.lY�UZJy���˲������wxyŝ#�=��{n�*�9��W�z�l�~��s��\f�+ۻj�*�j�Zkj�;a�\Y
���j��<K,-����j)��J�ŵt9��J��- ��q_w��V�K.4�@���;�Aڠ���ӥ��W�q`�k�\�� �zx-�:�i9���}�-��U*��w���bnz�(���]6B�Xԛ����&n�$!G���z�FdY������X�K�2�����i�ku#+�X`�5�T����|V�P��j���h���F��/���:|���2��g8���gҽ�Æ=_�JV��f9y�4`��`�x��kl�$=��&n�S�9����.�c���x�x�]�z�z�RPZ���/��:�Y�_K#h\���[� �B���Fc-�����f�aN�6V�l���`�W]JeQ	����_��:���6�]�	���vU���#/+��b�L���ԃ�;s˥C���dOK�0�8������lHL���J�i��c�%���*k�j���!6��Z�k�y�k��9%x_dٻt��!������(�8�l*���y}�D�V�;̬���M���"L�&���Nm[�JX��zO-�T!�&�&o��f ��we&�� ���͚0m�ϛ(�t�@k���.�6���
ܮVR��]G�����/��c���df1��Ј��z-k"��d�5<C����V��(���56*�
h)�ޗ�o����5G�0Gf���޺gFJ%y�v�a�7K���.b��~b&�,]�[�;+m��0����-�V˫�$*[�`bQ�m)+�ʕ�pu]�m�u���X I�7�Ǭ��E�X��xƊ���g),;>=�Z�� ^/Y�	�4��+�d&^3
k<xO�^�N�s��n+���'�J�EE��1�C
PyߑSg�@v��!gx�"������M@�凧+`���]��x`�Vw������4��ӵ%��0��D��C�ZUh��ө��݋Fa)��3�+��`Ώ�H��k�@8���%�V�k�=�E�r�
���c�^�ʌYO���U�?��
�ݰ�}0�Ё ���Z!��-��j�����d ܚ�lP����b���l*��/~���,�h���W��tQ�fZh���Y~�Z[k�-5S��:f�]��pЭ-�4C�s�'��p�U�&��e/hf
�YȪ�
� h��eh��%J��!EPX�$7��@��5�������<�9�Һ��t 0���X���
h���G.�ĳ�z�sߍ�qNr
�n�P*V$^�Ƥ~�1����;Eb�d�b�����ؤF�^��/�SO>O���e����?��L���FE���I9�l����9�"-6���ryy�ϣۓ��p��1;l�(��+0���rvv&���kݰ�iÖi���d*R��V�ؤ�^ �N�#�NGD$���h|4��暣 @�d2Y3�gv� ������� �_{~�����g��t+Y���N_p�t:�G;��b^kq�Z�v�X��B�/� �S�h�� �\�чV���@���l�= ���L,z-k[��r:�� �W7��B((�E���=���l�-����n�)�*Tc��,A�����Z�Dc��ZsR3��w0�1۲����*���yͮZš|��A�x8��JE�����V��砽�љm|�����>�S?����^����$ߧ|2�<O9b��jR��M�,������ ��V�cJ���CR�N��6~�Cw��H_��ߔ6iӮ"��h�{��E_n�
��`0N
� ��߼y#�^�
�`�)���T*2���L��\\\�`0X�&��}i�Zk���ah5	f8pk����&>C�NN����)R4�� ���Ѩ � Ђ���<���5Զn�4�mi�in�ۂ�����cY�al=Sn;���,6�<Gӫ}N�Y���x<��̭�Q��X��c^"�� �@p��Gw��{��e��u�l6e_�=a>,)W��> ���L.//���L^�~��JRZ�As����W�l@����hx~�F&�lc��=�c:i�-�R��Q��n�}�f3���-w{�^\[��Z0�+|�2�1)¦Fo�z�H�+Ҵa[�q���n�9W2�I��"��+Y�(6q�چz_�Di��),���QźqXũj,R�����/"v�M�*b�k�F�#�ܨ8� �f��D���F#y���<z�H�<y"/^��! @�3�����ޞt�]i6����+�駟d0��Q.���,�t:]cy1��o����k w4�l>�v��i{U7#p���Fc�Φ3��g������!�
�upp��5�eݠ����}Pt:���Z?̹;��-I3і��j4�R�2q�+�1�g��|>����bo`�6뀙0�;_.������_?ϩXfmگ�p�M4����d:�����C�W��򑷍]�����������ܕ�"Aㇹ���`�1Nxf���%�\ݩ���X��ӾT_�.��DRʎ.��Z�0��|8 ��v�rxx(�|�|��'���%���{g����6r�"$��=�e:?�B���(�G۲鹘*�����(j��Db)˖�zX^q��s�3)z<�n85�<I��5o	� T-��7Tw �R^��l6���sy��������#����	X[0���n����B~��� ���/�ˁ��k�ÍA�ǔ�ɛL&A��	k�}��uKV Mfޚͦ���5m&��jU^�|$HA�1�����R������c1��`I������S����y�re>K(���y��rh;:�r�S�V�&K3��<��h�Lx\9K�  ��^f�4x�1��Y6+��-�8�P�V�5Y�ד~��s�l�h,������y��I(V��5 $|�Լ�m�e��9hb ��ЖW�w�X5"�|�#H�\���3�.֟����T�ѐ��C�Fa?`�Ɵlr�U��&A_�4��4˶~H�m:���}����r���2��|�5�W��`�g�cEg�k2�6��Dr�i�>r#|�����J��yUj�Pd�r�9XN)�����\^^ʫW��ŋk&�jU.//�!������k:_\��ׯͬ ?����k�N?.��v�k��I��p�{���1�p�����Jգ)3�3�/40�4 �`h��=�%x�5,�Lq^ ��r�V��:����Ve�����T �}Y�G$�\-c}=��;T3�f���4�c��b���` /^����}988�F�������G��p8����5W�odX��XQ7l�1�e
S��T1��R��j�ۏs��1nY�ž���k>���ٙ,�˰��Z����rX���jY��A��>�ƾ;��`W ����J<?H��ҴZЛ$���X���$�P喱�&���:U������e�Z�n�4\\|f�'p�wfV[�֚5W�rz��1��s��!���5�A�+gs�E!�l���w���>]E��*���b��z�~��b--NN,���t�ll�cע���g�#�&�k\ی�=��0��kBo_��A'3�V1k�!5x�����}��z!C�se�3��>��m�    IDATj��N�Lsȑ@)���4�쏞��^�{V���R]B9��{\�Q:??��ϟK�ە��c�{���=����N#J����mLg��E��C�'�"�{h��B�u�xMR��1�x�J����(%_�9A�d�[i�MS9׽+�6W��	��,�\�ނ�� ��ֶ�lJ��,��VI=��c��11׾��*�QX��q�������=Ӟ�� ��Z�L�v ���V!��ٱ�
p�E�������H�vKr���L~��^�־�b������3S��+���=[�	f�dR&��\\\�˗/�͛7kŔ���ʂ�$W-eW�.�-)����J޾�pc)����<'k籚�\&���u��'�U�A��#��L&r~~
*��9d�]�\���=�P�"�v;~H���瘛���X��[k��=w��9U��Bo2��C�5_)�67P4
H�X�]	�=�y�O������X@�so(�ѭȦ�bSQ��Bo�c��W��.�+�GV[�0K��4���A�1�)���)g�b/}
�������4}hŬat�'ff�5ۣ%
�8�-�<�6�V��1P��˭��e׀�K]���z��=K8H�a�k�/���^u�_��ch�A�����R���T+�����拹,���˰���b=�5/����}���,�����{Px��%�eRY���|jO���sӅ��6�����z���n����"x�`���J�m׻�.S�1=i�)E\�\�vU<��u�c�6��I{r�m*@��L,3c2������ �`�:^Z�c r�L�a!S"�M��ӛ#��I}�*Kcj�@*=K)ŬlP=�*��3ֲ2`���2��5)�� �_���`�Tt�5ږՎ��լ^��kӬ�Uk�"2 �@�%�� 1��9���7�ޓ�eSK;�A�n7ju�b�P{u����zi ���ϴ�~��3j�W=nU��!f��9�+c�r�l.�����L#��n�+�N{M2�se��_5�x���f�`����w�JIyY	--A��� d�7�aJY>z{��*9Vϑۆ9�=�&\x�;s���|>�z�.������/�V��Z��WE2�)�e�r�"�$���� �9�`ٍՔ�˼��\�B�빵M&��Px�4zn{�]�lb,jJ,n9.��\n,���S�*v�B�zkBy�3�-���|�kV�7V+�+ڰ�I�ȵ_�w�X����������c���N�zmn�t�G�f��Z��3���'UQ&z�yY-��?V��f�q��3�wf��ɲXPK�aIV�h��7ͺY W�س�/�\,ײ��c�����r�,��/�0�4��1f?am	� <�la�K;m�Cn���x9lL��<���S�o��_���"%�.gx^r �~���e;@��� &��@I�k�,�����h7��ZnQ�\�����	\�K����I=k=��1��c��������*z��9?/�YkM���&���m�1���96.XB�[���,krs�A1�\�m����mQ��`}v�2�+���b�*��L�i�mk�ydvH�oy�d�,B��c��Yf�c~ۜe��4��:[nG�X,d1_�l>3[&[��8̟�Y7��J�a1B"�+o��Z/W��!�����aL�)�[w8�4m��������o�i9�2k͖��p�V&�A�l6Ŭ�+����~�֖Җ�V+)��k��V�%1�Ե��%)�}O��ҍ-؝F�?s�����5\���Ă���.��.�m��"�V���.�}�l^�����f`����#�獙�ocC�&ۛF,��3x�x�z?����)f��_ZCj�3��+Vx��p�W��a���������g[f$��d	�����K�����-i��O�9z�Y�B5���!ƶ�=���J?i4`�i\�7(T��w�T��m���ph���Zz,Fl]Z����R����� &p��}fc��Ej_b-�����w�c�976a�d2	k����>ֳx�:Nj�=��S{�'���%)���0hGs���ypc,��i,����n,1i 8�n�l��� !���Ы�;;��͛7���e�ZI��]�둡`6Wg�>&��M@�M�����DlONe�wERz�T���wWS��J+ĺ�hK�S��P�M-��l;�=�
=(Va�彪Z�����̵3���Y�iG=V�k6���tG!m�k��b&0pP�>
���1���fN�1�a=��l���ۈb�*g�/���h�9��֧�[�a�`-3��{N�6�1s���)4��D!Woך]�k̚�t�*�5�fi׭f6:�Ҍ1�0ˌ��>k42OB�\�<����8����5��&���_o��2�fNw������N����+���D=���S��^� �(ļ��c�y����㏲X,�O>	�*KQ4�`95|� vl�.�E�A}m�}�}��E�Xv��x��tL�hUX��	k����S�Qv��R�����.px��E4JEl5b�lj�-Q:g0�� uZ�S�Z��U�I���� �S�"�Ϡ�2h1��ݰ��2�=K-���-Ƭ��>#Vl���.WvON�@p�Xjz��2ł@v�n����I��v5��Y���𴫇�G0���Tk|�����% ���Ar�l6�@F�ΜX>�1}=�hQ����s�&��Җl��7�m�e�b{B�����0�ߋ��Vݳ���7X�v�-�rY^�~-��TF���J%��롫���-�·�ڦ��;�Y{c.���zE��-�o�f-�A���%QȽx�[ڪ��9�:6=-�D,"����غ7��7|�$�R��1�<_w(�E�gp���J{�t��gX�V���v4`�S����u(�yY��.��U��9��\��Ydi ��bd-g�*/���AJ&`����f.w�����]s�V��xz`7eOe�L�Q���vuVE�W�S�����N ��&&�ZM��LC�`�9M���9��x쓖�����T��(��y��k{8t��ج�㽒3Zh��4h�!Q��frxx(�����t���d�+��w��-;s���@[�>���\��6�5��[��صU7y�9�VQ�gz��ؤ����7�vHo�z��V�ٔv�m���&���4��g���	�"��d�t]}K� ��Z��V�����H�ݻ'����n���j<6���lǴ~8��s�u�`0��͉��lh ĩ6�'��CL���IC�,�<�k�Z�v�ŧ�90��c�
b���(���T����?x�'�񼴭`Y��2a��7���:j˓�*V��R�;K�Xs��h��]a1����ǲ{�� \H 3���e���Jl�O������|B�ݠՑ��7S6c|~hٌޛ����I��X�L^�����B�>}*�oߖN�s�bm:�^s�5�*���@r�}��k[r/�s�i�OAJ���@�٧�,e=%����沢9�@�B׋<�>�5�N�>(=�)��A(_�ץ��mL�at�%
�!yV<� �����K9;;�����5�".���nI�M���XW�T;�r�,�VK�����{�����AG�����-�L�0�@!��f3Y҅�h$��$�'��t:���0���I4k�������	�J{{�?�r[�B6�=���k�E:@yE��K�n΂0p�ϓ��U��^w6^�xi�=o���?���0�zl�@�jml��g m��r�Q0�Zw�Y�TFL�#p�54�,Wl��ϱW�`�Xiym�=V������^�g�][��vc㽐�A�ൃy�6s��DNNN�ٳgr��m��z��1/ maB�"3>$�ꝇ�� ǀd�����w����6ߔ�H�����/q}p���H�2�a���fc�9��B�V�%w�ܑ���˝;w������B�������|�R=z$?����������^����!��-��h4;�pZ�V�T�v�-GGGrt�H��{R��Ms}��t���Oχ/�R�ͦYt����mL�k��j�K_Z��E��u?E�~)͠C>L�><iV��^Q�����Z&��C3�����f �6 .��%)���Fl�����(k�y� \����Œ^�.f'�C���ٷ�x��:��Η�l�&�/Yo��Ϛub�`��� e�Z�XgƐ	�6����l2�Z:g1�:�-"��&ž��I�m�ᱫ��a�{ߥg�W�`fr�F��kN��Da��"�:�2bS�ǁ��ꫯ䷿����������J�����n6����̨.���bk�á<~�X����Qo��A^�x��Z� rut��Y��U"ֺV\��ɭ[���y��"%x��.�Z��\y�j���鄢��	��s�HY��9�L*�c1����+<L�x�W�{����b=+m_�VC�z���mH/�_�����8[�9�T��\,�s׌����FtY��ʑ��z B��e(x?a6za.�BQ|r���;��c���[s�wٖ�j9�3j1�
���˸���-Oi婳���l�8[ ��[���g3�9KO��Q�ץ�녎fz�Y��c��n�>&_ߜ��E4Ĺ82u=�,sjl�79��9]8<��w�Z(�}�r90���Rz��ܿ_~������A~��_����5��jcl�l��5������K�ӑN�#�~_�_��_���2d�ZI��\۬�1fݴ͘�V�Z���jk`���p Ӄ�����~?T�jͬ��r)����.�����^u}�c���.ZŜ�;�N���e�����g�UfY��HT�U�UkW~���H���$PJ��n��~4��_��cM�@>��b�[�T*_�5�緝��������i�\��jyM[��^��\��X�G='�߭t%�o[�VRQ)������<����0��Ƶ�@�2j�^[;劔+�k��V��f��{��P�I�zq���Rs�(u��T����?���f���Un���9>>���#�s�ܺuK:�N��<��-�}l�(��9ů���#�j�������п��$ƆY�������l6���@>������7���|���r��=���k`	l�������f�W̠a3�v��_�Jz�^ ��JE>|(�����Q]��.�[f��������rtt�BF|ߩ���W�VA@�ە^�'�N;�VU=_���е��i$	4Z�c�����Ns�ߥJl�F��ӷ���\	ݘV˷-\I*�����\.pşm5ȵJ+bţS���D��\\\��]���3��EaVPf���qb��?����R����l�_�}�@� ��{��%:`�a-���L&2�LH�v�k{)7� ��K7 Ny��{-��N�rqq��6���Y�qN�ݹ/W�cI-�0�*b:^v0tX��j��Xd� \ٖ��n�x<��|.�N'���n���O?�O?��J~vt$�n7�N��fʵS��r�-�bVc7%/�ԙ�#�\��Ω�~�F�!�$Xt�z]�ݻ'��ߗ���Z~�����~%h4��<�t�\��X��f���Y�ݻ~��nK�ӑ?��ryy@.�I{ޤ��{�8�...�ٳg����t:R*���L�XY��v�-���rxxX[T�C�����<�lp
�bJ�!�=1&_l�|�-��f����5`�Yh����2f��9u��υ*��h���c�&�� ��Z�fJ�,gf�"���4:��Zq��֩^����������{c�$x��24�`w4x����EK�tњn�\�Td>����TPmItr��Y��XE�O�1
�:��1����0���Nko�c _t�c�j�dooOnݺu�r���pf�?66��2���3O��1��Uo�N��.��yV�~�g�c�w���V�r������?���{����O>	U���Fk4�/K���HD_�b�vV�VK�޽+�JE�ݮ�j5������N.//�c���6��6,1����bÃ�L�ד~�/�~_����V�����8������H�Z��p8��h$��@��a��y�X~�)R���bN��*�����4+�}TW���/o��-��9��i�ĕ�ڕ@�>��yfvJϟ�P1��^�(d�
�"�]n1����Wk7c��G?OO����օ��x氄E*�5�iI`,�@�3�"� ��C9���K2�n���[\�� 4�+;�}G�z 7�e�r����1��vbA���X����f���y{�z���"�[>��u�
$Z]7��|��H�M�k�T�A�����-��+�;��d�D�Ul�l1Z����l%6�� �^�T���=��o~#��?�'���o���8T����D�Y@��1��]�8(�F�p<����A�E!%��?�Y�A ����k�{y�15� �'���x�B���������pH��f3i4����R���ӫ�/��^:��h��9���8�\������rZ[k4ֈ��E����*��3�qd]%�\�L9��K/�nj9(X�k-uJ���h�S��.s�$F���"�<�W{��zӚ}�=�n��g=�L�m���bN��5��J��-n��R+�3)�:�2KV�I�a��"*r3=�B�ss��\N��i]���zB��{"�y��e�v�AW��Í����MD@���q��/h(�k�k4�1��^��	M5��{�M#��>`�EUD�s O~�C������3c��wW�ә-�t:Wv`_ޗ/��R>��3�t:k:4�N�����3o����L�>�XT*�����7��j2��_�����������4�y�
��L��k�~�,5��ԝNGe?��ZM��y(D�N�2������+Z��ƗYN��4z1��
-V4�h-�i�jQ�r��j�ת��; NX?�����[[��3����pe��ޘ�Ļf��@��-���" �+��\+â�+�����xm~@����~~z�!��xV�d/�[b�M,#��J�Vk�;9������[�Ȭ����33�XS r*�J`n;��Z�?��d0H�Z�N�#��@��t�ݰ.����ּ���u��#9٭�tu�L����ͅ��1��!��h[n���RK�ޥ�nW�޽+_��|��粷��=�^�pLV���պ�bJ�Y��`��3.̀L᫯�
L�j�����@s���_d���V��:|�w�*A�P�T��h��D�)��|���Yϛk�<�ڬѳڙz����m����Y��xk:v�ֽ2`Ӫ��r�.�Dј>pY佴&�b��nU�����'n�����m���:���C�#�}��뭁eh���r��H��K�^�XB�a�⢻���_�}vΡk$S4���/ϑe�*/����^�u��C�?��T�áL&�5��o��ں^��a�X�ۏ�e�}����dV��`q
([߳m�cNi����~�+�}���w��6 l���l��7 \��`3d�Q�r�;w��F6�M��?�!�^�
�g`Yr�&���&�h�V���87�ږ�e�7ꦇ$�Mgӵ"�"]����y]L�.<��g�c S,���b,�'������\tǬ)?�'���ek0f�,�|���^&���VG�Ԝ�ls@���[��u���v;� �0�(:���d2	���h2���,��""��P���57�(����CL�le$R,��,s,S��=N9@X�ޚ�:�g�1�ܔ�I��9 ��=�UN���;eS��!���iw�]\ ���m�����b���"�Xꖻ������~���?�A>���ᶄ�v	l��֛�R ��AE*l�t:]�<�)�Z�&GGG����~M�8�O.��mpS�T�? w-��j����l ��b�X��F�_��|z���S���Ӽ!�c����ޫ�Ij�xl�%!�>�Vw).N�h�G�u�,f-��s��"���as5���'WS�[���=��j�;P�Ǚ��d"���k�3��
 ��~_�\._�������۬��S�������^���f�k���R$b��lq*#���Z���\���m�u{s�s��C�A��bYcҟM�������k�WՋ=�'�\ α�}��    IDAT:0�6<��ZF�~_~��������o+_��t�ݐ~�F+
��)5nm����3[�a3o4��t��l��V-��Q�ѐ۷o�f����������MX�Ԣfc+���Uat[�0�l4��*emr�\Yc8��N�2O�xx�66��9��}��O��5��X�T�h]��+�{�逭�����ɵ�`�CEl���6�O1|9��c�,���X>���4��]OÞb?u+���.e`�����R�ƵB/_dWf����%iT��p��(��E
�r��s+u�"w�}�j���cck��+O^�)h��S`"㇟sedT r9X�y� 7�a��]˼}�)��E�ଢ଼j�p����fP��|n4�Ґz��҈���}��������������_ȭ[���M|��=??��x,���ryy)��8l�E�u�\�a��۷��/���w�J��\��t�6�G׳���:t��t:��w߅ԟ���DS��(t�+<��d,��0��al�l�����,�R]��V+Y�2�Nd2��� ��-K�9HM��y����|L�ʹ�:l[U�ځ���+�I�g�Eݴi�%�~�b	�Nx���~ޱ�-�ߢ���f�� <V�ȿ�!8���P�Ͽ���j����R��ɺ�z�̍^�1�i1�`�4���&g|,�~�@1ե3%i�Y
�	sgPL���X;���S�9�� F���)L�:7s�e
�}�`6g��eq��MX�-Z�P�w}n5fK�ժܺuK������ܻwO����^��b-�us���p?~,�}���|�R�?.��p��J�P�1��R�ȭ[��׿�uжݺuK��������i�Z�&�oߖ�j�|�2 wn��.�n�	o��` ������� .�`ĸ�l6Zr��0_�b%�Yy�Ο����(�^
�j̟��6�PȷZ��i\|e�	~�ju���.Zcm�;K�k���n6=�-��K�u�7'7]�����Z�Fr��x��.�K�����x��rQ��e:����U�V]�Ѕl�Y�S�.RZPo��ȖM	 �$J�T��;��7�8x��t���N8(b"!�@������M �"�6���f��[�V�~6a����Z$�Iy�z�Qt�Bnj.U�� kooO�ܹ#_~��|��'���E��Z
�/�nց�����LNOO�o����������s999��xt��;�Cej�\�[�n��ׯ�5N�^���i4kh�f3 X�հ!�j5�{��t:�N����SY.����c��ص�ָ�������^����-t�C!��*���/�����d1���5��=��[lSl~k��%1�W3�1'˳�:8���= @$k,���J�4qqY�H�jTa�Ml95�c�.�ANO\��h�e�|� ��c���x�6/a����ׅ�2`����7�=�,Ҽ�M����r������
�<6�ߓ��sF�,a���g���;��v��&U�RvB"�Y��޵kV2EhlCx����H_��H�{�g�k��"ٍ7��JM����9�6�܂�X�4
��ۓ~�����P��{BJ�͛7���������[���?��ׯe8���=��-k���C�����իW!��W_���t�Y,2�޿\�lq�ic��R� ��۷��>�'O����I8hveМ*��:�~�/rpp ����j��=�[�mrJ�ӆn됳��q�++x�լǪ܋,�IϵXF�c�,&�rJ�f���Ơ�e`� ؍ףS�lA����E��6}��R��=Z��u�:P�u%���ϓ�^�;�Ŋ�����q6�?u�>d
�v�&w��e8���E(h��_�q�� �k[j��goy�{���ŏ�Ϝ ���Ę_n���j���D=�a���x�|>���K��������V��r:�5sFq�};w~�=s[���W���M�C�ck���H����g�T���Hb8f�K����)�e� "���y�������w��Ç���$ g��,0��8b����3���g988���۷C���` ��^Ɂ������^ �E��v1Ā�Æ	�� Vޙ�� $�}�<!Uɞb�b2���]��aN���%+�� ���"�c�r�%��d�	w���q��I<�O�����9P��cj#�E���z���0�}�`r�39��Z:�B@��?�b�'7h, ��[I�����X�㵾�Bb�M�T�u.X,�5<�PN��i��r����Z��l����~Ȯ�#צ1Ŭ�p��W�=��+��9�c���n{C�ۤ�z�zE "W��GGG���/�v�Ly����`0��O�����7�ӟ�$��_�ٳg�5�5�ͨY�L� ���B��_�En߾t��+t:��bQ3���z�g�R9.
 ��z=�[E�`E�\<�EF�J�~,1v#eӢ�Yf><�'�����Z�L��M�[�q��X�|,]��&[�dW�ra��\D�-�c.��2�?�]M5���J5���n6uh�{�^,�r,繇���[���d˅HI�5���kJN�{rXŞ*��6Af�6����X{�ʽ=�biy�Y���(m4kDM��+9�e�cSf�(��p�0MQ/��ɵ���S�����T�`/�:&��!y�tk��)��ߜ��/��B�޽{����<��L�S9;;�~�A����Y���?�ӧOe�ZI��u����@>�P�1�d4�����w���w���I�ە�r촘A��V�%�FC�����m�X��5��gO_�ix ��
�<�L���bǼ�S�n�ܲ����ܱHy��*�c��x�d|x�h#�bIR�C�����%�E�a�,v�c,@��Eh�[�!��UH�y9[�E��֟���l6�\K{�2� �~���=ˮ-&�ɑ6��YT�w�u]�c.	����wSPe���3���F��Uk�4�x_�^��N)`��M��X��_�5�&��M3�^�F��x�����C����/E�g����l6��ݻ��g�ɝ;w��ҽ�r[�Vryy)�=������?�I?~,��4J1#�{Ś"@v���9??�j��o���JǺ �Z-g�F#�ǁI�� ��@�Mn �'&r�>� S�9����W���C.vŘ;�! �A�&}�Z/bg���N�`k=j �[@�zc�x1��>Y��-V�
����'����^��k)/���?�qfp�`��2�: j ���!cO�|����N1�Z�m�g<��
4���5ř�3����c�����c���=�z����� �v�-�V+E�ׯV�0����q6f fS�ˬ�j�|m#?���&~湯�67��W�M�0����X��`	�w����t:�k��g/y���<|�P���;���e<W�m�M{j}W8��ey����\k^��?�!i�h�&`_v��Ʌ�Y'�&l9Ûh.���n����Ɯ<��;�r@L�b�`�
lS,ϵ`���+d��䰰��mv�������̬���
��x�2S�V0bI4,F/�z8�]z������Tʕ�?o�^܉N�Af=F>x���c��+����[������
�,@�S�j[�?l;H�J���岬d]+�ψ%F��c�����{�^tg���;8�E ���hk��[�;�^z�&���N: e�rxx(�~�8+�͜N����ky��Y𺅩9*�=w��)U1���ޞT�U9==���s)�����eoo/t=�V��ViA8=����˗/���<�W�Z@��Y]Kb��Q�P�A��2�jV�A@Nw���rcF�x~��5�}�c��I��]�6u��:��%n�sB�}�+��>���T�pLu���!樢C�H�s1g̭���
�bL�f׭�*�JY*�J`#Y��m�9`�a ��4����c�b��X2G��+VM���eF��X,d2����V�I��g �'��, ���L�dqc	��c�ԏ��΢{s�}^6q@�z�(U|fm����c�c���f3���lf�ٌF��H�á�|�RNOO���b�]�LX�K��iY��=X��h$?��������Z���ٙܺuKZ���Z-��z2�L�͛7����/�?� ?������_+d���E:��n"�8�&����IZ,�Z^i���n�t�6���
��"U�|)�"�X�9���Y�, ;Xv@���@�0^�L=��T�=׬�z�%[�i�1}۫�ҭ
po���K_��/zΧ,0h�<�9�gi49`�=K[ Z�V��xsVH�	�K�e@+^^��q�W|����/�b-��^��:O�wc�'��������\���l���Z�����Fq����2^����>�mn!�p���՜��J��bjS�a�Y{N'��i1t�999���S���d��g�����srqq:i�a��)�j�V�^�$���999�?�����_�'�|"��ߗ��#�N����?�_��Wy��<x�@~����z㐣��d�S\�18�!5�Ne����Y�Lg�5YI|��/Ҿ�9�Fk���i=ͮn��c�I���$VШ�<���ƣ?+e����{j�xvc9mcl8�K�A��+-:9��<��+��1D�k˛�^�^K`�s�:`��{6�I�^�<0�Ao
������岄E�)�7�[W�`)�˵�E�-������c_F}�wn�뷂c�{m��,�s�pDL�Ik������a �;�wU+���5�M(��(��=��խ����H ʼ����53Ɔ_�ץR��x<��` ?����������w�����Çr||,""Ϟ=������r~~s��e'w|r~�"d��`%4�N�,�����j�z�e�R����L�x:T���'��֋�tS��0�M)��1_���XF�b<��$v �Z��x��-)��_�v����+��9�}5v��0P�i�5��H�� A�{9g�4+s����0W{n�5���h^Pg����L�!����2U؝r$�������|�V���6J�[�87�V��ґ�c/8{� <%'���xk�Ad,J� �>4�����k'���M���������ַ���"�p�)R�?�|A�pzz*Ϟ=���y�������b��W�^ɳg�䧟~�r��_ >K�i���2EZ�Z)h/��#r1����fsXau�ap�b⽮4���z��X��Ai�i����^֛�޼t���xA�稐F�NZ?�X�[+��9�RQ*ۑ�A�^<Fղ8� �"���[�Y���v���J�k����%{}s� g�v���g�����*p����լ��HL#���T��3�[��<��e�`���d"��08��f3i�ZR*��n.�-�	�Y��w�����S����An����Ǜ�mu7��u��X�s��f�){{{��tBq�d2	-u���4�E��sЛ@X��l&ϟ?��hR� ��Ng-�+U=��턊uJU>[�#Қr~~.""�F#4���2-OC{P�G��)�c��9i��,���9^�:�`�i�2�c�=f�z���M/ޏ��y�@�mNzq��Jk�s��XGD����hW/0��
�Z
���ZI��Ú��4���c���P h-�Ѱ�8e�l�{�G��"���:��E��^�ro�I��Tց�1����s�L&�v�ݵ��&�8+����&gR��@P���}��qN��;�z���8��u
�$Z�Ү\��Q(�\Of�´�b!{{{��_����e:���驌F#Y.�W������Rk�b��K��;R�(@�k��^��=֢2��-����7��M�F���9;;�R�$�����v�Y�j��՛�>H�0�&�Ҝz޸��)�b(g���P�p�ō��)��W0�*�T���Y�9��,clL�J=U�n=�Tq��I��k K5��Z��ż@-�@k�����}�������j%�F�T
��܂��L���S��^k1m���-y��-�k�kP_�f����r�P�MB�e��3p��;��0/c���3�����k0P�ɯZ�\n5�>�R�n]��L��,�r�&�O�H}��֚���j�*w��Y����2�u
 g� �����M�[���`��0R��8��Ɩ�#�2��؆��K [��,�`��G� ��_�0K�#�fbc�n�w< ��êJ�E�Oz�,��n��
Z�B?�,����T���Mޞ����h�I%��l����d�1Kvßa[���^7#�V��ؿ��rC�c�}6w���v�����5��:cd��)�eS{Z,���*x�i�@k�X�Ӏ�=t2CC]�<rω]1�^ ����gsS�9�n̜��}Xls�n9��e���.wj� $V�^^�H�7�����y�䉜�����8=��*-Ms��p��t������Iz&��JuJ��ئp�����d�<����R��9Ѻ״��ǘ3��M1����,����5X�4+kiv��fU5x��/�6�P�w�X��Y��<X�ZZ��ə 洏����R?S��ÿ{ ךז~��-�8���sD{�j��)�g�[N��ԁ�C[��e,��7�b�-��{gN윍uD����r���H���=>c,�o/C����s U�l/���W�{I��t�t|�� fV�]�-����ə6�(�^��M�=_�M���R&�������$t/̫巿�m ��H<x�ց �7�X������$<	g�ٵ��1Ωl��qc�Ҧ����
��sEǶ�b!�r%��OE��X���C��S�����u��S=＃�]����F,S�����\;�[j5w�y�!kL4��X�X��T���{�e�t�"��[���%������ܡ^��J|�{l��b�;~<�4���
-	�H��6�&!���p��O��z�v��p�v���%�R��������������c{s�����VX1L��.��9�T����~����ܔ���.
��Iy��m�O��}��u�
���P��i�;w�����|�R�����ϡ��0ObN���Az)v���U���˟kB�ǁ�+ȍ�r��(�^P��9�ІgY��{[�ծ�����a{�1�`(9 ��g�:cr!OG�k��/�a���n4A2&�5���5|@�ױ>м�c�<��5s�"=^s��S4��t��u�창T���M#tg+{�@�n����%�5��^��Ys8���9�X�3�u�U�9�b`$eY�]�6�ZV�[������Lj��wo�a?���"זk�h�"�S��~�kI����EE�mS��&M�1�9,I��=��(��s4���ē
���b!������sy��� C`׃�/�j�*�^O~��_�x<�Z�&��X޼yA�,B�#�F��ѐ��K���m���l6��d�����.�W5c�{�+��X���������`,^�g����硗�NF��s�r��9�K���%4�`G���?U��1!Vz�
&R���h�G볽���1El�b���N�{�h�$[g��=��9��a��C�y�̱��^ki�Uׇg�ְ��b�αg���Ps��AD\�	M�����Gw��1���v� ��%��y�r��c�5M��9�� ��n*�C4}�m�7iUDf��uz���0���Ӛ֚����1XO��?99�W�^�p8����� �(|�&��O?�F�!�RI�������ɉ�����9XGf7��s���?�N�
x�6���S)FsSM�U���:��L��D����E{�ٱ9n�1�A
�)��X�\9Dj}�4�1ד�L&�k��@�k��yޤ�0�a���s!oK�|�~�*���ˊ^��U^w�e�~�X���c�����p�-���2� �����1��X�An�"ݳR�E��5g�fjv��1i�&�y�g#4��+&��H����g�f3�N��9p��HmB4y�ڻ���^�4j��~,�u�nsS9)�.F9�����t*gggrrr"'''��W_�����Z-�FAӪ�j��4���nW�FXTO�<�������e7l�RIZ�
��    IDAT����m���b����S���������͛���
�r�4lnc޶ށ`U�C*½ޭM����\�󹬖���9����\Z�b�t��.N�G��Rj-��X�!�J����x<Y���jnڋ��v[��H���ҎI�m�\�z{h�{c���c�
xmU�kց	?�V�W/�R�l�I�b��	�&��!Ud��Z �H�{����D&]�ƚ3��ZMʥ��䗬(�m��$|,�ӎȰ2�²<}��>�9��xy�n��\��h����jw<V�}��9R���{�F ��F���܋�c�n��tM���y���B~��G��ߗO?�T���K�V��r)�� ؃a�q�P[����>�N�#Ϟ=�������eH�s�Rvt(�����eooo-�`�Xȓ'O���X�>}*�=��ϟ�x<�\��A�8l;yc��Fo�xiclp�h7���rqq���ji�~,)�&N ^uw����Ɠc˗b�r�NN	2�`���S)����f�B��ZT�I�#/�U�ЉI�r�y^Ò"�l�b�c�טg_�B���b,d�ى5�R���[�����Tu�~OL�c�s$��a�q;�Ld8ʨ;
�~v !���V�R�V�\���a�A�� ��F#Ԡ� #XQon2��V�|��f.�j�\��q��f3�����ppF�*2�0��c�?����<��n�A1{����$9lG͑�dHm�F#y��T*9>>�J�"�|�ܺuK�ݮT*���Xld."kZ�F�!����j��֭[��e�x�Z�`0��h$��^�'�^/,FN�.�w�|��'���c���o�[`��ƌ�e�S��bu�﵍�����l�,���FR�T�Z��m��_�`,`c�r��tbX�������0���H{�rђ%ؤ�<փ�GO�*Љ�P�i�c}M�0+�{��,����tΜ>e�V����p��m<�0�%l�mn��6'c[��-4�̏��\���@XYd8���L��5b�Xʪ��Z�� �\.K�ݖ�w�����4�Mi4�?��dI��vg�7��Z�@�C�(Y�=��x��1�0�Go��"dYIP � �ꫲ�3� \;w��ܛ	��c)����{�9g��^�@QQEƽAF�� .
*t��6V�M����P��>x/������ﾣ��3�S�W`��Iּ/pb���p[�9ZL&�(���6�j�}t���捁��jE�^��?N���A�^�F���׿����j9�z��e����jE�|����x��^�G��`�11����|�Ѡ��C��>��m�����4�f3����l�߫̚�o���t6�m:�鉢�*���K���D��M�������52��T�8�i���<�}�ۼ]S�| �
o���������;�nS���6�Ӣ�m!��&�ے�='�I�%?���6d'g��9�Υ�����=���ί$�.w��C��n�Mַm�g#�h��L��L�S��@],��-���"�h���k�N��X,���>}���tpp@�r������ጐ ��$8����F�U���Ml]�>��,M&z���9����c�\Rg��|�������M�>�ޖ��ál��2�̌�%	alCX�yg�Y*�JF����SD�&k���"u�J������̂�"zYq� 	��hݖJ%�|��?�0J�5�McSE�j5�t:��W_��	}�k��e)\��6U���m�kZ-W�Z_�)�f��C\kAK���=�>V5Ċ��kk凶�l�{��͏R^<gR;�� ��Y�綠m����u�l؆�|̰���B0�*K{�B"�5p�=7R*�Iz\�UD��~C:"q�I�����Z.f_�[l�6	�?�Jg*]�{h6��r�L�R�����:�+M���(�����>��C��/I���&1?��&"C�h�Z.? y���8Ж�E�T���I� ���j���z=z��5��s�}<U5����[����%}m�� 7Ԅ��ڢumdq�C��4� �L&C�ٌ��>]]]�z��j�J�f�J�EQd���!�Bj`����3�xx�[�!���] �o�ZƦ�^�S>���bA���fC�q�ܓTo.&������L6_��g��s�T(6����,�3kkj��	qƘ���|�C|]��-5I��v���oC�1��:�bD2�6 �z��ZH�k��&YW۳��a��t��!���U) ��� ���G�b�m��d�m0��l]g�mhNN·��$$�-�/�k<�m�y��&�>v>��Q�R1��|r�._B�;
� ��j5�w�}��tttD�Ng�a������A`��YI.��K!�0��(��������.��5p�{�CՉ��2	��uV.��D���>�M�������O����!
�裏�R����T*e$Іro;��� @Z�p�[�w���d2�h4L��fi�X�p8���+�N��kј��!��nr�r+hh�o�O�%�h>����8]�-��AĶJ�_p�!�-��>{�P��Dg�3ɀ�4`$�u�u��x&43}۵q�C-�WþYWJ�����hϑf��+lB�"Z�j����`����� uuBB]�ݑ�(	uF�{�-��Fl3�ba�ۿ\�4�j��8�a�F�A{{{���O�v�D C�ϻ�8C'�e��p�}^_GP���r�]��F_���C30M��������w�?٤����Lȁd�T�@s�	�g�����?���d�Ï>4%Od��ג��<2����EB�
�T*������h4�����s:??7~������J}�r�qA���ۼ@�i���������b��ā�7[�6h��[���d4$���9> ����{��	_;6 ��+DllYW��˂^+�}��2a�m`ҧ����!��q���Z��:.��ob�s�b�m�/��}��q����������\A��u:::���j6��و���j����BR��+$mE��_X�;�f���^��|@��r�=}������^?}��xkWK,.;�yᆀ_"H|��a/^�0�`�l�(E�����"���,��� ��>6;%�����d21"�JQ�Ѡ�=����d�h�0x1-�w���!	���>���f���R)J��j����P��+������@��È���tE=�L��'��0-��Kjc���u[������Kr�Vn�s����'�j3���]����֜l�m0�6 'Ӿ|E�6A��	/J\"�m-N>�!�6f���>�_���)W�G���σ賹���)����+��}���|HZ��˽B�A����lR�ݦZ�F�b��������;2��q��m�_w��H����l6k��r�LDD�^���.M&sj`�?�T��=��3K��u��4ʢ���t�7g]9��t���)��4��=���1���rF�Υ��a�i�&��2td�^{��������"U+Uz��%]]]���c�-�] ݤ�y�8��X:��t&m�� ��xt�@��?��
�}��f��M�9k�<>�ȣ�eZ��H�t0M��:r@��ׂ�4��b׋
�P�� �k#���s�}��hr����rO���4���"_�5�Q���1����%�	��X[����}VY�h>�q���0Ю}��xrg4�x<6�Y��uI[����7���->��t�\C�!���;�k��\��(2�T�T�B��AL�:v��C�>���-��o6�/�+a�*��MK�8C[�>����pH�|󍩪��*�"���y�J��N���n��\[�)[�|S��g��{ʕ2=z��*u:z��	}����H��ĸ�m-?l��9Aڹ���x�,�B�|�S�a�m!r��7sl�(Pd̤d&�s$��thl^M-�-���P��ec\r
�@�Ş�k��4��|J��s��-����4y	�&<����J�'*�uݴ8f���m��۴c�(�m�/�~��>�������X��}�6�k{?�Zdḿ�����[I �xt��.]__��ёѮ�gF�z�u�
O�����.I�����n�NOO�������)��:4T����q݋��z�}|�V˵	�X�v�U���c""*�T�T(�JQ�ۥ������!5�MZ.���'�н{�(*F��M�{��'g&y���t��֏m3�d2��thoo�:�e�Y������S���ސO�*R��O�"�f�"+-mhL�B�����H�_;�Bl������{ ���� ?�8c+�|5�9�f3������~H���5�HkU�j�Ai���-YNc�$�� �ƎJ_P9X#�X�A,Y-�������z�QJojx��AZ�M�cd�U�������-!�qJ�@�$�"�%oq���Z���1��9�d ���g4�L�n����x<���Kz��2������A��"s]yF���D�$��)���������<yb�>�a��~Wv����w�����!�ެ���KVO��p�cBc}@Wc�/��R�X4�]�n�~����p8���Sz����C[���HFM�XL��Djy%���-:3�JQ�\�T*E�?�n�K�^�z�M&��.�A �8��ƕ���}[�Z�����r7
{�]BM�]�n���N;�NS�V���}j4����D\r�2��h<�)�R�d���gIz�t��á�q������9؆HB[�X�� 6��2zS��82�.]+�����S�R�|.O�L���j�L���Ö�!B���l6��}���}D�&1�
<i�(�XC��pQ��@�O:��WvY��l�lA,�����X,;FY���Oq6 v�kU�6���y�՞�sm���I�r����!bW>����ȯ���|N������K��-
T�Ռ��@�Κ�bU�&|������.�����^���������G��/��������,|�SG��O�۶���풄v�C5���"�c�ޥ�"�'��F�@���p�	1{ET(h�X��ׯ�����_m�������jQ��2��t���BƁ��/
���y��jT�TLJK.�3`�'� �r�x�v�>��#����^�G/_�4,5�"�����-�5�(�͈_C$�u�]w� �����l6�^�:�����T�T��j���1PE�X,�~U;ћ0��B��l�x ����tyyi�|�����r�g+L%��1����R�ۂ|y�[���#�=�y��!��lF����4����&�d:���V�����0b�P(P�Z�\.g��n�Kggg�����I��C��.�uC�|�^$���u�C�h�
�:6�"���(�PP��0��|����#J���J�j�EQ�A.p��d2����f��w�m��P��:k5���e�`Y�i�^[V�A��%�b����7�|c�3O2+
w:���E����6�;��\����O���#�H ?��3��������tsssǗ��R�v��U����i���'U������j��m ƕ��}�T ��	`b8�w�}G777���k��o�d��a� � 9��"zI��x)�J������0���k,�NަA��'�|B�L��>}JO�<��pH���N4���M��e|��|>��ht�Ư�O�⒳�L��@W��̰aU*j4T�Vh�}��!��,��������!��ڤ��=�F#�������0��{tڦ�әژP�Щm�֢ay�_Ɔ�������kc�$!X�QQ�R6] "��ph
��ri��� g�p��?4���0�����5���ا᳁D��o�Ћ �W�ͳ��~��r��}^�T[l"�3@0L�S�%C�9�Lh�^S�P�z�N�N����F� ����MJ���@����^���u;\U�|�<�>���\-���!���b�������a2����������w��esݵ申��z�֋�T�`�ZZ̵�R��G���}z��=}�����i6�mH�B��I�;���F�lC�<[���m>�Ƃ�3��w����'�����w܋���[�v� ?��y���|
��y�����~�3�N�DD�h4�P(P.�3�`��ÉM0�":88�L&C�Z���<]\\�h�L&CQ���/�^*i.��5ʄ��� �W�.�t�ys�}-j�w�t{��I{��A������ GR���E��u3\8���H�u�S�+�!�}����6ܥ��j�a� 5m�i���A/ⰶZ.�)�"S@��X@^�������C��a�R�^�G���N������D�,m �'#��Wơ����/�lVu��c�@� k�R�D�z������X �\͋�(�L��X˼���͞��k�1p��A ����G�D�wd8�)�	�Y�� @�͔,�K�����hD�Ʉ^�z��xd,�j�"Z�қi�����&��� �-'.�$�&��ēd��`���>]\\���)u�]��w	&m��.0��_�D�Γd��u1&!��%����|����T�]�V4�L�&�6���%���Ap>���b����^�G���tvvF�1����`2�P��#"2z0�&i�0?_�5��}�����|nXl�I��KǺ����6\+[uj�^՘D��3��Iɰ����F��Qܿ�db�i�T�T Vk�O����VI���4N��,��.6\ !ގ�Խ<`4V=�V��ʕ� M��ABH	���9��,����j�2��$���_B�2�Lh2�V���mg�*Tm@?�@�� [q���m�S[d�),���6��tb O�z],4�i0r��8/P`B���g�� )T�:.B'4%�7l$-	]Cx�6_�o��N^�N�Sz��]]]Q�P�b�h�{��$�}����1������NgҔN�.�3�k�����A�>3���%I���΀8�/�t*�����3�k�O$�>}�/��fbog�S� +����nZu�<�0����ﾣ�hD�������?��?��Ǐ�^�S�Z5���=!�,��Q�Z���#���������N&�⾋��g��0$ր��a��S�����EZR�,ld�=c�\.��~IM7KÀ�"�˙����e6�5�?���66i�����o�ǵ����N56�&	М6�-�N��gI2�hA�Es sv���`�xwE	�&��cn������ŏ� 67ہ���MKo�{��p��e�=���b��!M(��ƐkKq_�^���X(V^�\��]�3X�R�i���@x(���u�pk׉w��gVE�A���l1��O�K���Chh�+�v�p�������Q��:$>�V�k���'t�7̶p˿ީMض�پ�ļݵ���_��!�\�Q�)���U,��lFtss���,}��'T*���l��PK���N���j��Ǐ����t~~NgggF��mJ��<}�0�M�f���E�`�M%;��#n.��~��zwt���'#m������rٰ�x^P����5�b�+Z�'M������ָ�O��j&usI�W�Oq�=��g�.�_�E'���΢@���N\@w�X�Ѥ�Fc�C�4��=��u�h�a!�׵�C0d�d��������5ϻ``l��f�*���=�H�.��B�`ִt�Ѯ}���8{>g�1L+-0��>[�CH���ˡ@��B:Nh�Ț���Ӷshۮ�K+���af�'_�3��_�4��p���Cb��͉��.[)|:�fM�y��ŇVU�T��tJ�^����s���~G�咚�&������!��u""�������t:M�R���6����^�G�咊�b�o����c�j&-u��Gp�ƥ��O>�7��4m�6��s���}3��mmBj0�͌�z�6:>�r	���`�5��]�kSk?��@P�[��c���@#�!��ݜ��=��&����� �9q-�b���2q��W�_�f��W�ċR��I��4ħ���&�l �呂m���Rɀ�B�`y�Ţ�V(xp߹���6���`��L͹$��	6:/1`���=�t"eW>��b�w����n�9ͭ�X�Y    IDAT���P�vM��ߜ���|��kW̼�{4������|��\	}-������mpE���
�ֶ�L�����K��ly�6?y�,Sz�={��~���S�V�_��WtxxH�ry�F����8�Y�Z\��p��[F@�����4�EZ�V�I�@�w�V�!	y�6��i�@8/|napvp���t�g�8�����-��s��R��u�&gx�&���ъF	�d4r�>�,_n����~<Wch \4k4ىA;����XG�#���)�$���S��c%ر���kĂ�Y{>+9��Pd�C���&��4�H���8j �|��)�>|]H�9i�em�i��I�^M��u�R?�Kœϥ�N\2�i�?�%DZ��\YX��2���>8�%�nb�	:�����'��&A��Cq��?��0�6$�i���.D�'۵�'M�T[g�ۤ��`7�����+����O#P���G�t:T,��*o�s��ۓ�)m�
����偮�i�4|�(�"�ol��[HOQ[^�+�M�V[��sQ,`��1`�G�l ���}3y��4F�k�!cp^!��!�S\���wۆǤF����dp��m�#�9��k�]+p?������^��S�*C���LHL	�l�Cv6b�WS��Y�i���9�z�d���j`�0���񦅄 n:(�9�����`������9�����6�U[�ZB���~V{��>�:�H�ٜ��on���E��|��{�\�7���ڵ�!��m jV5dnIZ���L��H,��!CvI��;�M��#W�-n��O����0߃������|6 \ ���+z�䉑���|@�B�ӣ��̗`�D�"Y l� j\���H�P�d2�I�=h��(�sP��u%���E�qہ�[�x���`=�h(X�!"5K�sMZȸ�����̟�t�
^�p�_�~ڝ��Khl�榠�~� n�ċi���l�x�����oسB���4#�48�O|��Kf�$�i{�����uʶm�k����z��F�Z4)������i�OF/�ח ���{:(�q�=��;�(d(�.;���.�B�v���N�Ov���F���D�y�1�>ծ.�-;���!	=����_���Cr��p�,���	��:W��v39 ����}��7���C:::�v�mP� �G�������? .�/l`Tc�2ٷ�=������,��۬�ver͟;���-��d>����J��u�\/�Yܺ�����!�z�mk�s?Ґ���*Ű1Z|�H��^m��?0o+�d���yu<��x������,.4��2מ��rH���q7@%鉂|O��Ҍ{v����
�׈�J��j5�V�&����ȢS# 8��\.M؃�h�T���\C@���دl���!�����k,�.��@ԂP��{�H�|�mx�%�Դ�."��|H\�MRY����T��5t��YW�M'�J�ʻ\.S�R1��`J ����%���@8'�C3$1�����˅c; x��*t�^JK(X*!)�Z����m��$������o������� �㠃.��>����Z�q�u� [k8ę�v�C��d.��6q�m��8l����t+p�a��=C2�p�imrpE�x<��xdM.=�������t��N�<�]d�Kӧ=�>��P@d��p���)�^���z��C�ȸ-g��s�2k�6=�y�fwik�չ��K���l	��\.i>�o�i�l�(�]��mĤ�O�k����FWK� ĕ-�2C��Zd��cC��CY8�p�|M��z�n"q+���}���4i0���)}���F'OK��EDn��E�@��@mza�#D�Ukka
���*�,�1���b��K.@� S�3�������B�`�� h��5�vS�1��;��6=��X.%�����w�O�6I��qq7�Pv�g���%�i-QΤj��S��Cg���(�p���wY��.J|=ۊ����a�4!���|��,�lq�>�/Z��&��m��GQd,�ņ�j�K;
��>8��̃<8��:�!^���Z��u%��o��Si��]Pf�Ks�B��B��]����b��\�����.lV�- \øڙ�[ӡ]�]ܿ����&�<$qM�}�����l*��F�A>�����$" ��`@�ᐾ��[*�J���s���50Z�>����T�a��ab��k���ܾ��B�|�4j6���
6�ҿS��yR�l�,L|i=�׈����|:�R�|�d�K����IP4�`��ہ�m�Z,%�R6#}gm)drS��N`�m�qW\�\�Xp��,�l�6��(��������ͻ,X�� [M�`��!�j�!2P�2 �<`�@猖���]���x�ID�`WPyj���+
d�E<����w����?O!�;�9Tؘ}	n��&J��&��y�����KJ��&do�[^[�=D��~9T�É>�%"�N�+ ݆��Ul�pT���:�x���Юu:z��1��7��ǏS�Zݐ(�����ɘ��/���ƀ\nr#� v	p'�	M��;�.�I��X���.����_�F�a .�O�m����� ��׊I��+�|�34�`��� �p�*��v]8�L�}r�]0.�i��䬭,ȴ)i����wka��#o����p6`����l��w&�A� �ylP�P�+��$�D���m-aO�IM��>�"c%��������O-�!��h*���`@�^�8����y���{�3A.�tf�^p�X�s	��=�����]�Mn��%({X�]����6l`��\���t�Ð�}������8�N����_������ۿ��f3� }~�6=�M{뚲�>�m�1m� m�r�L�V�������t��=����R*���jQ�բZ�F�f��������/_���m[)xohm�u)�d2��hd\�ժ����@�QZ�v>��J�B�z�0���eU+?�l�C���,%��g�L&f�G�o8��;�綵�%�٨�l�x`b�Lq��ߏ{�	J�9/̸����f���,�O����%eK~�"�,ֆOB|Sm V2��@�k2YK��Ӷ�B:���'�ÒJ�(�"*�˔N�i4�p84�4�N�zMx���z���Ҵ����$v�qm9L�� �2y�-�V�[��J���b�0)t�Zm#�
%��~�OWWW4�͌�8"���n6�5g���f`����Hmc�m�Ӻ�ں�ki1_�`8�n�kֆ���X�Bbp�9C���U���/���I������̪��C+�jߖPdK���۶0���Y4�"R��d(��Q��0	6�^�...����ڦqZ�����VU�ۥ�hD<��?��>��Sz���j5���L|!"ʤ߲@�B�X�`c��$�6����`^�T�9�0\��[�����ѫq�g���o|��>�>��3���;Hp���L�S�Ft{{K�ш��I�CqV(��S6��~���k��תğ���(��>	s���?��wm�V�/���S�X�f�I�j�V�u�]T��M�v.����S���o
O�.>��������%6ZK4�Mr�J��3�>;2�Y|N/.�5X�j1K���{�+��AΝ.0��sD�� W M��	�/
�8�6��d�	�PV�e�&��f�7�EWWWo��	��+QawA"�J�v��B�|��7<�k倔(,C�d}F�����Jd�!�r���1Ϸ����bAS����V�E<�Ǐ��^�G����&\��W�\�����|N��ݣO>�������~��_҃�\.o����[ݰ�Z����K���jQ����c������3����f�I�J�6�O%ຆ�d:��#UZ��p��f����pW�\�s�f�`�R�P�T2�Θ��t�|17��3C��j�mK�.�ِ�,�\�Uf�k�c%���P�Zd��u5�N�P(УG�����nnnh<���9-j�ZDD��L�R4�L�}ĳ��4::� ?k�5�
���>��=�:l~mVS���./�P�$7�N�|&L.�7�"j6��Z���jQ�ݦj�JDD���H��^���鍢������8���׵��b�>��C�����.$ ���d|m�!�}�kg>�w^eC)v�{Aȃ�'u�GT,7O���j�5�t:���c"�at�u:���kHD���Sc�&��n�̓�[��Ʉ��4������=x��>��S���M<0�-��������I��؅�mb����l@;�5���턭��۳�C�$��;NT��zG�G�#8I��N���`à��n�^]��v�M�^�noo7,��(—`Mz�n�Dp7�%��ei�.�+�h]Q��PR�g�kT(].�&µZ�ңG����NOO���^�xA�ш:��z=3�$u��g��b�B�IE� �%U9P�V��z��ӆ�d��5KD�K��w��@��XS���$���X,R�ӡ(�h�XP�ݦv�m�ϸ�-�o��|޸4���.� �W��d>��oS�U^dK�ʟ��oͿ����gP���b_�Hl�ݸ�{�/�T��(���l������M+gP��ڿ�b���6���?71��r�^�xAWWW\�E�C�<���|>��tj� ONN裏>�G����1ݿ�����R��͑;p=+�����hdXa�w� x��S�V��舎���^��v�,�k�Ӿp��6��4�hL�Z\�͟�}�\���}#{��Retg�V3����ap��:��uc5�^�i8�t:��L!2	�%���:8mј>��c[C�|�4!�v��k�jZ|/�O U^]]�`0���S�b�r�ZQ��3���v���y�h�q�s������߶��'Yw	p�n�m>�V��"�]Ѵ.�k��"$M�V+j6�T������0�{�� ��5�b��ą�x�.����k�<������f���t:���.�_��O_?���U� ܌�h}������Ž)�(ō�P�X4�U5� p����홍ӱ�Ʉz�����lN<jQ^+0n����?��c�կ~E���o��?�v�mZ� � �< ds��xL���tssC�^�������tJ�t���6}�����#��ߧB�`�l��Ɯ�Y�t}6m��O2��4�0�ͨ\.S�Z���CZ,tuueZ�h[�R)3��8#e�[RΎs�5���M��^�sʶ��`�?�*���D*�Б�ڄ�,�]Cs�癇w�υ���rIggg��g��x<6�����,�Ʉ��y�p!IZ.�EU*���S��-eWqץKB�sdS�HO�V\�VL�mq�=C�%�H�x�`�V���=*�˴X,q����阽��A~���Z���j�p8����u,׏�Ǎ���kπ��Ù�s��%R��>��������5��?E��C�
uJ�3|�h��6����������d���ʲ���!�����q�x��[tpp`��ƂX�L&C�v����%����6�_����g}Z�����_���_��NNN(��)�P�$ ��}��5��/�o����ݮa!0��떑��Z,oX�F��߿OGGG�h4�F�s�ik���;M�n�]�i}08 +�
��mt}}m$)`6nnn����	8E���Z�R�բj�j���������{2��ƜI�P2�!v7Z��{��+._�6�7���v/9����0�r����SZ,��vM�h4(�Jmth�~�����r�4�>����U���؟����I糱���M�#�Z��ጡ���"%D�?�
��C��uj6�tqqA��������h���g2s_��[�T�L&C��ߧ�nHP����P�!��u������p��`�8$r\F�K�O��~bn�簸!]E'�m4��_��_�O&��	z��H�;&��1hI�A\�1{T��}�}���t��=j�ZVK�R�D�T�l8��j�J���@���JG��x<�B�@��������~������	�j5~8`AՌ�����Ћ/�ɓ'�׿��nnn��Y�m{�%����(��h�\��.�?W8��!�s�=�>��*_`,����t���P�ݦl6K����U9�h>����"��s<�`0�L&C�z��������<˰���^<.����ŀ�6�A�fY�b�� %����+�E���\ގ��\���b�hXzޥ+��_`��g�Y*A(��(hP(��o_��V�ɟ�1��Y!�})d�r��d}]zz�=�i�m���*.�K�F{(�"����$�Ak��f��𐎏�i:���ŅyN������.o65�����s߿��] ��� �y�R��m.#���(x�;ndq�����@� ^R�r�5���v�N��[r1���гg�(�����8C �`0�����(Tl��j�>��*
���C�F�d�m�����f�^K�J�BGGG���o�[T�h	�M�+�J;���3z��9}����_����F�ߕ�����G��æ�Ar�L"�O�_Ί� �1�|�v��}r��,YE�[	`�������>��#�������T*T��(�J����	���:����!�Cz��a��
煕oM����}�s���e�k�E�:�n�T�Ϥ^��/�7@�[� ��v������l�-��젷�`
�$<��2�O�k�4[����|���0$����p��� H�Zy=5�aP���!�i�>>dX�{��N&�4)�J������P�X���+:??��je�K���k���z�)g��`<�N��^Kf\#�l��t_���=�y�Wy:��t�M\o&��b�h!...����t}}��7�")��0��rߥ��f�T~bf�Ѳs�\�,_���aC9��J.�=��rId��u6�ѫW�h�\���!U�Uv��*��k�F��i�(9�E���Ç��Rr�+� �%�\�:in	�:@��r��v��o��?���_��_��W_�I]
\k�K1>gUr������...�����x���/���'�x�E&�O2����Y�Ռ���l�׫�jtrrb���"d:����5�C�V�U���G.��H���3��+�b�&�K�=�Z��|�on1&d��/���j��e6��(��޽{���#*�J�8��������T��42!�����6k�4��z���c�ي���c�I
4p��H��u���P� hmh� ]��Z�[����G�ѠZ�F��ǔJ���˗���SJ��t��}*�T*��^*�LW]4gC^������{���9�O`�i�N`:��t*���wuuE/_���ϟ����!�B ��wu�4�>����Tp���H��!Ԑ3!4��pm��!�S�hZ[kk`��M��x�>��3�����S�T�L:C���H���pK��r`�r�eso�o��y?<�`�^�j��(��r+\|�C��d����7�|C��_��/����3�w| ��$���7x������%���?Py�|18��p?�[���ɾ�=��G��I���@"o!��k�T*t��=���3���zp "�������ύ4��ϊg���9H� 0ɺY�pp6�h䐐khH��#�f�&��M�:d�b��0���tttD�t�NOOi0��<�R����v�t{{k�(���Hz�����d[��!d}�:b.���!;gqD)'�Ǉ�|��UعZ� ) n9K.�?��S�V3	��������F��%fX�x}�� b��v|>�����<�������g!����t{{�1`"M�y�vxw!Ox_���}_{I�14� �+�8��I@�ms�l���r�B*�m�`0�/^�z��~�O�ٌ>��S�w��)[��ۺ���l�flr\�@�?�F�7a�</_��'O�������/���ݫvv����������g��d|���  @�۲e�YZ���:ـM(����t���x_�R�*�
�Es?��io�Ň&����3���&�����t�?    IDAT\�)�/f|��Z������I_Z�y^l�ul���ip�=��l�!�y�]��x= b��E�V�T�V)�˙ �S~`���;$�7@.˱E,��V^D����*t�3�6X+^8�+�����$��"y��X,R��7� �������b�F��}t�O,� >p�ywF�w�q�|�}Ŏm�h�:�+� ���s��d21Cx�>6ra��t\����ލ��]�[Q�薍S�$����N,��l��Uqr� ��tJgggf�P�X����7ia���FJ��!�M���	Hd�l1g�A�}l��|�����~��w�Y���]'�I0�1#8 x2-)��u������������S�^�*l���5���p*�xW�]__���9�~�X��͍�� ���N������)G'�6$.Zunkǻ�0W�-/�B��B62��I �BY�9W\�tkL
f�Q<�QQ�ݦ�lF�R�Z�����y.��4�V�Q�R�J�B�j� �g��R�wց' ���eql�	I�϶�^�[���c�1D���z*��T��6:b��.//x� ��ɉ��[������O9��A-(��㾽�U�C�K�z��/??��������w:��m<7�Ʉ��>��}Ѯ�P�!V4������:&>�[_�^��H�V9��lRW곴������ ��
�H�bb���Ҵ�r����'ݕ���i�bӰ�k`�2r�'^�C���d����^�~M_|������?��Otqqa�CnQ�m>��vM���y�G�����M��50��]>t�Zo^+m��!ۤ~�C�(�LH�?��3�����_���ݻG���D���}���N�|�Z���yj6�F'�� IW`��hB�b���gX�|h��"X�=i] ���{���s�{\��Q�ף��+����j�J�L� ��bA�R���an1|��_*�(��R�Z�|!����T<��'����ׄ��\Tl��KslgF�!Z�<��8�a������z����:\��4�M7�Ȯ�9���y�8���kY�C��8d����ʃ��>M1�<�Т�{xwi�J��>i��'0����o�D�\oT��I��C6Z)K�5N���ژU�l2�g�j�JQ���s�V�f���d��ԬP�-0=|C�Z\�o�0;�~��a������qSHZ��j������N�C�V�Ls�Q���ڽ<B��]��V��d}S���#���	d�T>;;���KZ,txxH�F�0:`�`uss�&z7�6N�R��`v�, ��o\��sJ���?'�\l�k�ri]��Rg,�4\�X�^��Le�	�B���$���ij6�frk)X�a��zM������)Ҹ�\&\�m6�q�8��f�u�!��zNz(��L� p���������͍!!�p��]|��`9��5`N�A��'��x�kpAP�����w�l�.
,�Z�	�&���-�CH�8��%����ȵ(��	�i�]U"�;�z�|�E�>�왙�-�����E��m{oh�`C�V�F��s�������ӟ�D����MO�<��/_R�ݦN�C�\���is'eX�m��u����n�M:Z�܃��U (��7�ǚ������-\�Չ��;�z�N�J�0���E�~����yNj���o���1V:�T�j��a��m�`�P(6 ����Z�>�C��\��f�gq�v�ֈwJ�%�,�$���8m]
ts AA��5�6��� �OAD3@Q�P0��n׬e6 S��l_�𜸡.o�8mȸ�"��ڵ7��,ZK�0�?`+�틢�M������`��p�0"2�v:���1֗���hʵu���q��[X����xGS�=I�|�uێE�伟�m�b��,I�ﻷ�mZNڦ�iVC7\ͻ0�	�v�a�1�I߃l�ٌ�={F�b�f�u�]�����!o)IF�R�zy� ��V��Q�U�zzzJ/_�4N	�~�-��}Ì�_���C�lm�'�,,p:����P��1�T6�R�7�8ШA����DDk�I�k����;�fNDF�� ��v�{�.�����v������t:m���hD��.//�����(2b6�5A8!�iU�@�!�E�bm��Z����Nm��E��P�EY��ß�f�I����'��ej4���s�g ݌��KS� ��	�/f�g6����w����$>�q��4,[6}���\��g�`k:�6Z��|N�f�tcP���}�ǝN�f?��O�`FL�b�0���[���E��!4��vvK�4.�{�Y�AY>\fs�О3� �kPvWV^>��k��H¿������j�..��+nl�W�_�V�e���Ћ�[�\�.?�̓�v!|�E�WA?@�d2�����oKϞ=���3���g���O�������MkQƅ��W���y�����kz��)����?��^�zE�~���:�T�-���0�����2�,�٬	5(��2�~n����x<6�ޯ�z�-��Ҥ��B3�\.G�JŤOq����bA���h�К�f�&���WWW �{���}��j��U{`��tB�� �ﳻ\\�P;.В����Rs�[�6 ��Rg�]�6F��,�j5j�ZE�����dB{{{��Ş�ר�jtpp@ggg��ߚ8S�k���p΢��Zc�m��7��bhC}�]�r@bӓ������.¥a "�7:�Qpop>@���	��cO��	��ћ�_,�F�K�m�b"$!44�N�l63C�������s�#��!��I�J�3`�f�e��o���#GJb�+i����b�ʺ>��ɳU�!S�����,n��ι�����������ޞ1����}؆�d���,�����k��g��?���={F�n�0�I[��� �^�7������r@�A$��q=�!�V.[%�u�
��`VN+�
M�S��Ļ�xlr��&�r9c/�7i��f�-��&�"�&ʪ�0�X?�Х����r���~�s������n.���Et�8�~[ޱ)
T.�M����xL�z}cf ���r���r��x��o���րͶ-�^�b�B[ľu�$�J΁@[�uޜp@0�`)�
�I��pC���t:5vq`D��4�iM�"�����7)��׸�_��Z��Q:�6``���~�NOO��횿�Ś�9�������Ǣ�M�e��˲��	����em��+�Z���6 o�hm4~0��,J�6��J�(k�Ip�Z��Ʉ���Ks�N&z��5�7@��l>��x��.-�G����U��bAWWW��W_џ��g��/�o��n�KDd6�m��]i�^�����t}}m4��p���,j�٧����E�c3�y�<\P|������Ft{{K�^���5U�Uc3ĵ|(�L���E��Ʃ�CZD��5���Z*�M�dk��ATάiʶB��������-_���pC�^�g��l63�'Z�|r~:��<CDdl @��:��a�� ���$@W���u��u�ѐͷ��߯gn�ǋ��rI��� ��ril��,��c�f� <`����j���L�;�cy�]A�k�� �Z���h�
��xL�_�6ô�X,����s��PpW���������q:�����@z�k��s�]~�<���v��~��
k������NS*�h<�_��W��r4�ŋ��t6�4�k�HI�Uc����tzzj��^�|i��`2�h��'l ��k��vf�V����⛞������f�KK����a��	]P��b� l3��� �(�����?��-t�`L��4��c����Z�F���إq��v?]��z唾O�`+�nr��Rx���ٗŕCh����\"W�<c�?���px�=�f��3:�r�LDo���=�Bh�˥D�@Ist�M�kr�]ʾ�������u
q�@�{$UX�(�P����E�T*f���:�"��jw�����E<3l�R���9ʤ3��eMR%<�m�=!҄�9�*jg���H�C?h0��K:@������8���X�m��`��Ǳ��ڄ�E�rq-�|�	�P�f�����3�F0�5��ٳgtzzJ�F�X]��e���ňڼD9ȓl�`0�W�^���9�z=��Y��P��ԕ��� ��ꊢ(���c�ƕޝ���&�\q�%Ӗ8;�Ԓ��M�uPrk7LUCk��l>��%�/4|hC��Ǔ����d�ߧ�k���	�0�b�jj׎w]l�>! 3��v�j��Ŷ��O���̙X�}�e�`�( NX���� ��|N�r�<#�T�F����V��!�c�k�bݷ/�@�6�W��d^C|�C��8�ݖ���t����hDWWW�X,h��g젭FX�������[���^�|0��� \R��6��1�|��s�K2��������uu���%	�q}�� )�]�� �1��m {�����6�� ����S��A�Z%�V\!7F�i�L��...���*��h.�H�����v1<�+b� �����2�/�<a�;���= ������`Oe� �ϡ1��x�j-M���-�K�\	Z�`f���Z��B�h����t:�pM�5Ѽh�2Pr�Ax��q���#$�� ��$�����؜��=�.{���sk@�oXq>�ݣ�h#�y�\R.�3�n�p��յɺ"rC�xW��/eL���:_ʑk�s�?4�P<{ �XÐ'LgS3<FD�ȁ-%w��	�h�= 0�̠(�{���p9K����Ê�����#���;n6�ʤ�� chrỔ?�ؾv����s>Ɉ�����]�r�mF.��m��q 1o�s��b�BrfG�x%����vp��,��f(cx� Yہ���g��]ǁ��>Ҥ��?�Ӹ�Қ(E�L�v j̟l�p=xH��` �6��""z2�lj�B� Z�g�a�Pj��� �eu���$����R��Y��=KoP�4v��Y��G��B����g?�<� �x~���d���o�/JE)�g�4�L�F\ V[�.&�ОA[�K�q��F�J��/�-���^�	XH!e�C�����p<��im}쏚�� ��=���\��f�y���3��%!��MLu1�!��q��|�5?}m��K:Ԛ��K(�g�z�K!�ڑ�P�qZ6"2�6)��j53��2l�4�L��:Qn��m�8[�ߧ�e܅	�KFʞ�mh�Z��Gу�Z�]g�qxc�V�77@G[�oN���؄���g��(_	h�x<a��l`����t1X;�]�#�@�X,n<����(j�r'�"���Z�.������3��(��iE|���2�",��k5[���O�z�X&��A�� �8<�����^���y�\��q������CBC\{�,�4y�Ow�ɜ�t�3������}���F���*Dd�Zc@gG>���J<1��Ll�j�)z���A�@���3y������p[��J�h�!����p�!�v�V�ܕ|�T���Mg��b�Ѵ��C���8������+��r 
�>��ކ2��4��w-����a�CB�\kl|��t:��t�T*�ajm	B0���a�G3��4�h�1<�&!��d^�9�v�K�| )��� �[�q��f�7.�a@j�]]�8�z�;x�#����L�$� F2����ԧ[c�Mb[&MY�R��&ȡZ�]�x<6����on	�NF>��5�'xe�YJQ�˅��=�B��q��]A*Z���z��ې��}笤��s � ^d���N�9I�� -
���s���o�>kĆa�X�|>��phl��!���;�/\���
�I��}�$zO�l��nC0Lp��nHafs�
�_��Z���M�����o�����d+�[>�r���}>mI��`��]]g޺�Lob#�0�g���1�0���j�3_�헫�+;��c�'�,9k���%)8����`�k45&�:�.�n���\e4����������M_�b�3�}F����ir�� �͓E! �L��i�Z�r��pQp}܈u9�)yW��K��j���I�\���� /�ý<��&w���9�~y�]��}<�� �^�:U*�=8�P�q	`R�m��А���p����6��&��u�}z���F���ZE�pa�B�\l�&��bD�h9k7�N��5�n�In~�`��mG��t1L�M0i�K��%D�6:.��4��f��ͼ�s�A�T&E���.��q����l�\zFZ�@s]�����Xh�p c���b_�(?�v���6�5D� [�!�rx�y[;R��e�]mH�j���",�9o�j�� ���Cy�Z�b��S �>�k�k��Lx��;�$��K���HFk�� �^b�"�E:B_R��H�zk|}����mKB��*�"2�q.�3�Ҝ��'��� Iϔmֶ�>���wݕ��|ټ�]��. ��΃V]�m�%a��0'6{*��-��lm Fz�����sS�8%al5M��b�e[�d21�6h�ʉiC��_&����,��{�՚h����	�m��5��Z�������	��j��s�״����*^��-��5�͟}��3�wh?ρ��|����"��B-�|zO����j��(�K�u�`mQ��V8g>��J�*N4i�\��.����(�زP���{�� ���y��K���6@�g#	g��(
�2R��db�2�����	�\w���}$MI/rt"�����������F���:�ϩ��������`+�B���{��Pih,�o��/r���Z�4�����n��g�i丯��vUYq~�m:��&���B	���A�k����>��9������9]\\����џr�oL`Kp�����1��'rW��@�m��p� �̟��&�k[���s �q������3�k���x��BP[���X:�B�׿6��*rCXY��������L��f3c��Ӫp/1��u/mи���̹
a�������\h·M��� 0��z�HZ�¯#�
P�X#�����4���B���9�;��h�!C�ۀP�v��QQ�ӡ�����7{6����e2���2@Wv��@������ǽ66bJ�Q��?9'�]^��J�2��"��ǡ�nC��)�sqdUp�孽&X����������ݶ���zi�
��.//������u�z��|V�T3�l�wp��C!�?jHA�%h+s�	?~�-ښ��{-�R)3�ͯ/��`�-kٺvM��
Ai�_�3�Zj;�m������SvH8�k�B�N[��.%D�֙L�͐��k�3�p�����p{@���D!��Kh����hRF���s�oRr��<@@>WqI�� �{��_����P�?�;�՚Ɠ�)p�lH�}x=�:|k��]Xg��E��V�T�VM(��(�/..�|���h�QR��"Ζ��)����T�q5	�?q���}5.�iۗm����dC7<8�`-o<���v�ƹ��?c;T����xiZ���č�9���2ý�j��$��f3��zt{{K�~��[�6����^�<�]�I�p���BR� 1t�-���z=�v��sCW�(^���6�>�f�|��Ҙ��a&�c�Ɯ�
;ĲG&J	����f�&�q�e�[�ɐ�.M�ȥ6x��^в����3�#�]�x|�T��hVZ.�F��u�q`b�]�L�����@Ӷ'y�q�6^�a�=.�?��,�+lH�C���ʮP�wn�{��wDd
:�mpo!����|>7j�����!2�]�oq�r����bN����N�Kұm�A�����l�/�/����d	��$wi-��-0��|�ti�|>������=��i���@��|��dp I�L&D)�R�D�Rɀ	0q`J��$�3q�g0m�����`0�~�O�����hs�p <� q� ���e���\�V�=8�ύ��.�N\k�������kk@�e�oך�Z�q�S �#������qh�r}����^��r�}�C����ri��`a�]��rɹ�<�6��׫漠�|=b`��x�Ϡ��{z��2E��s    IDAT
C���pH�r��(�z�nbxa�ƥ���]�u��Q|b�'4��s�~�ta�g�x{y_�+Fq��].��V�QEƿy:��{Y,�T*Q�Ѡf�I�J�<Ӳ�uu����=#�����znl�}>��Z���î���R��K��G\e����%ʢ�P��H�A�.��(�v�m.��D߃f� �m/M�w�[3K~x�YК���f�+��w ��-�K����h�X�C
h�s�	n�����5���>����9�&�	]^^�x<�b�H�F�  hpe�ů�n���0��L���	}0�PZS�����!���Ym����kVR��^KF��Av.$�����tr|g,�^�\C��;g-y"!���2.��`k �q?�kpf��� _�R� ��B�8 ��i��#t� ��ߞ�f����	� V�z�c�u����I ��:��!>p�_g,������YH���6u:#9��� ��l�j���WWWŮM���F$e(CR��\_K=)��GI�����O��\Q�I>CH�;kc)�T�>�8�.m?`�>L>�ZȆj3ȶ�pC���y��T�.`lK+���� �W��ju��KI%l�0OG�~��gj�mJW���`�5-�Jf��X,��{��{k�{��?�N7"]���X]���IӅ�LJ����L~�l6V�y��������M�J���l�lk���hA�֩"�/g�5��/t�}��#��uIAl�	���BD&1�{7sv�b5�_�������,�S���yj���`Ȗ? 2R��[�,�Yp��>�!"y��J�B�V�Z���o�DG�/�{��rn�yB�md
�"���3�Xq����v��	�a�]q�K�GK�T�qZ��b]�^�dC�I�]L��l~�4w����U�"�u6��r�L�f� �L&c�N>q,cW�5}�#	`�����A"o!km�8#Z1"<��h4�^�gL�+�
�R)���6�\c��
�N�����p�
\3D��1��_+�$���~�ӠxW�>��b@�P(V\~/�R��y�0!o�ˠmmpM/��<�7�v�~Gȳm��7^<���G�φ��(�(���b�0S�\ �:u���&غV!{�,�%�q�A|��zl��6��eL�����z�jC^�r���?�.	��l�٤R���Y���3�Z�tȐb\�1t?p���\�wEms�v8�\O_P����{�-��ns1]����Ɛ�V:hr��6�M��N��%
���W�.m�`RK��B�W���O�s �μ�倐�A�gߛ�Ww��5�:���^�g)6��zm n�բj�J�f����iz��%�;q�\�����z?���/	�q����*��c�-I�h��xd����� JF��3yA��G��_�hRt']+�f�Yd./@;Z[�\��<g��g�&Rn��=����2M
p9c	�8����
�-^�bH����u��7�5��Wأx��?�`d�����ܝA�oP$
���;Z��Da�l�ϧ�vV�aި�V����;߰>P�p���[��e�ȸ \�k��y��K��Z��g��pp᭝ܸKܪ!�p��4�����\���]^�2�G@{�M�u�_�ơ]���9xu�-�0��:��7-�^�gx�XK�+)��ؔ��8�ωC�i>��r���1�����`��# *?"��@[�fl<Io	Ǒи�$���%l$��5�5��w"�������}E~!�.��V2���Iy�E@,+�1�uEF{�� ����4e�o�"n=�,\@4TsșF-����B�X,R�ӡj���R��=װ����6���gtP���JM;n�>(渖���������_9�4!�x!"*T�T̀פ�pR �@�4�͑(�����\��?�\���U<ۊ�8��w.��U6�@�\�I�@� p��d_E��(d���ZK2n����Kz"����Z��F��ڃ�P(�aA����4����ZSi�j߆��lL��Q��o;�v5�r�lLfqH��0 � �1� �`���Z�v�lA���:X�\jq�Z�� ����o�3�<wwՙІ��� 9�+ �]@S2�҂<xM^��i��4�M�u�-|Ci��jLO^��v����o6��J�B���txxH�|�nnnL!0�LL��!q9�g���W�`<����B�
���c3C`��Ժ�\��eJ\��[���y�%!�D��j����Z�R�Ӧj��a�(;v��O�S��l7}����,��'��$L���Lŕ�m|E��^emm���6�-�e���@���7-=(9��+P��m撉��B�5B��`O���7��*U{\W=�z�ʴ����k���"V��Z-3�{{{k�I��N��/ߢ���̻ ���E��/��h��V~I�.��Z��g�nض�[z}��h%����E�n��CD* �|>�Z��C��]��j���Š�3�KN��a 1�� 84P�!5�mc84�L�R*r����h4����߿O�v���C��IM+�,H���{���p�>7R*ͺ,�X(v�E�A,.7�]*�*!�Jx ?��\>pӰ��y���F<�r9*��f�����+��4 �s�j�h�.q(빋3�}I!�D�\TJKC�\$g��`"�j��h��ݴ׍���b�B/��J+�3�m!�Z.f��. %�M��j���mK�]�qi,D\@�� �x0�L��K�1O'�d2T������0h0P'"#	�ID6G���w0hE@�h42��-�"*��[��4���S*�L41����'���3�+(�g�l.J�:R 3��j5j4�� m`�E���-�c��������j�h៙?o�^�P�A�����Wy 0n�jƝ��l��=Ac��v��*�
���Ї~H{{{�����S�X�v�M�\�z����l�6�g�#m�ќR\�P!=���tj�"H3P-�4��7��|����k�y��p�%E!���_�c���M��ǳ��Z�V����=zD�N�H�xG@^��J���*�=6�����Rm�?��:�!���.>��Ij��/�~�������	�R�9� i`����|��ho4�I��>��@i�o���ed�*	����
�L��.i�z�Jl����e2*�&ƑW��upXB�zpp@�\�0Z�����h8�h4���x�a��cS �/��������l.k����wr���g�~e�����n�!'#F9K�%�� �!�����J�M�Sc�?����)���bLC,}�O��y؅|�q�s�g��Y ��g\��iA����ʩl�5���{��Itx8!@s{ttD�N�*��y����J%:==��V���;	��u(p�������.�% ��7�{����oᓍ�^�����|�`��f�I'''trrB�FÀs�I���o\�(��\.o�;���j������M���ٶuFw������f�:����c\���ƵSMb��m�q=�jp���ir#���m�#+q����@���X���ed*�vml�#��$9�>��셭8[)��qТ�ODT)W(*F�Τ��d2&H�\R���؆<�����2�@2�6	L6�ݐ.HY��8�8k�U8�6Jn��P�T�����2�岱X�%�J����Q:������PG��헦.FE*����ac>�
b=�X�kqY��ܒmW���,ۆ��g�dS1�l6�������R��g�(����e&onnh>�S�P؈���R纋�]�QP��fht������Ł��q����vو�$�
�{x�Ѡj�j�*db�� ���k�ļ`�H�|ŻF����Cm
��Bɼ�"7����7�]�����~e�08>0�p!�."Fml06�*ddK�����]��&���&��V�fIFk��A�6`lj��a?�,���y;���h��o��V��aJ��&�Í8L�*�k$��T��3�T�^����#���h�� �dlZ�]�G[�j{^�;Z��v�>|H'''T��)�N�S\Oo��Y.�tvvfbk�l���$sq���8��P)*Q�\2����8���|�Q�r��c</�Ce̑�4 �G�[*�hoo����C�",Eh6��\.������yN���g]���W(��m�d�E+�\�c{����b_����m��He�.E����rw �b�0
�L�:�IB���ϧ�O�#���	o�M�'`��R!�G��pq�g�k�<��}�pq<'Ct��T��K���"~�`�%�ȸP-�-&�Z��thchrO�"A\�!}�5P�����4��R^����= �|>O�v�Z�uo�&�W�,J�S�j������-�JFO�-����| G�o�4@��ي�m�>}�_nJ`.�|ttD��ߧ�c����שT*����5����h4�{M�
�����gួ�l���xV1y�{��q`$58���n���.��L��-�K*�˴��OGGG�l6i�Z�-<R[���u:;;�^�G��|C`�*ۦ8�s��s?Ox���F;� ��Y������dC%�L
(����X�T�^��c0�6+�$D�RCp�.Ȱ��E(&q� ����".f��p����V�&��$'M)�sM�!�����\C�|]ӯ>�I��Iz�>���U�l7�%�vX�
�}�9q�%8����4h8nxKj׍3V8�!ʿ�P(P�Ѡ��=����\.G�����U�.ن��ig�f��5�RX���Ϭ9r��ە��ͪɗ��5"0c�q��f�I���tttD�F}��](Ћ��J��)��.��ܘ���jeXӤkŶY��Z8��^� �ڳ�a�(�6<~Q��,�;`��=i�G�
:>��Z�M?��L�yxxH�v�
��F�;�X�h��,������z�u�v`C��6��R�r��ɡ<�덟��r���M�%p�s*T+�=��ehhK�EQt�|��I�C%p!��l�f�C��k\�!p'A��>K���sO��j]�Ўi�Pl��*/�v���Ү%en����3��@N3hC����\��{�B�ҡ?�i~C�(s�j<���-]__�`00�F\�)5j`}�&Z.����...����0�\Ϩ���B#�)��|o����|���b����i���揄/YK�� m���n�Mv=���0�������N�tyykO	h�ChkQ�����LQm���{�k%�~m:}<X+��۞��oC���E\>��N�C��Ǵ��O�BaC�Y�dd�(�f�I�v�ȍP������4�{�T2)l�{ }<w�����6�~�[�EQ��;)Ew ��e���yZ�
�#��"S�l|�k`N��n����Y�CNH��/�-n�<�y�DZQ�M�������&���H�|�]���󅶍����2p�R�*���r�h;�'�fm��2�Ʀ7�N����z���`3y�9� 0T�2G� �\.���!���Ӌ/���n�6��o�!:��ʵ�R�"3��Լ,��k�vX�5m:��{��\M��'R�0tׄ����rw�p��,5Z.���������.��lirh��$��ާΣ^�ʍ�{b������ؓ�C�<0�p�.׀�AÆmUh���>��D2��|�K�KI��ޢh�a�#Q�6W&W|ߊ/��GG��\ �=���PN�1�N��Ī��N�k�D���;��a7v�k��95:`��sN���F�{_�|-8�}��WWW��o���;�V+���A�۩��'O��e�__��{����,~���k��g;�/=�)ݺǜT6������;����5����K��U��>�=��8d�ul��9������C�/�����>�������x��	�H��4���c%�<j��}����:���)��1��� ;�=�Q��X,�u���{���Ư~�+|��w����A�vC��!*�����_���� ���?��o�}oVc7�S$��E7����A��HN� ~�C�=�|V�*�>��sNF��Q�p����r����DQ��z���[W�Lө;���`:�����_ay�ħO�����^�c�{����$���_/]�1��ߑҴ+u�ؗ�6օ;V�����1yB�$x����/�����}�v`��ׄ�O%�����_��i�������'c׵���Υ�v�ê5�X��$�|�/{ӂ�wa+t�9�;���必�t��.�Q�ym���eY�ӧO�����Ç�u��~x���>�јG�X��о{(�y��<���?���?��D�P`Ʊ��y�c����Ǭ��$��E���c�������,�>m�c�v-�SI�ZTotH�<�����n��=&�r߿�j��"�s4M�?��O�O��?�o�qݞ�t�` �eZ�v���Ǧi�_���+�
<>;�����C�7(�[�f��[�X���r�N� �1uC���|�e���7�2����4���ﳝ���o�ů~�+���?��Օ#�czԱ��<���w�b]����{g)�2#�����?-h��W{+�$D���(rdA;eV�.�Y�����1α	���kIV�����_������ӟ�y��(
��ѓr�>}6��g?�� �j����->|��t���޿4to���{�>�����ﵮ�l�4���dg�����߱���$�b��O~��}�օ;�����"����?��������������{αn�AP�\����C~��z��zn�s��#|O���&�>F\�q�xJ1v��r,ό�.��z����c���A�ֱ�S�����6��<m;v�������?�ޗ.��x(�������|>Gx��;��PQQ����kl+�`���i���5��wǜc׬��:�-��7 n\�Ծ��Scѕ��#���1]9�D��΃w���z��2���������o�����N�:��] ��
�M�,K�z~��w�����j�:}<*�K��]>�����ڙ{�����;�7	��ɩO�1���tm�rZ������}�~�_��o��|>���;�P;�<�1��]!���;|���>}r$��o>�d¿?�@�n�%��',�R3���t:�\�*9������B�)�C��E��{{yy����'��믱X,�Z�s�n $����_�����{���n��E�s�Χ�H}�����t/�wR�Ԏ�҇cNN�3Dw,u�?����S�9]~R�)$w�xJe�9��S��9��}]��,RƎC�q8x���1�v_��Kl��ń�7P]�����{�����{s��/~�<rg���ͯ����ܘ���}�����[|��wΞ�CL���1։���>���Әt�㤽��;N���ǁc�f�Ώ���
�}f�H�1o���sӿ���7�|�6H�^h���؉�o�d2��7o\��r�D���}q؟�&=f��R����?�9� �� �[v~������=��vr�Ҏ�Ҽ�k���������߰ R��E<�x����2�E��!rw��X���[&�M� ��O�f>`�U�R%��&q���3�5\u$�-��K���B��E%
\;&�����������������߿w1���SHZ�C�i��9�"����Ǥ�B�c:�c~��Ý���w���0���C��c��G�(���>�FB7���?��?��1{�c���B��,���~�C��C]�Cd�sl���� �&��?����������_����g���v����7�(���0B۵���j�rq���}�c�Zl��w�2�������{�ѫ�
���u�h����i���y,�G�~�����ѱ�{�q�{�.9$���i��t�w����;��j��v{?�'�p�;�� �l6�<'I2�+9|���!;��=�]۹�G?0�W�z�6M��(�^��e...ܦ����� ���>�JzlC�-�x���=��5���?�k�ҽ�Y�����A���l6����+�    IDAT�5�<�j�r�)w���cs�j�ǊE��J���m��8�Ă2"M�{ �yJot���yZ����PQ��9a!9d-HG��|���+�����4,��x2���:,�K�{��߿����������G�����ر��}},��27��篅���/;t�?�,������)]����cfL�sBr,�}����s:u�;�t���g��6�c����x̏�1{��T2��{�<6i�\����7�Fv��e�������5���?��o��7�|�7o��ʲt���8��\ۮu]�|���u�����G�q��������ޤ�p�K��)�ө#'c�u�i:�٩��_a�o�~�'�~�/�|,�����u��^]��ӧO�������1%��T�����d��*���"�������g��y������S75V��+,8T�w����UU5�c��E^7�����cw_��.�����I�N?��#�v�) �y����kO�z�uX�Vh��I�{�T+_�|�#��)�O��54H�Tk�]{�ܲpW)�^�*e����:��yjm�	G��u�w�޹�T�7-�)��(I�?���z��v�$Wck���1y����Os�OS=v�z��z���)���sh@�w�x�<̾k���1Cs�s��\|��>I�p�_����to%T}Nš�1$�X���~���co�&M?�K듦c��􍛱�?��ʲ����r�4l����{C !ӣN%n��֮7��V�/�X}z�M_���H�i���|�Ƭ�7��j�ɡ#6��cס��ƺU��{��1�ӟ\����f���1��!�wS���ln����'M�g:�v����r��i��ߕ�5_��+Zx}��vzm���;r�?��Kȑ������?8]2�1.�U�);�$W*��@���lÿ7�����:!��������3:�k�	�X���d�"���ԁ��=`�>6P�Xcf߉�om9F�ooo�^�'$J̵�j��ټ�V+��t����Q~���s�>c{��%}�/<Ձ�1;�c��c���:\s�{�U�5}��S�|����KO�>e�U �y�>���'cU�>��s��tŏY�c���c����Pp�"�e��v�������?��3���z�vo���WWWȲY�:@��I�}]{���|�E=��3mu�����D;�ڡ��igWm���������>c��{�T��|�1BŘݺ��`�Z�%��tl�R����|]�<G�e� N�1�cR�c�{��PIe1n����i��q��|��ſ��p{L�5F�YH�����J(6����󵢃�X���u8k2�`�X���T�u,�����
V���r�P����T��S��2�׻^_c�0z{��o�}�%� \���\�{���˽�ә�Ӡ��d���I�c~�Ǻ�;,8��|I�9vm<v��R^���9�H>G	nY�7pn<|��W��C<F2OU%�ȳ�B���d᱄��^��>�	�x��ƾ}_��X��� �M�o�O�y�7���Q�%nooQ���1���%a: ������J��y�H��t��T�kD��{��?fd�K���n�X.�G�`z�Y<(���׻(
wܼ�n���?�>�����(���o(�Ѵ%�P�6�C����|��}ߣ(
e��f�ݺ΋�+��Y��cO�9�S&���:H�N��q��7tv����`�OTi�C�ӷ�A$��k ���
9?�G��Ǹi������`������h-���d����p��}�Q�N���,�5�� �����}׻�1)k�����`��
P?	t�,�������CCJ������\�L�P�쾨�}D��Sm?��s8�!�}����6?�����2�p��~�/���g��_�g��7�}��cD�~�)/�S�s��>r��u�{��9�����s-�>G�����1���8h�۶� �S�~;eY�a_a2֍?��V��n"���m����A�pǤ�
�Ǹ�1����'�cZ�}׼:K�?��>��}G�~�;� ғϭ���ع߷Q?�^���[w�w�:e�N����S��/�Q��+��md��8B��E�V�E�sNd�yyl�P�Y%hc�Rc�_�����=��whM��[|m�X��^�,j(/�tc�{�R��v�ޣع翕W�"���/@�М��:�uu��#BQ{	�&��е��K/yJ|��~L��c6`�����}'8��Y�Z���n�6�e�R����>�;����v��g_��ox3A�G)�j8�2ٷO3���$����c��S�k���R��tp�+?�g�v���R��+��]˾�`�~�Ϭ��1�v����ߠ���f�u`J��con�DH���z�v��EQ<���#��e��Ɵ�{E;���}�����8wlpd_��c��ؽ�d�Gۜ給N��"�ڥ�À)���a�!�S�}��^[�	�9�{����W>FV��@E��d2qÂء�/O�t�U�U�j��,~�ef��Xw�9���\Y�Y�\J���>�����s�Lp�!q�u��&;�(?������|ˡ�������c���Lȼ��F̍�����O~��ç���M)���+e����P��\[���:$�xJ��s+��D����2�|�Z��[�C�c��}I4�:��U������l�#�mۢ(
��@m��\N�S߫����f��,]g�'��:�V��>ǷQ�=Z�Ͽ䩄���\ �{����=؁�$1v�iG��s����0����Ѭ�$I��l��|���M���������	�c���=�����/�Fw�4v����������
_:A�H��)� �R����3�䚤s_�/���A�_���SN\���;4��%�����>v�{B{�F�%:��P�!�����>G�˓5ܟ��g�ꫯGQ�� ~���?��V������l=v��]�ύ��7��ղ<�cp�ktjSY~΅}�&�Xz�cǧc>��c�9a�Wqk��7V]��V[\\^8�D������qs�n35��~�e��H��(���~��M�}���~}<�B�9��܁�1�����C�27z_W��<�2,�����A�ux-�u��ׇZO�}�7�+R�}}}���k|��wGuמ�~	r�%_�m�s�-B��I�������$�*��pD�s��]i������n�}���q�E`���ď�����}�j��b��s:�/rul��s��>����� iT4��͛7���D��7������ݿ������/��/\��Ԩ�C����D�)-�cZ��^_���Kk�_jx����n,����޾S�C��;8$"�L�����1��-���9f��<GQn:��!�*3ŋ�ݟ����կ~�o��֑�C��1�S����=�������d.����{��u�~?��'i_.����#�ۭ.�d�E��[����:���=�Ń�v����q�BQ�,�����O�r����-�8FQ�|�[?P&˲��#������!� ]�9b���9�O����C'�_j_9��:��5m��T��S��cy�S��$ ~�F�s_��SZ�=���d���͛�7˲~yy��ŗ&�O!�Oy�}��{��}II���s"�_�M�1���ڡ�˷�C���cy��ZGq#���� ���o�������^�Ѷ�;2���H^�p}}��t��v�rP�Ě�lE�����_��w?����f:���$(����سor��{w�Dd���#�O%�c�Scdv��.�ٮݽ&]����ӧO���߿w�EE(��d���X��^<�ցD�w� �a�o��?���7�������Kvq��^�n�Z��>�����.�A%Ac�~`�o9}=�����I����+���W_}�o�(���ñ��Cݻ1���<vJ�R$��.�ku?OEr�*�8�'<���b����w�<���t.�(ÿ��/��/�w0�������j���<��z�tz|OMvd�񤖓ј�>n�l9.;���q��?�G���j����?�(��v]��yT���꘡���UU��v�<�|�N�m���|���/��/m�_�� �?���+F�~� �.�_��C��4QQe-�^���ꫯ�$��޾}���������|�����o��۪���a����]S|44�䈝;vT��J�"��=q6Mc��"����?~t��D�z��pڰ �cFQ��Oj�۫nw�ok|�i���,�AȄ�\��v�F#£�^��N��>p'i�u6>��×A�$��n��'�� �쟃K$D��S��46��`B_C3h-dx��u����r�(3������\.�u�����f.����#�cM����n�������?� �������y?TF��T�=�L~�u�_����\��l�w����Ǝ��H����cS҆�"�H}M5zU=�)AQ� oQ1��s����\?Y���g�E1~���x���D/v����V�`0�k0���#B�cL�U����UU��z=ȭ���𺈢����d2�M�e��2]Svz���<����$y��T¢׃]��ؠ�*3�N����y��u����Zz�����`0�5^��r��ƥ�N\��X,id����j!WȲ�u��<f/��o������w=�L~3��&�����2�6SG�AB>� uv�ī�fc���޲K�voձŷc�_�e�%5���ŭ�`0�k0��U�1�{R�]���C�˥����u���<%I�`#�M�Do�q2e,����it$�\wv�T�RU�#5�R�MiCUUX�V����+\?������#��l��$�J�2Fp��!���p���8XF�- ����cL�(�;���l^�0���u����Y��vbEQ�i�KRK�)^�`"7�����k�p�{������W�iUU{�;��a��C��Fp��"����nB��Lݸ��iv�H���S�Mn���g��[#�'xü�2�C��8�1�L\�it���X.����q����\A%)w^�(����I� p6q��`�y�zW���Z-j�bM��Iu����%7Fp�W�8UU9���������n�[DQ���Kw���=ʲ�v�EQ��
EQ8]'���Z����!i���m�(�?~Ļw�\�+;�~lk�$H�=v�#9^�ר��3�9]!C�!�dW� �#�t�`���,vHny= ;9�f��v�}��()Lͮ�`0�k0�:��sF���Mݠ��}oIp�� \(���{�4���Q��N!��FpO���u�=Q)+�n�X��X�VN�@�&ד�$EI��P&[��k4M��t:-mxh'���,�ж-6�}��GM1C/e�l6�����l6x�������+�5��Nc#��ـ9j%�8�m�m�T4��DU�)CP�w>�	i ����:�bx�5�:w]7�Xs"�,ˁ��G�ܖe�R�(1i��jױ�l6ݵ��|�)����t:u�)=�䲫��˲lp�P��ug�J7^C���B[#���ܻ�M�}������WR�����LD��z\�i�N;��N����}�'�m6DQ��H~���k��6M�z[��/��(�0�N���j� �N:��w�=̂���]��x�S�b0��� �����-����e���� �ms�$1�p7?�6��S�jGf8M!C�6J
(C`ÂE�&�(P��X��1����6�<xO����MӠnjw
C����l6n����ꤒe.//�u���r�9h��f��`�`xu����ڶu�ڵU3x^���V�7����*�e�:��ӑ[`ש�N���Ǐ!����L����QʢŎ5y��,K�`84�E�j�yoRkK[8���A�͛7�N-��i���t!�%��o�1�\��n&jl�hб��+I;{��y�;��z�v@%@jo�����f������g�����v�։\v{Iv)I�{B����@�$��Y�9��˃r ��>�m[�V+�i�鋆������}�c:�b6�=���y�zk~#��Y@�1A���}�зS;!�,�fh]��!TU�d(\#ڷ�c���3��NvR����R~@�K�5�������s^�:f��['����(=�������1��puu�֚|�|ߠ��:m#��Y��a�� nhL��j�)d$J���i;uH�W?��{Zh�2�N]�u�Q!��@l�<c�N�S�{[U�#���3
X������8v���x2؁�y6�������n���S�MYS���`0�5Ά�C�G�UU�)���}�͉����_F�2�J��v���@�kƵ�E�;����(A`�׎]�(�pqq��$q�"\O ���OJI�'(�����BQ� kA���5SU� �PO��\�ᬈCء���񃞘ڥ��m�T��͗VUu]��1���h��Z�q-)5v�@JH���n1�LQ�ί��N�,˜4!�c,A���[���-N�(B>͝^���\K�ׁF��';����p���#z��idIr)k��G�H�s�4�\>���}�FM�������6m��GrC�kx]��&��O+?�3��|��a@dQה1#��\��I.T�,CY�(�UU=������W����K��]�G�4mS<X����G���0��n��U2K���p"$��찮�kGHy�6M�=����=�T;$������{�k����`�`8��i����qd�U;6$@�,iG�\.��l�&���-4����{$dG��� �%��ш��t��t��/�����4w�Av m�O���U�A�2L�Q�q켬U ��*7��X��:��\���j3�}�$W��5�~��b�\:�(��w�(Xn�F~N[İ���+����,F ��:�L&�i�����p�R��R�Mן�b�YE��
�ۥ���|'S	�I1O NE���$I���yeY>�1#��ـ�9�z[c��>�
��Ǎ���5�;�����3�T1����o*'�/*m�X� �\uh��;�(�$���׻�|��q�g�e;��NvĶm\�i� `�G�ޯtK��:Fp���N�WU h��y�rsӮ�~�nv<�V#yn|���,�z��2P�3���XǨղ,X����=nyNb�}Y�N�׎�t�L��M2��7���6aQ!�# �y3����A������X�~ޏk6Fp����v�E���#%��Аu�s�:�>�YT%�L�Ř�����YG;�:���:��p	�5�)��ǮChAŎ�.+bN��������c�:\H>2�`��m׺��A�^?�df0�5���q�6(x�$�a���)j>V�>8�0z0�s�7�d�4��?:e<w�8�d2q�$X������B��,^�X��ɶ��uiIhy�3�y@^ @0(�蚡*��7��g�ͱN�[n��������}2n�Fp_����+��A�A�u����y�?�:�Cp���Y�(�P�%�M�|�#�bw=0��i��k�u�BE�I��r]|�l��`0�k0�tSb��	-�4�A탘n��Ӑ�\�_a�w�y�p��Y���إd��sdY�5$��nڊi���A��<�I�q����(P�%�<!��8��WZ������m0��g���`x������&�t$I�nF���PF��&�9-�`����q��ԣm�~��P���"�#-�0b���k��#�iQwܭ?���8�$��O-��<X��`0�k0�T�W�厐��\�Ӎ��_*���Q���v�O�Z��U���>������r�~�2���l
x0���)��q�B F��6��D_� g�����vA�+���(�`��&��=��`�`8[�C����I�:���o��ѝL&�n�߽�AhCH�B��δ_�z$������=;��� @۴�K�f۶�L&����UU5��^zϲ���t�˫K$i�<�Ip5�cl����{Y�� ��#�ë����z����f37|��g$+�@Ə�i\�#^�K�˟��V�d�    IDAT�����.4��v8��-D8�F{(%�$�V��K������)=��E:I�X,�ܘ���{琠�_���\UU�K���#��Ym�eYb�^;�[������o�c���n�$	�FQH���|���`��6�WXk�~ڞ�j��-u���EQ�m[�y��|����.
��:G�x`8����1CL&GL	�% 7 �����k��d2A�en`͑ܶ��^����p��"po��&��]�.�b�Q;"�XW���!�ӯ�Fl]��2���C%��A���&)bT/;�M�`�Za�Za�^���N_�P�T9���G�5�����ۆ�ж-�����p ����(hh�&�}��A����T���P�����'�{�k*I^����F�a#aSw���Æ�N��R2D��X��뺁t�k���z�b��[�`���5���)r3K��M���*��d��ٔ+hwO�C�n� �Fk�紅׎���3���|JL|�(������HrԁÆ�N/3�A��0�����Ĉ:j=͡��r���͍2�k����3Fp�׿�d0�BJz��1)��H-I�~���k����y��{���u]��`�N�7�s���- L�Sg�knk{�uf��nQŽu<ou�r_�AB��n�X.���0�%J"�\��,@"˩x&Wm6�u��ۑ%��ɮ�8��vqF�NG|ʲDUU���u�Hj�f�iTa����������v�u��p:�C��5�"����}�ݫ��>>�����J��1c�^�k���23��gEp��?�s��Q[nj�m�"��{ޢ���j2���`��D-��N��}��k�w=��q �-�f�qn	q�i��vr��G]��~�ap�m�d�����^�h�����l6CE.&�Ԡ�����p�&EB��-����m����7A�%�y��u����`��pl6|��q`��)U�r�_<�&!��f�A۶���<0���\^���$���%...\�u�\b��b2� �����=�>��^]]a�Z����r��f38�1Fp������RS��;�t����Z�dN&��Mn��P�X{�i�6\��A�~�Å����ԭ�J�s�4�8q6r\c>w]׮�K�l8�ZSG�X,E����E=r]�����)7Z,x��-��%��%>}���@L�b0�5��f[/ �[K].1�L���p����yjd(7L��s$��"^i���������u֩��:)Y�?��w�sRH��#LZ�@�4�u�e ���1���f @�7��=O'n�Ix'�	����"=���`�`8���N�+!%9�67Q���n���VG���u���򈜖b��������9���@F�iu�0!���]�;��Jn9��D׺�����Ous�2���u��k�c��u�ڶm�m�;�����t� ��9���]�$��V�`0�k0�x<��� �J�廮DyR�@rZ�%V��{M�|>�y��`
��#����)I��1��q�_c�I�UƠ��|�����sB؆N#�� SPw������Vb���=v>�c>������`0�k0�Hx�,�YrxDɮ��y>~��
EQ���,�\GP��t�۷�2�,�%1m��z�Ȋ\��*q�n���=�Π�3���ȭ�13x����xu������d��<�����EQ��k+a0�5Ά�A�,��1ʲDQ����Qu�4N���$K�*����te�i�ק%@UU�y��[��GI.����eaT��*�C=0��X�(m��JY�XQ����~2�82�B�1� ����*�;�2^ �* x�L�s���?c]׫���%�*?o8�e�A[��v;�o�x]���'N�� ���5��&��C;�<�a �}�b�/vIpiȮ�]_+`�/��_����@�)�����̿m[EqS�1������m�$	=Ѕ�P?D��� ��;��Di��'<:w��:�H��0��j�,�K:�˓���^�]׾�:\\\���܇a�:�u]��*�E�����ہ?6�c��#���ݪ�P��K�b��'�9I��{Ef�����m�t��Oz�}8tbG��%��A;��Q�@�	�������wx����j����c�\<W��v[yRO�1���]<ט�؝�4u�sc�;牻�l1�|��6Fp��"A�� p�$�7��H�����z�}�ݢ�V�``G��S�d8�a��O_�0ֽ��Ht�}��!����i�.j��N��L&Η���eY�"�v}z}t]�,������, pZ\���F#��Y[.��ǜz�L��v�h#���ڋ�{4Tb_���2k`P���:O��_x��
t�����C�&p�̊�ӂ��0�I��\��mQ�%�8��Z�h��若�뺁T��[-^�\��,�6`$7q#�278Dr�a �I�:�I��rH�����[���\�Tj��y���b>)�����-�Һ�� Ϯ�y�N�Ӂ}�z��I	�-�&H�z�kDC?���(1~a0���Dpٹ%�� �nd����ˍ�q���s�MؼQO��JP}��1����-��4u���p"ʲt�q�Ӯ5�[�Qk�Ø]:)�]JזD���z(�=̘߱p��`�`xu����$IG��(U������5	/}n��I�.�k$�t���M�U-|����q���P��ӯ1��*(�e�.�q�/�$eQ��n��-����E�~�+^[o����pf�Ig۴�`���d'@������OJ6����NKn}�CBm�"
��]_,$?��>�[+dNKp�ˢ%MS'S��ȅ���5���@�HpY�<vm#��Y�v�C��0���N����u��$H�	1�l �Pi�ڃ�ka���3B���M�>��U���%���G����u�U ���j�ƴc�I-5������|����|���1Fp��$�������d���q�?��Ѽ<2���p������YqM�0\�K�]L�- ��T)J����f���DQ�����q��ӑ\ BJ�4��`��/z��C�I��:�����\����\������'�~��]W��;�����O;E�lǙ���'1&�d֡$W���u�|�4��F���j�c��:M�������r�:����� ��l6sZ\�p�N�enx��1$�6Ph0�5Ζ��XZ����(�!r�J4��wHP}���'� \�����T�@�����ɭrp�pz�t���r��z=��}�������y�d�~�i��\��U���t=C��#�Ѯ��h������(XW�Uح��b$�"�� �W�%����u�v��r�t��a:9�IQ^�hE��X��ɑHdIp��ﻵ��f��6�����p���7Ci�x�����T�����G�Fv^uS�,KdY�HkE��n�v p�O$�����5M��,�Z���l�t��X��%�Zt�şZ�����1�iڍQ���k|Pbl0��g���6-���-��G�$�L&����� u]����FNCz��A����p��J�]/Z��Z��Z�v��{q���i�N�Ȳ̅7���ʘ8@ȟk�(�\��,16���W׵����z�R0~�~����ӂ]��d2�X��?��Ns�U�0���}=�{LZ 	+�<�1�L\�6lC�Ҷ� �&vs��k0�5Ζت�?m�x4�^�̪W��\�$I�t�f#��ćE?h���7h�2�o�����<���`����\`g�Fg n؏�I�Y�a2���HZ�m�?�Q7[k����p�$W��H��4hj�O �)Ǣ{9�_ŀNO~���k�n8�_�&�4q�C�:�$@�%���F�>������u[�E6����&Y��:v�ּwI�5�A]�\��l.7)�P�7��T�Ŀ�ޏ�Q]����c���ӑ۪��u���aQ=�-�4�C��U�ٶ-ڦ�6NGp�D��	eY���S�b-|X��e���ןQ��k0��gEnuS����pD�$�c|G�M���u~�!Ү����]w-J8h�G�c�l%8��$I��4�}��E�����n�(�­���i@z8K1_G�0��\o��Fp��-6E���G���R�W׵;��R]�X�V��s2�`6���*�n�u���i�XM�󵶼���[~�����b����t������j0Ƶ)�ґW]� ��']��:��\���R�*�j��\�M&�����,����[���ׁ��~ǖ���Ѯ<��vQ�^�#kj�9h�?����Q�1-����d2q��:f�.z<�iq��%�Fp��&@����!n�<�� q�cM>��C<����k;mC<��r�� �������Ñ`��!�`��9�,sr#��/P}r�'.L�w1�4��O8SR��g��l0�5Κ����<����D<�n�M{?L���� \�����3OG~Hl���<�m�z��GG�tvC���(.�S��;  �8B�]�/	.���}����H	�Z �6���c�>q�yFp#���[�������G*�R�	`��i�b2�`�X8���������;�aW��.eY:}%�aY��q�c4���ЧϮz�ν���N&dY��G㳵{;*9���U^���1Fp�����m�a>sIE=�bw��^���`��`�Z��k$I���k\]]9�C�!Ra��P���/}���t:]s^�c�_�]<^KFp_���{X�9'IB�Q�׺�ѵڮ}0���?��5�k0�5Η�F1�(�P�I�;=nUU�,��+��r�ٝ���q��g�'cc'@��?~t�8v\UG�Z N����z �j;�Tg��tPُj�YT�k��Q�RI���<щ����Q�1A��`�`8�Kr�ǏMӠ�V��Y�����eY"C��U���r�l��)����m���\v��<`�5����ƅ7x�A��o��\��^�N�v�{M;���f0Xj��u]�ہ�^�BH��^6��gMt�'	N�u�{].5|��t@xf����k4M��t�$I��3�����z�v��م�$%,D��qk�#q�p^J|Hx�8JX�y�{�S���VwʪD����7�L&�B���:(k���~δ��\�������a��{�����u��;'5��Y�a�X`��8�D�����ǎ�/j����k�מ��8�8WF��#y:�b��b:�Z��+��~h��h��ӫ�i�q��l�<��e��kȢ�W���#��Ya@p��v�8}��=��%nnnж������I��r�&�N/C�9�O���טҒ�m���['�Y_~@�����vj}�c%���Y�!:,�۶�u��(��ݩӂ:��[�~�X5��gInIp��A��u��8�WU�w�ޡ(
��sG��$AQ�*��{g,��H��M��o�Q< ��v�'A����B��K�$���up�$qׂ�t��v[U7K�J�2.�2��'�U�4M]qJ�
I��#��Y����iPV��/�	f�����R��I�>y��*����Z%�+J...0�����O��wz�jw��v��<Xh��TGV����&I��|��l梖I��{��{�Q��e�j0��gG��$A��(��I*Y�6CJxĽ�lP��`h�UU�NOUU�n�n8�)~×'�///]�t:EUU���?�������x�x=�|���ؙ%�M�]Բvܻ�C�`�������j��6Fp��"?��S���E��l��t��b�;IZi�5�N�e��8^&�y�9�!2�,�4�b�p��� x����~��6�^�ʵ�)�S-R�H�<AS�(!R�[�Hc'��:m1����s�$	b�W�'�7��@��HX%�:�n�� IGp�(
E�H�&��U����׌�%%���/-V������0��]�b�}�Cg��7�k0�5�~'��У�^ n����4�L�Sca�	rh�*�n8H~ �,KG���BY��fSZJiȃ_�h�&i�}�{�Em�ڶ�z�v
Oj�!B�T��vcjC��C������p��(�U��v����	���۶m�Ϋ�+�i���Gx'|��6�R&)iU���N��ch��u�_I� �2w���/D�N��� @��#@ � �:���r����p�#J~�߲������ 	b�N\�}��|����
���C�p:r�`� 0�L�ڰcW������֪��GvI��__vQ��v�k%�cP� w][o�y0��:��\��,�G�:m�.�*��i!�g�s(m�ٸ�̲WWW শ�����u�JZ�$u�w �����j�5A�������e	.�C�� ��F��c1�~�>��{i�G�6��`0�5�<j$)%�Uͥ\���͏6`�0˲$g���v��!�څ��]�=XO���5sT���zN{OshP��x���uW9 �]�l�,CY����W��\���AoK����P��T�(@���'Ŕ& pDV��UUa�^;2l8-H8��,@H���J�tZ~�<��򚱣�ӯ�~0]���<m��b���:H�ϩ5�a"�c׽U���`�`xuPn��6�8{,���#l=U��W�B�U�u�^*#ᚰ#_��[�(�G1��qŉZ�EQ�I:��`��բ�ި��pZPW��'�������3�S�᭪
UU!�2,�m��(�&)ڦuג�`0�k0�:�3�S������Ū.������� �}�4��/�X�����5��Z;�|��Q!�7� Ax��[I�q�^���# �`��,C�e�[�����-��4ui�}�#ID�لFp�3���?Fl �B7���7Fv�tj?�2G��ú{/7T���b�٠,KG`I� `[����t�I6A���-t�����چW"�Q�x���P���}��j=PK8�ܶu6��g���0�OB��Ȱ������v�)��p���AuU0s��.�h�m�:r�u�>����gY�4M�����R��[o�ݩ�� ���������Z��꺮qss�4���ܢ�#�Ù�L^̦�b�_��Hj>��t8)�"w<M� ��gxy��I��>�����f\'�a���ka�����]94����ڰHa���,���:X|�0�_}��f�AQ�l6���Z1Fp���/�N���˩�{@Z5݌^�enՍ�����In�4(�����!ɍ�عZ��Y�<T��@���`�=��	n�$���uvw�y��j�5�{�z�;�og0��gC~xL�dV]HZ�$^�K����EQ����"`/��\Cj��4�G���8q]�1m&p����׈f[�ӯ3��΢�'�9A>�A@]+?�NՒ$��&�`0�k0�ݦ�oP�Ī�R�P�(��:Da�Wf� ��cP��NK~�	A;��j�E<�V�D-'�~/�>�H��t�)	׬�{TU5��RS��u�;V�Pw��n��:�2�th�[����p�WӍtB�^�L2�L&;0G^�7�1)#<�����i�)w:�1��(��.7��� !�-��� �Os�y	 l�OKp}		���S��Jz�놅PUU��֮G���im0�5�{���6cWӍ��0�WC����%�a�k;GP�F�箣���f�l@��\w{{���[�@�'����{�Ɉ�9X����7yw]�$N���a![��#�J�۶E�wh;�(Fp��6In��²;Kg�����40�G�6�ɏ��\��b��-�qc:�:�??�:I���)����/Va��vu��s� ȲlP�6u�A�۝/rQ����|p*�1�����p�$�ƆS�x�\D���08���&%>A2�sz4M3�w����X�L&����$K�:�;�$�ג�t��O�_��`�6L&�y��򤆃gY.���Y�9r��m�#�ù��8�11j�]    IDAT�L� ��u]���.�w$'MSL&Gn���}PcMZvi��p�C������vR��n=;~vL����:4F��ͭk��	ڙ�u�\.�^�1��������xT�k0���JhuS#����1�_�&��>�L�����wZr�u)���������޽s�J�O|g��$I�S�,���DU�#�kӿ�X᠙ʐؽ�)����[���������׮�o���\���.I�X�@��f<�ֈVv��OW��Cr�,�b�@��������ߣ,K\\\���z`��'�y�펦��94��Z��:P=4��_ױ�B�mVoc����{��`0�k0���I��)UO�G�m��Mw�����i�6Q�_Qa�X`6�!
��/q�4��
�7�6�˧>�,j4<@�-[�m�w$�i���X��k��V�\g��e���9��������С�`0�k0�%ܴu�=Ӎ��Q��z4u3�d����G���ӭ�%��͛7����q4L��*;�~�����}�b�k�[��hlߓZ�O#�Y��i��|��m����#����@��
�O>R�ӦmQ�$��x�g����+�q�u�������fx���Nc�
9�PN��N<Wr審���)P]��w�����~�v��wE.	.m���O|�~6��gn�c�T����I�u@Im���:^#��_��UUa2���۷���F�u(7��߷F��9(��+�r����;B�����/�N�1�UU�"l�#��y�vuƢ?9p�MT	-������'_���:�V�,�J솎��S�Z|�E�_��m���\���d��:�n��ZY���z00�����1ݭ��}߻p+V#�Ù��]��nV����yr�ȗ2p
[?�1�������r�&�ɠ Q�/��D�������P���i�]����u�����<V�{���\���I�ߩ����몽�%
�t��H��{����a��b�Z!�s7ae$O��F}��CpI4��b���R=���qy��/�~�j=f0��gM+S���ͼ���)���� �� �\.~�F�N��<n�\��=5�I�����^'A�"��{RE�\׵u�^i�ٝO�Թ���}��*z�j�	3�����n�.�?ǒ�#��ق����h��$��ծ�?U�͓�)Jl�ܞ����tU�@b�{#��Zs�(B�e.���lxy��i�q�,���=�(��$I�,�W�'�^/$�|_��7���|�;����p����j�A�ug���]W�O3#�a���Q������8ƾK��:�4V̨c��8�]ҙa88<Ȑz����"^�b�9X�u��ۻf~��15����`0�k0��aǆ�7�n���%�xv�h�A�� �{{�5��+��0��\_}���} ���IW������>�:�>�L&��M� �2$I�.x?����A�k���+�r��u~Y��ć.����pV�'e	��g֗(��Im��-J��a���NW����?�|>x�v�T����u֠3˲)6�<T��9...�u>|�� PU�����m`7,�v��۪��i�V+�u��iJ�h����`�`8;�[�%ڶt�)�����!�����7d#��#�c��J�8���[����m[�e�'�.µm[dY��Ҭ�{h!:�L���,���u_Y�l6,�Kl�[7��X`�N ���DQ䴹,Z��v�y[Fp�3� �����6Q⤤�d�ฒ2��#L#��b���N��Q@�����\G�]=��#�`8HZ��$�ė�4;���EQ��ǏH��)Q�5��i�:����]���`0�k0�%��?�������t�];���U_\#�'�}�# w��:7,�G�at,ݶ-�n��u���9�4E�e�#o���������}����']/�
����drc���`�`8{��wm٩Ub���cl�FQ��y�����D�`Џ][�������T�S����}� CɃ ���v�a��ڑXޓ����:�2dY�4M��sW`d3�G�=E\��Y!c0�5�c�N����Ѹ]��K��9�V��h�Jt�Dt��εw�j�\�Z+�����É6�8v:h�zh���������M�`��kG��~�a�`0�k0�%���σ�]�6��Izv�$��k�m�|n#����:�⬠���	���n���e�,�L�r:p����a����^꘰o���$ƚv�j��`�`8�P�f5���c��9pB�]%J�������3��Z��Z���O���<�|$���+�(
��k�ij)W'&�i���^?���{L&��:�~�u���b����N�}Gn�&�`0�k0���7=%1wa�&��t}�����g��N_.��Zgݓ� �0xP�h1�q�*=џg����ﶲ��z��j`��i��D�]��]�V�n�������`�`8;r�M��:�|R���&;=��|>}�M՟Zpp����Ԇ��Wv]�0���F��z}�a"�2�������L]ר���	����UO^X���˥;���$I܇�`0�k0��������sq��Ϊ���s脛&7��t:��������bPZB�$u��wk�M� B�#��P��D�G��;�Nquu�������UU�X_��2,*����aO-X�}e@�!��ߝ�ܑg:�����y[��`0�k0���n���#<꟩ݸ�(\����\I��X� �d�Wxü3����^��pmH��~�EA�-�y�01�����TU��!�$�Q�F,�7�cL�S�y��mZ�M=�gf�c��3Fp��"��Ѵ���KI0�����	�����l%��1���� MSW�L�S pN�ĺ���.y.����	v}h����$
�+V����ZԐ�FQ��l�<�1�L�!�آn�m�\$�t�U�m0��g�)�Onb:��K*���u=��i�z���U���k�Do�w���ԥY-�K|���I����F���$=M�`�^��kk�G���VU��,��l�m�t:�l6s�yJ�f�����#W�	�Xud���{��`0�k0���6���έ�츙jg�����Ъ�\Ɉ�묱ڷ�i��t꺫4����k�?�(B���T��f�u�0m��.
mۢ,wE%��t����δ��?5�,ti9���p����9����pć����P�N̫�Ώ�Ux�q�[�n8-Hxnnn��l��]X\=�V�)>������}���I}�i^��$�\vi���n��)g����x��IXX�hܳ��\��,�4*ٶ�u��97�F�K"Cr[���FQ��b��,Q���^�������������۷o�e٨�`н�z�� p�vR���i�|WU�m8�%Y�P�a:���eIi���{<�%EQ�(������a�dI����pVx0	�l�ڮE�~�sʣi=�l�f��ϭ�kl�[$I��b��l6��4�{Z��w�u�(Ig����@0���r!�L^/���/���S�p�"F�����z�v�~��Ȯ�k��}�oF@������FQd���\��<A�$�J�4(��u�[��1�
�3�)>g]׃)}%[ܐ�!>}�#MS|��Wx����,sI]ר��� k'����U=o?�����k����n��t�~�Z��� ����v�����庳ȡ�m[��5�k0�5Ί�jZQY�X�V���]���#MLeO&��q5%z�i]��\(o߾ś7o�e�#E$'��s��a�#�����H�0�e�?�Π�����V�Z�x?gY��b��ݽ����  ���ynŪ�`�`8/h��A����4E��H��gS�G"��*���4EQ��>�����e	.���I6谻x޻�]x-@�"{�(�%]�@��n(��QK9���Y�C:�ǂ�	�����E��ѣ������ S��b��v�Ő��\���{���S׵#��۶EQ(��>������!���\gG�-=4��^�ͺA����P#���8��4�>���0�Q���n����Aʏx3�W]���d2AE����s�-mۢk��dIYʚT�d0����
r�9�DrJ���HpI\i(?�L������.2��zD��_>�$��n�g���G��:jJ�%��.����Zҏ�ē]y-<�~�I�F���� M8�I��`0�k0��m�]�t{��p��V`
�6Q��
��Y�!�s\\\`:���|��ܗ
:�m; ��RE�'~^�^����>Vo��'��pa�5�い@�-�Ujp٭��vm�$�{5����#��ّ?�^I�Jf����.�K��ɲEQ�0y�E����V����@�����d28�Vh�nw� ]O|x-���@Oz�E�^���u`aJIA�$�� (�O���fqD�K�Bh��`0�k0���1�����2��sãQ~pӣo.%$����=�:�X!�Q"�kA)C�&��Q��n�م%	z�:���2���ʵ�ƚ�:;�u]#˲��]=��z�Rbm0��g�(���c$4�$�}��r	 �q ���.u�c�$d3���r���92��H�(a�{�B��"���߯����:���U���_�M]�(�½�@ Il�$�:a��/a�"�`0�5�u]w:(�M��z�N&�u��f��v��f�8�1��1�L\w�'9�����^쨳�{������]:vY����{�fv:��N�����1VH0I�y��8X��}��Fp����?��ۛ������A�H�t@t4�H�$9L�X,�c�FY����RNZӀގ2O�0]���{q�]��#��e�}O���W}��kxy�K�tY���q��.˲X��-`����u}���:�f3׽�l6�k�vcFp#����y�y���Y�!Ig
���h��^�N�������w0���#�1��r�Dɪ��a����!�� ���AyAY����#�8�b�p:ZZ�i��b��y�� �!�c���=6����f�q�+`#��Y�믿��������,��	;� ^�a"
�/`�Oq}}�:�<�d��l6t}�ˁ4�'��UPNB�B�e�� pG�~qҡX�	,���1�#�,*)9 ���^eH$��_��/��%��z��:E���[��k�XǓ�0��熐$D�{a����ww�	��Q~���t:��������=-���Tͩx\#Y���ZRb��i��)!��}�i�5�L&��f�-n����M2c�/Oc����z�ƧO�P��0Q5Fp�W;y��dW���j�ݎ��y>��/��u{t"���No��v�y�{�����_}���R=Z�^3MSL�S����eJ�%&:��"Iɰ�d��0�|>w$�m[�V+E����eaC�<�g�O�=�(
��k׽uÅw�8`��`�`8+��Z�\�=��t�HɊv�8�E��� Q�D�C~L��ܗ����c�x^v��dLs�?I�x=В�?Kg8�� ���uUy/��ܸ{UC\�F����sL����j�r_W9�1�\��Q��;��a!=�$�!�吚���VT !�^]���'?���������*��B&דn
\sZ@��I�_�P� ����5t��L&dY6p�����n�PJ�(Q����۪�\�zm�0Fp�� 7�4M]�QUUH�\�̨˥|��k,�Kw�Q�$Br�	��eEQHbҶ�@N �i�˲t�.<�� �����ϧ��FpO�1���`w뎮뜟-R�eE��S�Z��^�k�����:��\��6�$I0�N�v��̨6��8��M3�!�n�N�����#M����u�T<		�HnHj�����<�h���k��ć�N��?X@��kE�ֵ�k׭'���`�;�������u�}=�`0��gnP�|g�F��JpI�����˪�P��;�vvc�p`��Z5����q��l� PU�3짴Dc]u��Ib\׵��c,3e�,����4�n���,�eY��p`��8�0�^��{�/�ݿeYb�Z�j���:Fp���?|�Qz\�1ڦE�6@��`j�3�4 ��5��n�f����3�׃v�$�l6x+�s,����d2�b�@En@�Rv��UW��k�m��lv�I��x��j1l0��gGn�C�vtW !R�jr�5n�$8� N&��)l���W�Л��i�y���\�7�z�#j)\�,�\d3?ϣo�(���i�8�ő�O�e��t�B=4����(�N-~Ǹ��ra~3u�����p�$���"e��vm��c����f���8��4����(ɲ���uV����M�0D���]Z ����dY�4MQ���~� �Ӂ]t���N�������>:C�]��܊V��+Il�$������l6��/��H��`�`8kr�$W��6u�<�d��������n؅	h�2����A}%��,p-��u��E'���E�_�	;�>=����uWٱ����f�����t��gqp/A�72I.�4��A���i�#����pVP+'%�$���S�^۶�(T]8|D�.��@{)��
��FQ��v��(PU�#�<���o�[�Q�.�.S�		��N�K����v�y��u�,߲,�b�pC�c��oH׎.�O�-����\��l��؆��Ծ�1��ir9P ���sw}� ���i��ז���%(��r��m[t}����e���=������߈�i�_vfYhrM�,$ّ�����s졚|~�9�XЃ�`�`8gp��:�v�:4~�N��9���)��)���ޥE�,;��~�{D��j5=P�f�$ߥ@?��4AB#ȡ4�@��AKЅ����~ޏ;���t�q�`V����ώmkm[fEQ Bt}gėWٺ���f#�s��'!�3fy�U�!� \x{R�n�<�����h:\?�(lS�r_q�����!��IHp�~x���e���=���hoADp�f@��x]^k��ӵݫC����d$1���k�������ׅ�.�o�}������u�g��x��cE�a���	�>}��xD�u����w�}���Bt��=�;�ab�'����^g�!��G]�F~A����y>OU���$���{>���9i+�@�m��:���g��e��A  �䰛���\R�zo�۶mQU������0;�$�����Y��||�/?�S/"��pS���C��:��[E�?{���F��r���ڄ�~q>wh۶5��'(,Z�z���Cf��&��Op��C]���J+��}�������^*�� �
VA���'.	�����H�k.u�����I�~��'l�(��繭I���q��:CDa�xV��6���Ľ/t����g?v��zg��-�f�����Zk}AWn�0�g?L��wj�I�'�^���<8��AW��#�t������ۀQ��2`�$=�4�3 l���0DQ�V,X�$���pi���,^��h�.�wW��� ��
�M�� ��%֕��ݽ����A�K�"���$$��2��I!��%��'��쭻��v�omE(�EQ��m[+@�!.�ϔ���{��.���4	� �+7����Q$Bi��;�$�LNZ��g{�h���� �uN���ZZC����y�DR�.f��%	�- �	���<��WY���v�����t�\��@��מ��w����F�� ��
�͓  Fr9$��Qy��JZ�7}�8�Lm�}��ז�����X�����,ˬK��|�����5I�죶[g\#�5+�,�)׈����b��+�5���
�� �4�e�������3�B���l!4�8*� S���Mn{�%l��,@�Uv���� �u?p���<�h�f�}�U}�^��`|N�K��ⲙZ�I)��K��`�w���C�k}�H� ��
�M��u��}�g��3��q�h���"?����2�����4M�c=ȩz1+%�    IDAT��}��k��@�e�o�4V\z�? �;�|6�45���t�bh��S�!"��p�䖇��&�[��R�駪=�]����K$W��uݵ�֖.$�^�9M�@�Z�E�Ε�8~�u�w�4���ja��}�����[�=�_����kK8A�Ć��	��;�I� ���j$8Y��p8� ��a��H��`W>�cBbd����uԫ���d�5QҺo�o���Ï?����Bv�}G�[6M����񈪪��~��焄��Ԉ�
��\��@~^�
�EA,d
^WɃ �<GQ������քZ��v�Q����A��k�¦���6�����??��Vk�=~���w��o��7�>}���bdG�N'�mk{ ��3�.	mY�(�Y�a�;��D>~�u#"��p�`��d������b�=	����ϐ,����"��>	_>u��$�c�G����f�̏a�O������u��p�}�}���HF�@_b]vp���t��(�Һ���\s����p^� �� ���4���~�I��e���$�+l~�i�}��~�� _2������$IP%��ٳ�?wd۶]t�|H�8$)�b,���@Ǩ�j�}a;�0�5����w�Y�������aP�5�qD�����i��AW�O0}��:�u��mS� � �Q�(�r��Yc� ,}V�/�j���ܹ�}��#x���@� lm�0��׺��q%Pw�v8�Ea]yvxY��㈢(����+׻f��˵�r%�� �+7O��@?3��k���5���"^wzk*�<\�/V��9\�/�(xoT��4�4N���y���`�_خX�V`]��L��:���_�!���}���?�r����� �� �	�S�[G}%����&��iI$K���Vf�s��_m����0�%������֤(�2�Y������s��}��&Q^'g�
n;$I�dz�¥����j�>��Y�P%���kEal������ADp��H�a��ѫ�:�d�kt�<��/�{��xR�I�m���L/^�"�Ғ�x��4Mֱ��4.���<�Ij�뭨��8~���wA��C�\�K����=�N<����=��@��f)���:�� �+7�(� 0=����UU�i��q��i�e�pM�ǥCVw����#I�3)���w�kHb�`����8`�W���x|��~��߾���s~H�Ã$��d3>^v Qa��ő�ep8��d� �+7?	�+?dR�5���a"���mQU��#��=������oU�`�	���{"�"g�LL�>��Y��u�Z�y~~� �l���!t��^v����v[?���p�@iE���4�m��x<.H��(� �+7�����VQ�M�a|������q:�ć�㥄+aP^�e0�8,\���ZS'm�x���/$�q#�b��Z�P	W$�Ahvmk�0�G������w{9�Ɓ4��AWn�ؒx��^q��S�x�� �n	$>$B���}�O�¿0��uq��ksT������U���3�5e'0�"�QhO����cr�� \��z�bOn9l��;� ��R��u�
z\A�x����\_=z?M�Ea��nI15�<#�$W�n�In���2�v$1�ȲlAd�������Sk�-���?������Ǐ_��ѷ�d�Z��p������Pʑ�`�$H� �+7�y��y�'O�� ��&gR��J�˃�it]g�?���u��u���-�(B������V��8w�1�_��٭�]Ox�7�8��뽏���4M��2J
��1�?�����ж-PUڶ]�2\A�I���=�����#�%�%�	�ap&���b �;�$B�W>�ۮ�n��Ce/�4M_�1���p����r�z������Ou]�@�06��}̵fW����R�5>��O�>��k/�� �$.uR/�Z�[�iF?��ʁ$�!����Wؖ�=i�����k2����� 0�0~����
��eӺ����G<<<`�g���㫯�Z׵�u�h�ֆ��u][z!�-� ��
�M����E�0:r��fו��<�h�֮��׭��^��מ�v�]ֵt��ʺ����uu�iB�	S��ql�
�zwi0M�\�ϟ?���=y��L��mݰY�u&?�#�~��amGI��A�����T��N���*v���7��9���}�Pѭ�#<\O���4Mh�A�,����[ݻ&�$?i�^L,�zo���i���-b��d��$�~�Em�&cI�䕌%�AWn����hS�a����	�<��� rX��H��z�)?�"ҳ=��I��P�0���(BF�������D�s `1U�����o�n��o�~�w�����/q8�4��O|a���>�(�3�}�����m����z�� ��
���Gx>==���	o޼����iB]�FX���@F���L��������	������g���;���1�8FFl���4/��Ql��$Q�/d�8�~����=���kK\���c�ynE��z'S��~�d&"��pSכ���2ILӄ���x�:cF����z��/�c��u(K8�mGr��To���,Z������kO˩$I��	h��0�t:a��m���^��<Ͽc,�~�GE����qDUU�@W��X/i �eqKڊ���WJ �&LDp�v��MY�������~��u��B��y��A���<�8�B�+b{r��׾�$:6x4�Kk1�e�+��M}������@�<|�2��\�a�Ͳ,QڶE۶�3�����UU� ����K�""��p3𱜻��"]�qD�vg�sw��F��ɮ�I`�,@0�=q=���K��kM&���޳p	� x�)�z`ƌ(~�|����bN򄫯������;� ,���q00�EKF?���$�މa��&	}�g&�Qa���͛7(��|��<-�S=�a��:�δ��8,�@^qi�^�rX��u���-n7�"�Ѳ8���:��֡ŷ�~�����=>�����6�wG���ѥg�n
$��s��(�eY"MSu��g�:���sV���¨��?��O(���?{'}2�ru=0��r����!ʲ��:�~�b��ˤ�~��wg-�����!r{��r�<�]���u}�"#�y2�=�Km���v���CY����Ӭ�UDp�6I�?���u�$����z�K�%�|4��5�����l�a�����ijGMӘ'.��Ip�i�п8n�S�|��H�����8�Q���mq:��4����v���R�I��p���i��$� �+7/Q�����'�N'�]/���rp�_���_m���ս���g�JH^|Z�_3ߍ^b���$R����_�u�88��<P[K���Dadjo�������h2� �+7Kpy}IO�al�$BL�t1���i�E�S�kr+}�d�k���b��y���]{OX/IJ|r����5Z�m��]3��1�Q��z�_���0x����@z||���#��X��A�����5Mc�@<ԦiB��g�Ȳ�<	��D~B��ۗbzE~�_kvh}T/�/%\��+~���zg���8�q8LG������������u�XF�=%�SA�q�����\AWnk��Î]���SuZ�y��TU�0qwwg�*����z2�c�m��$�4�����^Y}=�s��$y���(`�����un�$����;�#��#���n�[�_vy�4E��V���\co7���mH��c� ��
�M��i�E�N�N�����
�]�y�Q����(Ǳi��M�d��	�.��-�忻z���i�.�s��3q��%	��R���Kؖ�ך�zk��u߯���x�/�}o74�1x�ADp�.	K�e���H�z��S�^�p8 ����-j�q�����H�/�¶����O��%/�g+�5���H��묵_S�VƵ��۔u�Y�u�Έ��}|�� "��p�!5���p]�P�[׵��n�$I0�#���iP�%��������Oz���w�0����:s$@$�`�E����������5^?M��/V������39�0�=�i�U� ��
���M��x<��vo�&�i�[�!�,3��-��94�"`~M�Dv��%�6\��� ��W��v۶E۶F�.�KIi�6��h?��N,5����m��,_?���A!���}�<���V�,"��pk���!�sUU�isHH��&����Kx�E���� }�[����Z�g;P��I�s�0`�F�2��_q�/�>��mk]��u�3e$��u���(C�MM۶f��&Q������)_��A���������<m�<�.-�4>��*p4+�rA��6t��'lOp}7/�"��{������Yn�MӼ����^�sM8(棲�?Y��"�:z�;��P�! �;��3ADp�ȭw7����[��|&6�>�ŕ'�4y�Z��{�������v�K���F��_�/�Q�"/���Ķm�v��J��p|��,��ܳ,l�$5?k�4���g�s���ܞ%
�� �,�e����n��N= ���쿼ǭ/�۶��S� �s��wm��$�^���+����ϝ�(^t�8����T�\���ah{��� l�鉛g����*|��Y���oFݽ=K0��"�Y\A�*�M	.����Ұ�7���i#^��=:E~�E����ڤ$0� �{�$�+'������f����/~�|T/ +V�a MӠ��E�����҇�3AWn�����49�m�8Z�r����wm��>&��n�\�JI(-����-mÞ���(ƌ�ܭ�ƅ��ڙ��\mKp����������R�q_������!�0@*�PDp�E�a�J3�cS�J����C%6��|ty��y~vRx&W�R�Dr��7��1�^{K4�0=���e�l�2~��K�j�m����pm�[ʹA�um��1��<��k��h��^��+� ��
�M��y���mt/��̭��I� �##�M�A���eY"�cBѹ��يN���1N��@�y:wo A���i^F�H]"�|&��ہ{x��g�6�2+N�yFUU�� �6��*���r� ��
��n��I���	/ �xq^`��䖃(��TV�m3~���'�FR��y\v����~����'��ہvo����� 0
o_�嗷��Ѵ�L1���å|nA����'��d�Cg<���?>�[O���.m�8�O2T��8y��>$�/��,4֤��1Jy�q�I��Fj�f�]�*K���#u��CQ�N>Ё�ʼ]��;m�`?��)����t��^�j�AWn��p �l>����u'=�8y����RڃEa������%�]:vp�e��� 7I�ynd�iw,�X�0�Ç_I�X��}���/I�/\ٝ�~Ք��a��E�5ADp��OEȲla�σ�[���<��5|���%�|�َ-��ӡxEr�׋��{{"�m��8Y�#�i�i��4�)��>_s�m���===YǞd�����3�$ɢ���eY"I���e���vb� ��
�͐���k��5��C���v$�>��vD2��HpH`IRر�]�(�EH�&H����qD۶ֽe��g�vc$[~pM���������N4��* sP ��鴰�E����(�� ��]X��p[�0
1�������x��پ�_�E���]�1�,{����8���^t�L��u]���'?�Y�p8��
�!��{�0 �c�v;��{��r���(��p�>���ub�؊�
�� ��Y[FQ��k�K���<!BdF��#�m�|ԫ�������z]�����1���_voi-E�1>3qq����۵eY���;A`�7v�o,f։w��^*�A���:�$�����ђ�]�0�����A����,8DƎ^۶�(�S��a�8���0a�2�0�@I�iv��g�]ba�=��ѺQ!�s��{{Hl)U΃jeYZЃ���
)ADp�&�m��^�$�����q�0���OO�H�����⁨x�/���um>ǞА�a�qM_�.��(�A3� ����g�/X���$MSE��,�BX��}od�,˅E��5�]'�	� �+7Ap}.�%oK~��k��:?����k~f���A,lCr�q4��4��F�E����ĕ䕃cy�/���t.z��S�Z,w����&�2 �=q���ZA��m���w� "��p����ú�����������5G�g�[8���mۅ����Yu�ؙ[&$����}�B�Âǻc��+�_�o��ָ�(7M꺶�:$pm������Ss�"��A���$?��%��׽���5��ꮻ�+R�+��u.Ij��}�����"v��,؀Q���k-.��"u��Cr�m
�t۶�2�<%��d*�MN�45'?x*�� ������kw�g�G�����=��vS�+N�z$�k�d+v�<Q���<-R��z��X�EѥWa;x�F�}��/T���,X��1��/��ZDp��t<�x�	.�v��p��';�$��0n��Nӄ�m�eق�A� ���<�B�Ex��u�Z�	n�L#[ܾ�_��B���p��[� g-/�؂ ��
��������,zz4��)V�.�}VEp�Gd����Z�ҰТ#����8��<�����������ym�$1�o�$��'�'�C�.V�|��<�AW��8(�q%qM�t����qy�M��N�u�!��[�gv�|g�"�#@����Y~ xE��m�}��$Y����dB�p�G�z������g�L�@\A�	"kds�u|֞�뎮O�
� C?�
�t�k�.-a{���G��]0��1�a�JF{I��5��~^kp�N�k��yMd/����縷��\A��kH�8MM�}o]=Z���h�i�ځIK!چ�$����:d��(���<<���a8=<L��.���	���z��}=8�u�k����gHb��'��r\A���#�������n
 ����x��D�����^&��y��-�����{�a�g$�R�M��/��=�����Ô�`��|�_3F�%�m�M���Rڰ^oADp�f�����u]����Ai���/@��]a�N���E��$	��kab{��K���M�sm|ZU�u������8	.�mךE�勞��q����@����O�y����<Ϩ��~��^� �0A���"�����(��Z��,C�evx���������[$lO~�o�輸/�g���C�|�x�u��B���4��_^vpɪ��)EQ`��#���՛N�04�K������ ��
���Kd�]�4�u����W����zݾ�Q��"�{l
ےܟ�ў_��Zo�E/D�O鳸ag~�۽JM��&#z�\� �2�e���� ���}o�.���Q��DADp�f���Q�ǁ�u/4��
������6Mc���a�5�:�k�C �i\���}b
���Q�0��k�yn��>"V2�m�y�1��B�Kb;���^��(^�]��\C�^��c�u3#"��ps��g�Sn@��	��|H�@��f�< Ip��&�	��j\�����
Hr����|j�'LL1�뮿/d����Z��ֶ��-���]סm[{>���796��, �!�A����?}�ֻ%�ӌ(^Nͳ��F2�kR���]��`���!?�֒��0�KѬ$�\���Q���n]׽�t
���uxW�����O�}��~@۶������nQ� �+7�� �������D�$߽��خE�iB�4��m��&��S�#Z=����Hp�(�0h��8�i�WCI��Fē\�Gم�qc������P�?��g�  IDAT���n����R$ADp����<m��ut�$���������(����kL]kn���+K�&�$Bk-�2@H���z)y���5���N*����U�d7�"$i�8�E�}JG0UU�,��͍ "��ps���ƘBƃ�z$@�ݒ�t]g�>z�fY��^JI�,m�Y:����Ү��T��Q�K�DI�JR|D�t��3\K?@Fi����������=C�y����
����\AWn�{�A�eg#x�xQ��i�[���a@UUxzz�n��p��x^up�	H۶V�������a"���ŌOǚ�	q#��Rup������zǔ ���Ӗ�ť(���{��W������0�E�� ��
�M�ݞ�m��C��a�8���L��8��kA��,Q�%�$�Il��&��#� ,͊���֖a�uGpY�P����u��qD��H�t* lOpIn��I.;�� �8]��s��|���iBQV�p_��L\A�)Pb0ϳ[���3α��l�I�. ��n�����n����ڮ�rYOjI���\vj���O�Ǳ�h}�p8>�cp�o���Ǝn���q��kL�?,���;\A�Y��x���'Q�z>?h�!�,�~����y�,���t���<��VpI� K3+P�v����.�=|3��;(�@�t���¶{��Pv�	�/x�0<� 0c���^�Р�<a��͂ ��
�́]Yjk9,DBK�C��Q%I��܈�<���q���Z� lGr�hǱ���r=Hh|�=MR �L��(B���͘p�u��$�����g��0���E�]�YJX��bH�YDp�Do-G�u~���<�Q_��w��q����Q�UUi�k��L/==[zM3b���/|�wMp�A$\�R��������KK��}��E��eH�\A�Y�c҃0X\-������W��7�k:�'���G��=�d< �x^�y:8��:b���PI�`��#�"�GTUeq¶�)tI� �2�P�!�g�$g2;����?��!����>��΂ �+�Hp�g�u�;:`����/I�����(����*<@ؖ�R�����/:���fqß�R~�4�xPg͟�������4��X�����'���Fad:�<��uN���A۵F�9H PЃ ��
��e����W���Ah]����[���,�F��0\J6�|��� t=�yD���Ȩ_�u*��  ]��3�G��m�x���\�,J����0\���q�N�q&�I�X�����-���-`�F\A���"�����Id<������/�yu]�a'8�2���K$����'�������A}���z��:��b �u���4;v������>j;x�.~�'�<eI\'	�a�<��ݝ�Y�!�2A��mM����@Dp�����$�>����z�ƅ�������`ƌi��V��)��xe ��8�8�N8�N����(]}���P�v Am��
�8��`y[��z��8���9�iB���,�poσ���"X\A�}B�мG�϶_��/2� 3�c~2[w�B�][_���n�@<N�>}�����1v���#?`���m	��d�f�k�N�[�z�0~=Nb�ٟ�������
]�u)sAWn��x=?���@$2�j�:�ud�e���W�R��$
ے���M:BY �4����k;{&�(BY�8H�d���DIE���9��mK��~�5F��r@�[�y����䪪L��u֒��� ��x��zǃi��gS�!Rk�ˮ����~a9����יkA�����"3�u�R��v;��{��p���V��mיds�&�]0���%Ё71,n���FƧڭ;�k?�� �$(`G�Q�$D!�>B7wF�In�$AY�6}��mF�H�*�튘$I�Ղ�X��1���,��6RQ��(l���*\�`��0�u��$�sA�����q-����4YraEd�$X.
� �+7	V�4�R�9�ϟ��%��wyp�<��fYf]C?���϶ćޥ����:��k��ዞ��Q��"q�~�&TU���P�5�4Րٕ.	)	�������4�b/���u�,r���ɎDpAWn�`�Y���%��j�9�h_�|�"ȭ������'	��]C�6�~뢃^� Ѭ^��b�߯��B��fnOp}(�/��_�u&%*�ra+F�e',T�iBQ6t�N@AWn�����7��Ł�5��z���~�����)��:ćD�w�=A��$$�mۢ�:�mk_�������*.B�G]a�}� � �͸���f�gtm���z��4M��(1
���H"�� �+7��u�.m�|\�����+?�}��m����@���d��!@��P�µ�a���� �s#Km��x<�x<���5��Q�4��AE���뺸�n}��0�gM=�4�0D۶�B��B�����-��KYԩ\A�I�ˎ�~�?�q�u�i�NΥC��3��"qh�D����Є~q��:vQ���k49Aρ1��z��{�N'|���:y��ｐ}W_؆�z����<�@�W�mA Nb��������<v�� "��ps�$���$2u]/���]��������5	�a;p}�k��ջ[��+���p0�T3���U~�_؞���Ļ(��K��Z3��y�~`��x<�����ĳ,G?���A�����	�������u4�%��$��DQ��m]�<4E~�+b�>���퉭'5�k�4M���di���'t}����c�jJ��zs϶m�8�m��$Av۽a������� ଽ�A!� ��
�M�Z��O^W�!���MgɎ;�|=�r��g'���mי�m��5Mc�y����ZLO�|�?IdY�,�p<��W�u]�x<.�
¶��� ͻ.*�ש��;o]���ы��V�.�B�� ��
�m�W��rP��{;�8,����� �����L������շ��ے��:Zz��<ϑ��B�����^�BB���F!��2y����:oOp��	��Y��ah�	u�Y�پg��,�3�R ��ӓE�Nӄq��ZDp��@r��y/!XH�39ʲ]�!�2�:e�w���S���p�u���n��7K3[���_���ya�?���z�����g�I,(�0�.�Z�ri���Y A�����v0C�,"��p;XO@�����MK'��i�Z��׿�.	.�5����=���j)�0�"f�ij���e}�� !�l��9��{�+���-b�qD�4V�xG�^rD��5��4M&U�s\׵��AWn����������Vv��%	MӠm[{��Z�$��Dt�]cvai�5��{��?5I��?�+9�rdy�y�q<_�w�/v[����ӓ�-o^�<_~v]g$�)u^W�4��#��:{#g9�i6���﬘AWn��D���G���M�3f���v;3�����7�2�yn||D��� �����Hp����s(���_����p�Yi�"/r��gǗ����'���s���y��e!�e��,����=���d���(���"2� �+�Gp��.��w�ؐ��yn�F���X��u|�r(�����e��ng�fh��t�2���S��$	v��M�@�4&7���<e$i�{rJ�2O�9�/��:G�$0���,(��Y���E����4E�ux||��tB]צ�堚o~� �+7��o�~���~�>��w�c�$��S FL�8>w��iv>@9t���B�0M���~�GQ��H�;\�p7 �>���`�����֤�*4M����Ey_\�7}��(�E��a�.˲wEQ �s���a�߿��`k�g�p8X�GUUFn)C!��1� �+����8�S��ڙE>���<���գ��?;�#���.0��8Ư~�+�i�!��Z�/�����0Q�(��p@��W~&y�|��y)Q��AC6y{9a|��7����}���|1S�%�<�<Ϧ�eW�Ä�*0����M����!M�va�0���5� �+7v[ٱa�W�$IY�Y�`�#�NCJ�t1�Dr���[��߿���?h�,�4���4�IX�p=�,�������GUU��;��)A`��"a�e�N'�;��%%,F(G!�A��[���1��c����WA��� F>}�����V@σHY����ޮ�۶�A%�"��=8���^�q�Dܦ�y?��w�<���
 L�Y׵vf�}��t���x©:-�E�6�y��mϲL2�-�g4�7�L�O��a@UUV��T� �-	/�]��H�+"��ps��;Gi��y��	.;�Y����V)W��ha���A|��X����������>�w$9�\�}o]]~P���{�GTU��}e��,K��0k��i�j�7���}���{Xv��\�9�򒵗�&��%MS�y�|A���A�|�$�;�v�-�Hvi'Ť3 ��cG�Cg��v]���$	��=�iz��7�H���C�4�"6�������'$G��x�(�a��z6�3�4E۶���+��7�R�IY�6�i{x���a��U��O�@���M�{ww'�?A���ï����O���p8��a�|�� 7����^�3f#EUU���a.:D�Mm��n�������v�wMӘ\�< ���&��8FQ��a3j���d���n�u�������8~���;��W5�� ��i�Y���P �1�S�!���+�^�E�D�� ����<����/~�s:��vx����i�e�nGTU�O�>�ӧOxxx��xD�4�����-����o߾�0����,m��[E��TU��k1��60�������n�� ��z�B�&@�������� v]���M^B�lY�fH��E��+^�����}���&H�?�@�?� ��7���(��4�t< `�	� �J�ǿ�s�(B�4fO��l����~�p���k�(�L�y:�k�#����q�$�������g�du��������{�ei򠪪��{��.�a��AQ_�Z�o�#B{6�<�4M���_J�""t:
��]5���8�?��{�ah��
HR�q4�L �|P��$�qD]�F�˲����Ȳ�}Q޼y�01�ioIl��f'6L�dZ݇�#����E��Dh�&��ZOӄ��'<>>�m[$I�7o����q�m�ƊoH=.}p�0@�w�}8p/GA����۷o?�a��(
��}zzBUU���H,���z�(
�
��v�գ�����qdrև�,E|6�o~������7olPȬ��EQ`��a��c��c�۝������?��?>�x���p�,��a�N���/�B]�+�׿�� �)��ޢx��t�h���֌W�:]j���1����CQ�ς�s4��O ??�<O���C���P�-����zv�h�C�IM����Y�a�g9(\�;�:s]����n��p�k}zz��tZ\c���R��k�7o������zWD۶�8�Ȳo޼���~����
q�x<Z۶g�u�e43e(,h��C_���1M��gݯ "��p{Ȳ�o�8~���{xx0��Z[�S�J��l=��G�B�)\������t:}���h����C���=lM��u�9d<w�)51��ldY����	�DI�+�"<==�������g�s˲�,�|#���gqDi˳ۊnUAWnf�|-��8\t:���v�۱#�8��o��6I������G$I�������o~�u}6��������ݏ���hߟ�OOO8g����4]48�D"���e�uy9Pxww�$I4ttE�˿�˻�������*��|��?����?���eY�o�A�刣�ЛɧR�4M��#N���8��
� �+�J���i���4�%]�m{�����-�h)Ef̋n.I2���	�����g��� m��?�����<�1>����G$I���{�hRG�u���������	|�O�ˮ^Q��]�$�;�Z�u������'�����?��a���,=[��8����f��s��T��;À��'<==Yq�����-"��p�xxx�ǣ��SV@��y�k����|#$qb\��(kxxx����e٨�mq8�$I�N�9v��*�N'L�d�MӠ�*��v���� z��9���s|]�a��Y�}�������T�����r����MO͸^&v]���Mc���ۉ	� �+7��,�i���W_ٵ4���q4�BO\��8��+�5��М�9̲L�܍qww��$I��n���(z�upww��o�� m���d8��� �8���\�����~�����7o����4��(��=<<p����	��#�i2ّ����C�,j���8�Z�� �.v��o�yF�4#M�IV��7)E�_��H���<ϱ��h4�y�[��o�����; ���������iFj-����%����b<ofG�8�=�y�]6" Z�+���> ������m���$IF���45�I�u���H0��%��`e�aEQ�ZkA��� F(Ñ7�    IEND�B`�PK
     w�O\Z���N� N� /   images/7e39c2f4-a1af-49ff-bc26-783004b83469.png�PNG

   IHDR  �  �   ��U   	pHYs    ��~�  eXIfII*          �      �         (                  �       �       �   1    �   2    �   i�    �                    GIMP 2.10.38 2024:05:18 22:57:08   �    0210�      �    0100�       �    �  �    �      �M]�  viTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 4.4.0-Exiv2">
 <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
  <rdf:Description rdf:about=""
    xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/"
    xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#"
    xmlns:GIMP="http://www.gimp.org/xmp/"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
    xmlns:xmp="http://ns.adobe.com/xap/1.0/"
   xmpMM:DocumentID="gimp:docid:gimp:af2322b1-529a-4b8a-bb63-8a16a68440cf"
   xmpMM:InstanceID="xmp.iid:e2ccc7bd-7563-4995-8bdd-ee54e5669374"
   xmpMM:OriginalDocumentID="xmp.did:abf57cb8-2880-4205-bc1e-6b7909543b7e"
   GIMP:API="2.0"
   GIMP:Platform="Windows"
   GIMP:TimeStamp="1716065832663280"
   GIMP:Version="2.10.38"
   dc:Format="image/png"
   tiff:Orientation="1"
   xmp:CreatorTool="GIMP 2.10"
   xmp:MetadataDate="2024:05:18T22:57:08+02:00"
   xmp:ModifyDate="2024:05:18T22:57:08+02:00">
   <xmpMM:History>
    <rdf:Seq>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:1c838011-541d-4cc5-97cc-1bb3eecb47b0"
      stEvt:softwareAgent="Gimp 2.10 (Windows)"
      stEvt:when="2024-05-18T22:57:12"/>
    </rdf:Seq>
   </xmpMM:History>
  </rdf:Description>
 </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>B#3A  ��IDATx��k�-Ǖ%�#2ϫ��%)��=�i��mذ�?]�0����	����a`c��xښ�Zj�!�o��33±��;2/[�0S$c_V�y�#2K�b��k�ҪU�V��z�����xz|8���t�qe�Q���{�(��������?|�����jժU�V����V�Z�z���e�����Ɨ/_��>��q�r���t�4&ܜ�t1J_ n��<x�����~�w��Ӌ��E�/>��?�I��Z�j��H5�۪U+�o��GϞ=��n�}���) W�ۭ���jO2`[���^V˕��(1D9�l����r�\^^__I�~��o>�g�g���jժU�V����V������_�~���_~��7�׏�<�Zn�o���F�=�����d�Y���Y��!�E�'��/g9@�u���W����_��������Acs[��*�*���t:�����_Ä��r?v��������g�Z�b5�۪����<���������G_���9/ v�Z�W��� ��������X.�/�k�`;�b�A`��,	҅ps��������ܜm N���������q��?կ�k����pz����b/j]� � ��������/�E[5hժU��Z}�k���t��{Y������Ņ�z�J�no����o���܋T��6�g��� ����L^_�,`ϥG����t���`}����������x}}�^�x�L� ry��.N����@� .�/��|���������_�e��Z��W��Z}O�����x��Chm7g��G����t14�7���V�[9�Z�Z�ߒA�sY��;/ 9tB�[ ��v��������i�Z�7ꗿ����ۏ��c�h]����R�@��r^&L�d�]��r�����P�A�ܟwww�i��\.W~�ŗ?1���?h�V���� n�V��z����˗/?.����͍�����������@
v���a8�a��z-o��� � ��_@ܛ7I*�s�8`���W���me�9�,�������~��u��Xhl,����x�{��\� ������^���ÇeQ����l� ۺS�,$4�F��]��]����o~��ٟ7�B�V߷j �U��a���? \Pg;�Q;��/_�g��N�={�&3 �/��\��7l.���j�&��ec��$
pḰ?��8��t�{�����Q�X��X��կ0������!��y�hb����`O�rO���˽x{w+�$,�=W����.ʽ��q�>{�L���k)��Qy�_���}���_�{�U��Q5�۪���^�xq����n{'� ����y'��V�no	n�ڢ�ү�2��/�Pv-���^n!��W5�s�E/èA )�s����O>�ͯ>��?k ��Z_~����W�?.@�ѓ'O(�pŊثׯ���#��Z�{	2��~��\<���z;:~nMVW8�:O�~��~����z�я~��O^�x�������s�Z}O��V��g������Ͽx���s�0{N������\��{.��)�j�"�����	@ 4`״/`�����.���+�6.$����`w�7��w�I?�G�|r�쫏���8�����_}����G���w�^��½�u{w'w7w�LA��;�d �Ϟ>#�����s����ϐ� �|�����~����'��?����^��j�=�p[���g����v��d{w����'L$�
��ƱT����pUX-t�7��-?sO �>�F
|�@���
J6�!�,�}���|�������٣����O~�럝�]���{�B��P_?��r��~��~����>�[�8&Y��ܖ��x8�ļ���6<�",rW�:���x�B��%��e�^�=Г�\_Sv�7g.�#%6���]��<Z���T��Z}O��맗�W�_]_=z���GY��,WK6�y�U^I�R��$^ 4�f��ǴB�l�\$��0�/��+�I��z��������p{��׿�??]�m�6��fXp��$"�h#��8�r `� nԦ.�.@:P����* �e?2�$��$~��"���L����Fu�ȳƦyq\��4N�}\�7?����"3B���G]�O���f�<yp���W�A���S��r�a,0>1�r���Q�/#l8�tM�����5h=�(A �1cC$��{޳�z�~Lƞ=&o�������=��;�@�V���� n�Vߓ:�?=��^�~I�"�  z E�+ .,"� 4�}�2�9'T ��Ҥ�U�,�ϙ��9`2w�������u>�<{pqٕ}���z��P��0$�4u�E]j�?pO��l�T�-��A�*b��	l�g�.�>�cߗcI~>⌳�n��1���s?ץs��"�>�`����o��T3 ;w��s�qm�*�$���_��Ӳ͈mwe�#�e�!*�n��*�ݢ�ӝ:T���?c�F�^_�z����F����2�
r�, t�K��v���I��S��%�����X��8d[��@d�� ����{f����ʄ�ls�X�۪�w��m��{P����?�}�����+9���y�B��<�m`rA��IHX�L(������S�:��s�J��E� d`��>�� �����|rQWd�HVK}ĸ��a%uw�%��#��Uy,PꁖxW���E��
�x^p�BJ��������Eeq��q�Wuq�P͕��&x1�e�c"� s�mH�xOܢ6�	l��L@z���K��G6���C�K��m�c��ׂ`z��FP0�����կ�|�Z�#�ʯm��{�
|6Y���g���Еc�t���{x���������տk����e���V�7N���8c�=�!t귌�a���=��p�����Z�$#�`��B@���l�����:I�V���� n�V��z�ů����d{{�h���M)g�5m��$vD����T�a'X|���@}t���g3g�%����@����Zʑ �ݕm��8�p Dp�o.�8���=X�m��v���<�w�~[�.�����) Lqw �#��J`�����`�&7�X
�
�^e���9b��?��	|��,�>��L*{�l0�I}�+�k�6�.} �e���;�Y�q����L�:ql�N0���Œ`R�y0IAj�Z���r��$[ۭ*K�}��x,����%'KHO��W����i���o�n�8������i��{�Bvϟ���t�"`�q;9�h~l���[]����B�{M2�Y�����9
���>����������/����ت�w��m��;X����t<>��\��^�||w}�������Fe�� ^�.��G� @�H�Dp{:�S F, R++�J����Mg`@'Y )����L����^��� M� .��FVRTǋ���N��P��#���m��/��]p7p�w(�8�|����t|1 �k^Us�hS�q'R��A&A���7+Zz��Z�-���f9L2���	D�`BK�t�O�)�¿xPv��,f�â�h�T^'�Y�A5�Q?_� ��T�Л��q��$�����{m�g�.0��z_b��н�y��-���=�k��5+��K���}�Y������u\�� .#y���.��_� �Ӡ�6&x�:�.�����ӧO7}����O�_>����k �U��h5�۪�w���}�Nǟ�z���q���y�Z^<{*�^�����nn	>N���H3u��re����E ���I���\�`�加�P@���H�K��Jb�HAs<���� �Ӡ ��.�S,��`���N^�Chؕ\�_�كs��cP)��-�,������B_��ž �qj��sN��}��5�m$�r�F���`��yR���|<�ZN�Y��4!�et�@�s*?�A�-v�'|c�q.0��`<Ǳ#����H������G�8�1���A�����j�!Q�c�����ńcq�{4���ZB��Dd�\$�k&��轼Y�	���Bʀ}O��� ����~+���v�c�t�{v�~�x?&^���v{�����G|��'7��}���r[��.V��Z}���_��e���_�<}���������� ���M�7�ljr��\ l���r>���ٚ� f}�27����U�� db�a�o���.�A	���4�5C��K�O0��/x�v������_U���@��Z@ϛ
���U5�#�[9���r�?�;D	D^y��`�`,K�y�?z�U��K�S���ʌ�U�˷�N�VW��3ҏ�n���P�g08�gq=$!ek,���<�����ztaiA_��+q���c�Fs�:]��-�,0bXo����-������ߚ�b�Ư5�f*�8�|�ϸ��xR����q���fS&$� ���U9�c�k>7�c8��n�$h�Iʂ��\���<x����� �b\�ƞ�:����z�
�ܢ2��&�c���,�r�w�[���O���<z���'7/����6��V��k� n�V��z�������鳯��p��^^�z!ׯ���� �\�86NK�n}��VW���c	�50Y�G ]p�Y�c�s���:���ܾ�څaIk���� ���C����bC�uf�,m>�yC5��yb���������yڏ��^��d_���0��w�zȐ
�,Z�<�&�~��5�c�au_��/^�W���Vu2 tױczU���XǙg߭�\�9���S�,�&Θ8D�xNu�C�	F��~m�2K�R�"�ڣ�n�|�*�2޿��q9��n�}��2	:�z]&DWr��
 =ҳ8��XAn&�\, �U"��.�����^��z���=�M�:�}�1=�σ����:�e�ry����=�2����' �|�h�a)��f>K�7p���_H ������dww+_��KY��>:۬�7n�V��j �U�oY����\�^_`���nn.���y�՗rs�B��^"B�P@��G0y lᲀ8�xF��1�y�r�=v�.�d�4 �BLe'� �kT�/�wf��K�D��D�7[g|p) ��c��Eesq��6X
Ĭ�FӋBWFq��p,��Zn�����!Y��م���'���M��l����\\�k��-�!w��З ?@&z٬ֶ�L@6���o՚R�lbf�T��k,�>y�p8�1G��8>�� q��s��R�]�@���. X�590{���틗�/_4��Y�^�L�xJK�jg��g�Ndzm���\�3�r�l7,�L����C���,I-��U��-�%^CTo_��SF�~{_=X��q��A�݁ �"��RfJ�ߍ݉za �Ճ�������X �� ~���|��?��&Uh��;T�j�-�ן~y{u���O��������_��els�
�X��-+0^X�7�&��})����ɴ��G�XEe/ŀ�A �Ղ�� ���Pv
pu����B��ZL�ԓU ��N�L������jU�L��GE_Y>����AV��Z��݂ɽ�� �ۋj7�~��x�YlΨ`�t�r=����2���A��H�Mpq�L.�pg	=���bg@ښ�$Wӆ��5p��^��.����0��yc����b�B0{0�N�r����4�a��r��d��J�/_���K9��(3�j�L\E;f6��\�������	�+�c�'C	�)�0�k	M�t��u�C�d��r?Ag;��.�;ڟAf&�t>T
~��,���-�m܇�QΡφ5Y�����_�������g����~���m��;R�j�-�����뫏_>��ɗ_ʫ'O�p}���0��*_�ʞfk��~7�wpť��zXa�|��db�MH 
0����`����H ��T�	btd*�S����^zp8v��N��'�8(&�g�Za������.�kz:��\�c��2��<�Ͱ���2jx{����ɦ ^�=�7k��f6Щ�j�f�N�Â#$����
��\�Pճ�:O�����H` ��&Z���n�7�7����Ε�=p-9�e��9)t	0��i���h+��|������8 d�<�`xu-W/_����ܾ��c��q�}��;�'�qb��L���=�%�_,(_��$*e�R��@�_�h��	�v���L{���������n�F6���J��~4�5����l p�|Q�r<�>�_��������Ń��|��?[�����w[�Y�V��j �U�{^/?������'/�<y����N�_<�E!?�8�e��X�r)QI�VL7�+(�GȢ�É�j��qy�aH� p�%^��h)ՉG���v0}�LzRsT �8$}��;6*)��̼��!t�^��	����F���*� ��,huE��������v��?�;l�b�9���l#Kh;�'��r�~�r���s6����wa��MI��Th�ν�K8>з6�\l&�x!��Mo����j�U���M�	�ĩu���2��L�]���=arb��&"'�p�@ ���>q[ ��+~P�� �-�%y�%g�t+�C�D�<����m��Oو��IE�i�����H�8g���\�)M�5���}��(�댙=����Y��`��BNL�x�8;�x �o���zs&0�qCC���kz+���������n�������G������m��[\�ju����������W�=���崽���B.
[ay ��D
�bX�a�U�^7���c�L�:��|�j�>���	��.��+����&��і��W�B�d�'m*�����ЫW��F�Ԅ��j�V� ��-޿^-e��	n �V��D����/\���U�q<Ȱ;�u��u�P
��\�r*���m�^˦�� ��.+ p�l���2ڷ6�A�<���Uӫ6j�q��
<�`Z��ֳ2a��pL*o ȭ���k`�N0�Po�<ؑ�`�o9�������f�Q^�����D�VS��F3w&���+sk,�/�u� $M������\:�X�<�̾��+kn��{�����Dk~�T{m�ߑ>��3&ɂ)�4s24Ѯ�ϱ �q�c����������6 ����x�h��|�����Y���O~�g��m��[X�ju�+��t���X������Mg��hO�Iɘby��V 1hJhR՚ �OP�կV\V?�}�G8���9�X҆���	�#�¨3��4����2B�*�;.�@�y�T��
h�X������WY���-��0�� �� י����Fdm��1Yl�P��A�}s��.5��l�s�Md{`kWb#�;�r���*,��' ���dJ�����;���#�	K��0�2�Mvb���1mT����&�
[Hv7�r���]ߒ�SP;O�F��q9��Y�[0�Q}��5�f6����]4�Uo�l~A�v�6k`Hv �h�����+��I6��u��+���;D��*�=�)�|'�@(>�H٤��L�s�!��=�~�z���;������L�����ۗ�p�|�����}����hln�V߲j �U�{\qǮ�Aޔ��]�,#}ح��i�e�����B�����)��������=��򙘗� �菴c�|y�l��.� K�j� �!s� �@��y��ӥN�=�k|���BoҤ��X�_����M䉺V��Kh��<e,�K`��R��  ��k������n[�O���y��'�	�N���]�����N��/�����w��^<�̂�k2�3ծ���X�Wt�����C�n���p��|uT�ެ��L7��xc-�ɼaqm��w:��� �ׯ���y}%�8p\� �޼��[xT�t�d:�5޻��]kj�)�����t:	�L�T tN*��;���[����Yei{c���������
��#XN�ɵ�vH]8�{,����I�E#��/��������ѕ{��Y�/���_�ճ/��~�h��|�w���������?�qcs[���T��Z��n w	��3�EԨYF�B� ���MzI�F0�!V@K֯�X��%�?6��G�/	���e�S��u�g�3��q�:Z���e=Nl`(�t
�6��~b|o��m�\�]� H��f)kX�-��\Ɣ)M�X�H� |��9���*4+��y��K�[����'�d�3 ,*� ���v���d����zm���v�h�ruW0=l5,�l����c\F�m[�Z\
z'���i XcRv0*��p�K���HЖl����X�sY��,-ko��ʶ#�xt�&	�'�V`H���h�*�t�&:؀�[���%T~_��0
<�"��`�r�L�f5�B������LR�������{R��yAj�$_>z4�8��z�Ž�_Kw� {6�G	�q'wۗ���J��������t8��Ջ�������m��[P�ju�kD��pb��;o�{?π�vѩ��e�K�X�z����\x�Bb��L�K�]e׫5��sR�F�S���� 8G��ǘ;Ջ��2E��؞�]
j՘`��EC�\.g{S���:'[����� 6�a���ae ��r$Ц@�	�o">�VW�bi�
�r�6f���'��m�����֛Àm�l���b�u�_1��/y�"�
L,�Y@&����8�}d��饹mcD;�|EzW9�}��iw�x���R̂�͙.�jb�JRp�=���p9A*�=ҙ��p�a���	Q\`���ń�����4�\�ֆ	�I��H'�dNJ!��Ǳ�+�x`u����H�� O��	�7&>��cfJa2��x)b��JB����}����<{򕜝?x�X�>�z��o�z���juϫ�V��qa ���r
�Ԥ�^
�2� k��_��A�>��Ĝ�Z]��銟��3ڒtO�vVH� �ر)�<�?(��H�^F�t���ʌ2�
 ��I%	5���إiS` i�e�J��%V4��3\�Q�j�� :��w�wU� �Pʹv���֠��4����vlWcm{�*�6�u=`2�����)[;�0�3��Rs�Ҵ�h�[�����fㄳٿ���ԤZ��]���&�@jX^@�ԩ��+��x�A�"A>�0�$�����p���qPF5�l�d�11Y�KZu�-�UF� .�(:l�� UHQ�w�Q(��O ��t������N&Y�kAP˄>M��X%LҬ��
i��`�!���c�6�����s�D��0r� �2�_</��Z6g��EK>k��[P�ju��3���(�/��t�dk�!�0�) Ƹ��g�p�u�gP�^���頰 ����`Mh<��MfF|�+�u�.a��`A��;c�u;x/ 
 �d�W��e3�Yj9��&U)N6b��sk���04��K�0��r&:�T)�6�)㪢[����3��k�m�]����[v�k'.��aX�XIH% �XiC��؄_/����/,�	;{8�Ťf��:әBg�����j�F ���q�m����P���7F�c5ͳZ�3=͵�&W������y˳����۔\������-e��~`,2&�I�uw�5�[�L��I{�؀�:^�\���d�˰Ã���#:�b��G�෯�S�LL܋�NbǓ�
 ~��%���H6���'���CL">�z�������ju���V��q%5V%�)P�,^N�P��ܠ���!�XX~e����Mٛ���G�>�6@��[�e��C|?��"�8ܝ�S�@sԻG�L�lNfu��1Be6  L�[Xs�q���2p��X_;b?���V����kK)v������ͦ͠n��Ѳ�$��t���B���� ����d�x����:�;�n8�\�����5 ���:X5at.�NY�Zo�^��0!o������ɧ�3����������z��OW����b��ll������`J���5�{��͚��'��<����o6D�Vk^{	�N� #��:[h���X̪�'��Lhp�I2����t���{iA<��E�Y��I��*���������UV�b���o��w������������4�U�{]�ju�K�^d�}����VH��:��Qn�IZ)Y�N�vx�/����P���to�i��eV/�h�]�w.u9 ��[�.��6�!��h�Oc���0�GS�HR�H��kvQ`��m0׈��STӅ��n\%����H�[I� v�(Ѐk��LޔdK�!��`$͋W]]2�$�Lst����}	�=r�6��8v=����ZZ�;h#��tVX���R�c����һ�2�x��-\$
����$�,u(�4[��՗gz:d�C��+%M��=�m��2�t�N(���^��H����?�����m��� �� 7�s�4��$���wv=�(�I�4\�1�N�8k?�c2��2�br��"X���(�r>f��?�~�o^TS���,��\�|�kq�V�Z��j �U�{Z���.ׯ�����&MX���>��4@������ۊ�g>����eX.ӂ�����٨�U�v���|t	�`v:*��᩷�3���,{��CR�*ðL���u�����ӳ�MT ��נ��@�B�%Z^�3����,A�T�91�B���!6�B4�L���N�qnS�8&�yL�(�_���e�}�Ke�G��/S�m^�u�b�K��2�x0�-.	(;h��d�1w ��d�'�G������<��V`��緧N�"�Oh�:����,�nW�+k��8�d	�Be�sЊ�D۵� sd ��ۭ�3`���x��U����Cp�������`Moz~\�H���l2v��C�	�Hwz?�
���I'S�j:Ħ{
��4�Lf!b+"�wYY|�&����w�}�����߮�j���Z��j �U�{Z)�ǡ�.	�����6Yy� V��Z��0ɮr�1�p��
b�:�%�N�[�r�I�y
֔fD�5���1&uH ����� �X`��V�G#̨u����'�2P� �,�B��ǃ&:)��xE����:jjA��AAi�t� ���F����at���op����D��'�g�����q�34byߏ��hZ�r� {����ZC���;�s�]� �Ԛ�\۪x,�A�܁񽰂��3�tS�eG�Ebz�FN� �Өzܓ���ڔ�f����dn	fV��;�!���^'50��$��_���Y�8�۝�:q�ݮrm�;��Y��z����'>	�[W���Yu��z��V7�L�J��Y�5qz�f���nw�7�f��~}�d
�Z��j �U�{Z叹�� X`�S6@��Eo+�.�͔�>q sF`�[�YoF�� p�"�X������.�5 �F��%���koP �Vp,8u�@��'���b1�����+9g2ӱr��ُ1N6������ő@�A�^�т  2G6����e���ޅ��5�w��ɮKx�f��!��F9n�e=�X�8���B�� �`�V��X-���9GA1�.�!��b��Rޡ�=�ޚ�	�~C��!��(X�/�����MwiD�o���~uVmv;����s�U�}5��G;��ՆB��:�	z\�]�&8 �۲O����r%}�!�ǲ�햀�h����\�h�Z��6˝�d�5߽�B�������MXLO�Q��&D�n��9ǽ�~���WWe"�l2�V��q5�۪�}-���8�����ҭG�ڲj���:)`$����*�+��?�a���C��~�쓩=R7I���\�0v�̎�"�\]2�cY�V&R��%é2�di%����Fc�	,��K]:;�du	Em�2�ݘ�^�Ơ"q�4`�ĸ[6.����3��X�h�nɖh6Ћ�br�9;[��ű�9Oޔ78�Q��h"iو��t�R8��E�� �	��;���T�I�H��f����mb(ϡ��3�,�K%�z�`U�n���r������Kˋ�$����'�zR� �E�`Jl����L9�jŀ�{}G0��Yc|k��݇ ې��������L�0��x�v��>�,����xmA_a���zz ������t�B�����&}���X�N��$���r�����ͳ'��?j,n�V���m��V�I�[E�h�7��V: �3��,�.�w��F]���J�Ygm:�S�&���֠�"P��9���,�'b�t��6N�_]�+h�����)G��v�K��ؙ�-�N8��y��C��NJ,���Tِ����S����f:1��}��Åc�-U���M�iO�56㑓����cv��X�T��\�%�<��E�����d
���M[�1��E�km�K__�47ڋ�$�C�3����y��6��/��h�`���c�{��	��q�&���2$�лFS]�`����w�m6K_���<?D����[Y�f��	��T�e�Gg�2�J�,�ܡ��xRo�q8j�F��U�ɅG8�ECǪ�V+�n�����$��=\�A?���v.O�c�)�juO��V��ii��F�*�˧)I�D�n�	��_S�L_�Q�Sڃ�V��rem�lo�aǻ�����E����uV 
I�lTiB?(��6;��F�Xٵ)]ʜ�yN��0?@4fg���4@n��@o�U�fr�d�ή��@elʊ��eMJX��X2�6�נz=����Y,W�+�|�݌v��Ǹ\u���o�2��2�&�,����fCy�1�a����߰�i_C��h��`j���f�v�a�&��������v_���NH��ͪ6;��F4�w4�{��	\��X�}�T�L�<�ʰ�u�P����q��w���;$��Vd���2����Y��?�>5H�%&~%s֠��hc�a���x8�ҪU�{Y�juO�]��Q[-eQ]
�u�P/�D SS������:$(��¶'c]�8gw�n���H6l)��2��icø��v?�S�殙��,m_��]�͙ͪځi�2k���V��-����I�v�{ȃ�,D�R5���_=�lI<��#�1���@�-���� ������ ��l�޷oc���}ØAO��gR��q�Ā��U?�|<-�8��n� ��ȡL$����F��v�VԴ�r�$�ټ_�C\>������,0e+����ŃQ�8�rm �
Ѓԣ뗒�N���W|ܟd�Ћ�+`�� ҐE$M1�[�c�/0�e[4���z�p����s<�疷%� l��L��,�ON&�ֈ]�����˟���s j�v��)2D*�j��~V��Z�ӊk�g%]��n�[�ۅ`j*�0*��/A�m-�@��� �o�`6�i��:� �/��	���3e���`if~e
��Ic�d�e\&&�kM@]��'�A�j'�44��}�2�4��42��0N �<L����6�����i��c�䰄 �V1�b�5�%�TP��%�r�Իu`�����ɼ;�<z\/�V*{ �IĪ ��ٙ6�%ӫJ0����<��(��z-�d��Q�d�e��Q�NYǦ�$l�;�(y-��X���Ƕ��%�c�>���5y�"��G���� l0��H�c����}^��vr�P�2��0F2ϙ��Mr6+�X'�YŹ�6X#�4O�uBܱ#x�������7i�uR�k}<5�۪�}�p[����U(��b��q`�A���\��7@�5���ݐs�W�0��w}�����n�jZ�%�A�Bj�=�N��ݾ%nC�N	љ5o�
�<5��\T����Ic2�ȴ�	���r�TST�(��;�%�9y��o�7���6UG�"� ���:�z��_;��\���P��Z�Џ�� �|h�evh ��.���L��5�� i�6�ԖȠӽ�W[���Ƃ8�ܬ���\���y�<�[�2Du��<���\n��2���� �����n��nz��[wP��@W8*�6]0C<�_Q�l��c@	"tOp�А
l�O��C\����e�����	aZE���3��M�����@*R�A�V�Z��j �U�{Z!dj�%�c�zX±h�u�&S�Cq�2�΅�X��nՐ�7_�-��|��U�61@D��o+dB���,�f�o�Ĭ�T4'ц˴��ܲ�I���y9�����p���1��V%v�2��2�
&a����ɴmT2�+�"K4�<��7�ܮ����+�NC�����*�s��P�P��V�vU�f6���5
9MK�}�l���Oj��C;�S�z*�J�n+��`U@(��6�O�I?�B��gg�z��$�u����>��a��ͪ:)��n�%w2�{h��A��Zw��>���L�$��@/�޹�+*�6�2�f�@,�胉��Y����L�uו��M��*v�3�>�{����	�2ʾɚKx����?��?m�f�Zݳj �U�{X��__���q>�	���\ �z)8(�5����7ųƣ:m���c���eX'G~���`�=5��7Ex �~��m�ceQq�H��TA7�?k�)zWd�h�>�������\~��ǵ����q4�A��3]��M��U&O?K�-�ME��z_����P�����Fu���:�Ϯ�3�e0)�J0������Ng�Z���iXm��#<LMfئ�j�r4�����s2������*� {������|�����C�F�{�p0y'"��u9g�8��+��I�x|#��δ�ƚ2ٮ�l�6_sszp�6w6�s2����0f��Gu}@�_��?���I�;��f]��d��{C>�#DՉ����Py�<-�$_��MsRh��V��Z��z\��^Jp���y�
{c[�u�'T}���P5�����y+l����N@�Mf1({�wk��h���#�����)^_�ʺ� "`sH����� R�X�V�a*/�$<�YcXv�.+H�&�r�L���P8�u��v�|e�l�r��^l\:]�b���|�� �!4�Q5Ǝ�F����@6)Au����hzUm�J�H�%�$��}-�C�M��ҡ��ɚ�N���Qe1zKN��~sQ��2��\�_�E9�E�2+���[H���� �� �#o;MOs�0:9�5�w�w�:�Y�K\��bM�������^Ǣ���
�\_ɐ	��?w���r�lˣ��[�ju���V��ce�{�Ko[׶:�	�pc6`�?Ə���@6CYa����(�lX3{1��nRߛ{�G�d)_�v��{�Љ�ITʖ��C%��,=wQp�:�(6X��)Z���:�㬬R������D���� 8��?�LMp�p��k��I kR=}g��t�B����g����WjC��ku��~h�#M���&��!Xx��8`F/WO@�	,�`�R����,�6��i�M�$D��W����r� �0T�6�����él�Hy��(*��\c:��^;J��i��̤7\M�j��� ���4x-���Cv�[Ns�)���#�
mb�+
� V�=Z�ju���V��aQ�izP�˞�e`��@p���_	/W!��POD�7��+�����D�4��v*Y��T��%r��(�ⷣwq�)lv�V׀9�u1O��81/�N��T��)_R�Y�
P���w�-�CO����6�ӑd$	j�7.��5�k0[�ޢbGd�R��!�%n�z�r�{]���w}g�u;��O�3	
�y,��栓����^�	�:��̶r	�OD��K�
uR0�D��n�Q��F�l���1��Y_�0A�\�*�s1�& K����ǉ�q-u��>�W&0m�� *O��dӏk��6�)��v��h������;c��.�/N����;��œ�\��I<��hN
�Z��j �U�{X՝�S`��W��Ɠ���9@Io�N2_�-�7��������d~�1�4�t!�t0W���d���Ć���<��G�*��hz�l���2�4!V ���\= {H�R������w��У�����	��'œ���)�6>�������N�C�Q5��gv.��7�bg�+��W��RA�J����:�3yu��V$�1���'j[5V���gp;0;�9Ύ�R�мǆ�\��10x��v���/�xy<�A�*�����πzǷ�=�����)h�l�<���ޣ���VlˬZ��M̭n�&16n�&^��O'�Sá�u�4���44��Y�j���U��Z���d�e`!(9�N�P�zY��c9}I~ڀ8И3���7b+)8�q��Q�D���  C�Vt���``��˒�\��	a�}x]f��۪a��+=���`����� t�Z�Oa�UYN�%tvҏ���Ru�>ֶk�+�W;�@���$f�%.�q���y�>�a�����,=�'�	w�i��jÓ�b�Y�O��������Ǝ������4��^�s�� zeu8�
'Jf��׳��9�� �a�dQg�eHX�W��Ө �|t� u���*�N�$Voؠ1��e he@��|�����b�%�͝/t���t�\��Zy�[�ق���p`�����w������?l�f�Zݣj �U��Xy撚UGxDt/$ ��h�l�*���� tƔ�>!;�p[%�x'F���s��$�BL�w@6���ը����+���󀦕Y�������}�fW�VL-���Eo�� G���!*��4r�@-��i	�Y�8I@��;����t֫�1��A�����,��6�c�ٝ���D�<cO`&e��|x+��b̒O���UC\y����0Mvr=H�\h~u��d�1���-��vv.�G���e�U�)�3��)3�Q�q������2�dd�5AD��zk�G� f���m�^O?_�扙�F��͔=��	�}���27'�V��]5�۪�=-���fUh��OT��m�0�9���Y2�e�i)��Wu��&.�U+�	��_]ڶ� ��\[�|��k��2p�� I��C=/z�u?�ΙN}	�N.IG]�.C00��tNV/�x|Lge��i�ج�!��l����S$��D��Ujmr�t�&z.UpP��d��1֤����<��9N�����[�¢,xH��=X�8t�����E��:1
���h��),���[*�*`�c&�=�e�g���!+��p5�A��"��f2�z�&��q]!�)3��D��`T	�M��,ML������ϛ�Y`а�h�S����=���B�V���m����"��3�KYq�U����u4*7���ͥvsum|C*��.���̣Dez���e�yw����	FV�E9��C�L�I�4�ӗ�]�8I| ̮�ҭ�T. �]���>�X�I\c���&��@���Fj�s���;#T0c2
��YI&c�/*C�ͫ�]>ؕs�9-�
��sLb@Ώ�'b�ߙ���8���7ȥ4�)����Շ����jǕf�K��)6f]����{��S��ل0y����I�8�CG;e�$�����4HN�Y��͠�]���U������6�$:��Շy0��&Bm�I%��P�eK8��[�F:ɲIJJoL�Z�ju��V��aU-'�����,S��d��f���?��58�-Ju�u���������>?�Ê�\����泱g`P�� �9+��xҊ��%����l��ST�?;�`:[9Sw;�VҦ1_��Ml<�L�rp��f�=��z�3��5�}~�w�ۘ�=�A0��+��$�&C�&����e���iba���+.?�z��nc�s�b�d��M��*W�X��1�b��Ҕ01�� �I����b�Xo���ؙ)K�.���e_�$Ot������t��!#9��+߸/!?�C�n^�w4w1�r�U�`ds�U�4��1�D���d&L+"v��a�p�`�V�Zݯj �U�{X��
ƶ'�I�ƥuw��r���6��4O�����Y���Lb�:\�owz"�ҵdJ��
��@Fԏ�DonR��>EӘ�{�u�Un�%2s:�՜��&٪U٤i͆*��!p��q��1� Fc0�+�Qp�5�uL(���
�WE�I�t�sA+cɦ�~Η��&ЪVI�L�db�=WIVT*Zm|5 A��i�U��l�Կ���X��=���T����g�-�4���Tʶ�W޴��
��]b��0��r,c�-4T��U^`l�M��a���	�N�/L7S����G�m�=�rc�P�'��Y��ӑT��_�n[���� n�V����@��nT]
�?�*��C?[o�7O(F<���ɰ�L��?�}'o�����o����e� j������� s�N�`���g�g�\��8U.������8��ͤ1U�g���9�lg��S�B��ْ�عQ��q'5r�R
���^����2���ld�\��P���h�nP����s8˛Ń0r;�-U�NZdz�&/��G���Y��43�N�9ݫ�%����#��l�7)��z�8�����N���P��K7�-����ujF��k0�X{�*#���EE1.e��"�wb�̕����p������?�Ҍ���3�ADa`��'\�~/�TA�kX?���Ə���j��~U��Z��"�$���i��K�-7�5�T�[6[2��->��I������'؅��|��5���/:����C��&1u�WD��QsjE��]n�?�����1��N,�:���� ��!?8[�e�X�0	��	/8O*o6-�f�^�)$�o����R� `�Z��@��}�p�/wWy���r���bj���JcS���g��C�$_���Qw�`��M�>�����Pw꓏��;KkV=}m;�0�I�|�Ɂ 2�n0\��b*�H*W0��ۂ��O�9�E����c�l��+�=|���~9��B�޴����Sm�;R�鈭&�$��W�vbtc��|>��m��U��Z�â A�8R�T�'�\���F'Ve�Nܞ�`�jjs}�e^ISG�\[0;2{Uǩ��Xu��r:��DZR��rɵ��b�#�;����	���9Ack�Jm�ɵaM?��X@,ԎpY�U��z�|2����𜂪%Y��T�r��E�� ����Ӵ�`�a��$�&Ӕ6��#�
�{��oE�0���xC���p�|y�+��TT7<7�N?����&�X�3I^���d9&�9*p;/�]e��NpT���u74�u��D��fN�&�˸aZ����J���|;��uq�G��m��lR�`2�L�a��u	oL|��j�ɬU�{W�ju�>�s�
�̾˙;ǸїsgR#x]#�#���u�6�2�P�8Dh�&�7C�[3T`s~V@D��j-7�7�� (�.��:q��)��N��a�|r�V�B������-��,�#1�=�v4Ov\��\/lJ��i�ԝ�B��+6�������'\* ���p=�7;�+�s�W��K_����:��vY �>��uو��n�Ҭ�I�@w��}Ό�1��N&�!LG�e:&��0�ڔ�r	�,��%1�O=}p㘌���;�^+2���U�K�By~��wc�p���282��X�=�]��S��G��,ȯ�evm&�T1L��&-ͬU�{V�ju��e5�u�^��Ӂlc����u�(��!�T߁i4�S3X�ᇔ&=���Z��Ǚ;�$�P��c�Ù���Q����CK
� ��-:����! ��k���hn��
ڥ���ZMk���ᵺ �	��,��I5̝ۈEK2ˌ=��!�$�Ԏ*rn?��b���,K�XĪ�eJ�L\C9dJ�rׅX5��J��-az�"�4�_ב�QČ�u%�4�|����\}e^�'ֆ>�Y�&���<�'�89��0�2~�,89
���i���,N�,��?�fM���� w�L��t�����������`�q����!��f6�; }ޟ�'��cn��6�6b���<<�_�_�|��o����Ъ�=�p[�������^����E�a_@d�?�ƪ$���y�����H�qǖ�����U�h�ǖ��t$k�υ�r-�@<���8uy�+�_v
TM3,f�`��T>�F���C
�~��8���
�����3Y%�O�XØX��\�A0g�d9�.�Sa=�k������W�`+�iX 8�����Cklwr�I;�^��]*RG@�ӥ���,!�����K�99��k�M2��(}�G��zgR�0��Qۦ�tг�b��tܚ��d�^�7�P��+���6�NƹZ4V6r�nd��:�Dt�f�����Z�*=pwT�N��3y���\��5�&�S����GxH�]�chif�Zݣj �U��X�:��e��X�-�K��"d�j��/o��+e�v��d��>���Ė���������3�c\P{v��b�'He`Z�W��i��T��_�j�]�6,�>'��]W���V����i���W@��2�+���6CH�h���,-�3���մm�'������]F�`�s�����DE�H�80�M�$4e=�f��%�>A�r�z�����_e��,�1�/	sen�!��M*<��AF^����	�x��˘��lZ����b��������gc>-����2�4�B�4��RCᨢ0لȌUw]�y��p��;�Ediif�Zݣj �U�{X�(���?�X�G��3�cvYBy�v{Gv�WmeS�=�
�UZ�a��K����+����!��}�p�.���C_ �f#�����N��[H���K�1Q����w�P�����i8�q��=S_ -u�x�c���d�O�'�,�M�k��|���:cpf#RÂ���ě���	��ʢ��5��N��:tvn�ƛ��t�u�D�]fc/���-~��>�	f�_�]`�h�9��a�����瘪�[2��z�vc;Ǒ�V�^����m ��ѵ�z��Jȶ:h�@��}�Ɇ�����Agjc�R�څ�V�vkM�C���zeC�~��F�<\M���V�Z��p[���5���7�D��u��\��, �Fe����ʴ�I�Zc=�Y����r�����J�#ӥ�hVf� yB���\����+�����UШ*�L���n+��Gz؂�[Ğ_��׀%�ق�k0������5�)�\M^��u���6+����Ã{g (�͔sgNo����\��A��Gp�K�p�k9�<�X�z9�:��m�k��]gM�NA�ÔB�S��N�-��7 �t�3�/��C�1�9���e,v,�@�0�i![3�1��9�H�OL&��OFU�ZB=z�[7�~���n�ק6lگ���{���C*���f��e�V��O5�۪ս-�y�{u�K=!��5�+�dQ�lRe��s��l�U�кT� m��X�Y����26@�+�M�~�� H5s�e�N�s7����$��2��x�2����vr�����n	2�h�2�8V�N��B7;ל0Ϛ���.xm>N�x�V4�mO0��8�<Vm'���Ԇ&0�lb�@	�?����Kʸeڵ)3)��{�=��cc�n��9�Kh!WVz�Dl$�O�8PtDg�M�K�J���u��0��rַ�Ľz��$��ӱ*v�'Z�N�lr`�U\�oN��S��ڌF>��m���k��ں�^P�5MtQ�;���4I�ӹ���=�w����y�V��A5�۪ս����ܩ��]!�!9���YY�����?�����-iÆ�U Ҩq�<�^� ��`-���1�8�h�V|���f,�}�vq���˾��1@¤�tZ��_���[��ZF��2��W��`,	H8r����9�eN�]����8%rB:�~�צ��IFTb�����d�%r���9?�dL�xR�k�sq���RBM~�uH�[W��M �4L�����}�	F$�T ��8�Ӷ�i�%���~��
u���&��my��� G�3�Y��k�X����O|�B:�C����"�!a�+�dhB�[�Mpf�zOV�
������k�|�� ��09�o^��Zݷj �U��X9'���KGo��5=mm0��l,�/��d28 �U�UB����}�j.�_��J��$��Ԝ�9Xc�h� ��yƂ�( ;ڱAL�7��
��؜�|�B$�P���)��.*��r2xI�.ZS�M��u��'�ڙ~�tv�+��l��8�~���������8V�����o	�L*��r���AtT�Ǔ�Zd���W4"L�ET�U=
\nP��f ��.�����v��M'�5�9؝���GT�m���{�i���E�aj��o��%�������	i4	� �{u�[.*$��$£�EYsgѫ�-�َ��9N�k����̶Χz8"������N*'�H�V��O5�۪�=�|��R�Ǵ��'/��� ���5�I�Q��;(�$�R� 
���<��$���k %X��7�YVz�<�V ��H�"X�H�~�ijZ������ZԬ��Óv�^�q��ȩ����Z6gg �F��l�	�8%@�ރ	e��40|���9�x��7XA�˞��@:1�Ķ^���9�q��s9.hw�%xg��E�5��(�x��]���ܗ2�b,��|eyjf�m�|�J\�Q�po�	3��wƽ�,�r�h>�*���o���%�@�PPکZ��ʹ���a�w�����N0<�������^����tѩ/���i�]0/gS6�w�i�b�I�br�o�c�X�y�[tiC��Tm��Q.�85�B�V���m��U�7�~��a�q䷳�&q&Ь� lH�d��X^<�t�N,�gu����(i�#�x�.ԯ6Uk��'�X<��Z�G$�J��*0��h޿�[f72X N6�9�%�Lo+��M�� p�;��/6+6��c~�;0Ng�B�X�}��.%�3�¹A�ݚ�s�W@�h�&Xe`�2|He0��w���絜�*(;-�j��ۊ��S�Y3�D����J/�c;y�*	>����0W�����9[�^���{�$k.\,W������&>�I����BgWU��ڞX�鞢�0�}�aR�4��n�f�4U�`v����r�:��/<8-�kL+1kr?��j{^Oqx��3%5&�Iv�Sʙ��]��m��V��ZݻbNWU��ig��ї�I]�p[�XN�]"k�Ӵ-����� ����}�|F�U�7��w�Z��=�hg:T.	�H3�{U� ޡ�`��ĝ��I�����x" Ǿ7gY���°?RÊ�3D�6k���U�%Ė�-�!X;<����K��� ǆ=5�`����4
����ir'H��^���<�s�ɊM�J�6XT�in]�����i)~|�常TK,���H�`��il�=�����(�x:����	���o�ɇs�~ �h�����K��`�z��,s���4��Jt�-�t�z�w�,|�I ���t��t�i�ꠐF2��ޯ��jޔT͎y���=�g��!&��t51_�o^�V�Zݏj �U��V5���X]z�(I��͖�5��T �`@sT�˟}.��
JlF�5�  Eh���*,�E�9S�7(`��'�Y����mF2�@`P�l>�`��ف2c�,P�묮�z��C|� �}���X����ݖ����:�A}�>��@����q���e6��;���54��.GG���i�]����n����?���@�x�]T�������6��
��&��������D�S��(���N ~[���v��j�29X�u�!�]j �2� ���R�.�����?:�v���9\�~�q�q0��ƖDV���%�������\LN�=�s=��<��V𱨿s��
Iet̻v�^�V�Z��j �U�{V��T?�@}�5��Xǻ2�9�[��_5����S�?�����K*a0��i�Ց94�Ş�H�+-o�3Cb��h���W�����e�7�D������<��4;ۨ�\���N �N%��Ǳ�2w{[��_�z�d���v |˅���Y��
���4}�P�j�Э!��zEfq��| �ry� ��x`C&�i1}�\�;����4�T-�i���؄�R��0K���0�6�хa���Y���H�K~�D�S�x�ڌ�?��E���م�]�SL�pRm��G�Ǳ�����XQ�M���t ��	�"{͙CE��&:�9K�}��Z�%K
s�n�nlR5��.����X�B��c�6�� ��j�r4AB�1G���&���n�m�V���m��U�k&{�����H��jrT6G�IYjYv�S�Gg�<`8�DL����u �\
_`��t������7�M�E��I����g69�ro�h��`�X�����bO����n�9=vww;9lwdkW+�`��v���|��͊���b�>�vl��ܩ|���3��P��եx�%N	�w���a��"Ɨ�xy�¤��߾>�}�ɇ4O��@�kM]��ׄq� �ԩF��ܖ��#�W�� �$/�>�:��
��y@3�ޜ��������������e��ɤ/��Y1���x�9�
4��&�vLgJi�Ǵ���-^�8ݓ�F�Y]���s6�N7
4�9����ub vp<�Q�Qc�� h���gOeq��w�U�V���m��U��|3*�|c�]��K�2KJ:I�� #���d�F%��?N�������}[(D�}UԮ�Tת.
�$�l+~������,D;�4~C�j��à���oE6�-N9�0�d�ZK\.��^�к��(�8�8���3Y�m�Y��X������P�S�bB�0iNi�}�f,���XL~�Z/ed��k�3W����5,U�\1IB��R�� ���f�l�o2�G�15M0� ��ӝ����ff��_ڠ� �.�ۨ����Ie7sm����{�|�#&��� ��&fY�#�d���r��"J�C�꓌��6��\ 7`����Ҡ�p�aR��ɍM�\G�IVR�1�����	J�����o8A�j��~T��ZݷJ�f̐�0��<�!�;@T�%r�S���E/�79B��deɂ�^����@p7���}q�zn�P-���L�.9����c݆��щK�db�¬3�a=m��v`ײ���q���N�gl&�w�=��� ��$��s�<�����.�w�����g�� ��YMř�RA)XQ�	p�0�e�	,���j����9nP�B�ce�u{!�&6Vj��x@�I&-�su0[,Ģo���j����
�jo��U5�������H���@ ��cg����`��v�Ks}پ�74�ęXq6��1�o���c�ݮ,��<�7��� �d�N���38�T��F4OZ^�	����6�$���S��v[�ju���V��]�O�_ڿ*^/�<����m$�X�x�8�_��*��_ՏY���S��	!hG>�-�/�:��>b�����r���-w�k�`L�tpQ4=��X.X�U�㼱�B,�k�*u��,v�� ��Kχ�I��J�i!복�?| g?x[V�� 2��lu�G_�5Ii�ӛѾ����R#<�^����Z��$CbzmdP�h,��q���ꌑ�~/F����ڄ�%#�@QK�hnL����*l� �;s�����%�����8��	OT&?�q� ����/�b�u��c|�R�x�erŨvr�J4�A�6�6'�'f6���H1	�(�dYg�S)�� =ت�Xc%/�]C�/��ewg>�2�]_]�\�����.�U��U�ju�*>�ѿ���Ӑ�em�r&M����0�5��i"����2ف�	UN�
�̒�֔���D${=@VP��~�����8wlIW=n�D��A�ϡ�v�C� 	�n{g~��/c���R��F�P^෤W.� 0X��DRʼ�c7p��W�'+HU�`�����X��X��l0��'˥l��]M�r;)����1ΕQ��{�^I��Jp�#_�Y�"K�e����� ,�@H�>Χ��!	j�?�?4f�Fc��eɢ�"����|DĜ��^'N&KjU�.o�%3ofddd�)�:묽v����^����ܙKM|��*�uݚ�����	Mk���X��FQ{�ڻ������f�|�"�"C~�b*�~&�G�<��y�2f��on_�I��0�C���`6�v�&E�qx�-͠���;��*' ��^n5�����bɁ�~l��C�V��N/�{��ǖO"�z��yCF2K�c���@ pm7��P	w\����\�2����6\Nf���k*���L�������C=Ѐ�E��;7U��*���B�'/��%"�XU~\�����ӂ8.�W�K�倈h�kz1*�kW�Qz�$���@����D���m0'"�Ln�6pը��@��t���4%<�@��
���u��gJl������§[P�s�j�mF�M�Y�s[e��ec�l��5u�,�Y�4���Om���\~=z�{���[��}hW]J�.P{S	%ك�&TE��j��Hz�J�o
�Mr#�9����C��.~���(�s�?���8�B���	�`�m�I����V���79�9O����*���o�?C���	�Ap�k��.ո��Jz�oQY2թ�v_�մ�ν��dAF�%�A2�3�g�!=��[<�~����Ɉ����#[Nr�W�˸ĭ����7
�qR��M�XIJ�tY�����,X�g$,������
���:#��j&u� ���?�C��]i�t�+Y_^��G9�J�J��$�d@�<��5>h���B@^j��Gb�����GK`4^���"(9���H�H"�����6@�Cn�lo���f0+	�5�V�2ŵ�ݪa*��`!}����������Mm�1	B�3���y���B�ݰs�#����	}hE�/���vMu^�Yt^՛%��$Yr�и���q��6t�j��dr����N�{�������'����TX���$7?�?���퇼t�U��x������C�B��Qt]8�gUΔFm�j��A/�߻bT�	��e�v���|U/�j���`aM�W�J5�v2��|�`H{h�mL D�n���ʈ�9E-�T���k�4ua��M��9�����ڍ�/�d������у�έ)�z�<s����3��i�mo���a���/B콻.I���U"�P�'�LY�����boN*_+�J3t�=���ƞ�[�`T%��TJJ던%ף���?$���.�2���2��Lr{��8���f �=�;Դ��Sj�YFY���$���$��.���=�+
�`hUv}�1hބ�~hk�F5��q2X�4�sps�]L�6�''��?�@ pm7���v��������Ή�y����	�[i���Ý���k��;�*__ffk^U�@&5�ԈL&N�@R�堲�}�:vS�A�µ{`{W�M�3%Xɜ�
v��;���Lz�s���KΝ����Z�|�2����V�U[�NmM#�zwH$���Q���pi��t]�}����������:�HxZ+��� '�V<��y�z�ί����ޑ�_�h��X#�,*"���@,�O��Z'9{���>#�����gΫpccI( �f�f���
-.� ��ه"���h�d�2�cc3�w�UgU�.��T.ߪ�[5��k�63{9�,!"wISaI~{ZP0���>!��@��8']��S!�w��Ԍ_K]{d�G��k� ���5����/�V\���*�Y�T��ǃU�[��Ҋs��9m,F�,wp����rnܞP�2��,��W�>���ŉ�b�q����j�,WS��q��mk�n�Pb��ֽ<V�v��*���`$�Kd�Y�$���W�ZrYo'[����.�C�Un��%��"� $�uK�ڂh�v�<υ�m�Qrr��A=
�	�N�ʭ	T��U1'(L`*�
�[�]����Z�ҋv�k(��
����6��0�}ň�A'U�Dn7������jn�qU@����Nrԓ���16����6ආʊҘO;����>���Ш;֛��9άn�l#�T�u����?�a��P~%�p�y�+��k� ���5F��&Q<{��e�rG� l%��'��_�:���QT"�yDXc/T_���_��k�-/C��`�̌f�-7kw'�LD�I���Oӣ��ì��A�5�7�Od�NaE�6P2��8����_��v�HT�kU>^���z��±�F�Zd�*��X.�����52�$�jĬ����R.//tY}:��Az|6�)�Y]k��j��O�Dnճ\k�
�V�\�H���vn9P��v���Iy���+�ڊ�Ֆ�:�ijW�}�Ǒ;_�vi͉�G�V�V�_.�k�y��H��k�Um<�ʫe�8,Uo�D�a����*W��`	�V�))�P��)�TYm£�sW2���S2z�H�CG��餈{ܲP��!�9^C}�~G�(\/��!J��$���?�C�����H\ںDr��r��u���wV���G}���5i��LTbmh{��2� ;��צ���&�ʕEdֱ̈,���2$ψm��@�Lu��,1*j��b)Y�zaA��μ�(�b�k��d�U�&P$+��oz�����d2Mܭ�� $U��(f[�{��5��6��>%�N8��-�ʩ}o��e�XN��՞tQ[�z2U	UQ_�i�� ��N���;g�>�%�ml���,jCpkI��-�X�X]�a8��-�Qd�~���1R�s�'w��mݦ�u�{.�X���m�����u��{Ǽ�S���F�5�������V]����L�	���������j���$R?�/\Ș� �#�5kl�մm$(�Ap�k����6��nFd!<���2hqT"�&)hf+��ވm�*�>�����ex�����('Yi�뫊,,���'����b�'h=�U�o|ٞ�*�Wo{S°=�H���7WI���DO�0
�V�4�6m���7o��ZK���r�Yk'3#?�U1�k	r۴���з	1ex�,��B�����TE%��v��E_�>�f���vv2��OU[d�Bi��.�W�,��^�΋��.Ѩ�$H��k�K�z ĉ��^iS�$B�%[B��#�e�V-��&�,�����7��/A��6m<m��uP_-��4�L�U���lp����c;��ͷl�0�ME�c�ꐋ9Vjo���Ε�|U��t��a���#x�#���í5�k[�$Ɋ�8pi�f�N�x�L&��\3��%H*�3�%����h�� DmuP�٘�Lq��`c]�d��2�)e�x�ޛ��*.}���0m�(g�l�֬�$N���D�9XWo���ɴ3�C��WJ�Q�t0�&������;*�+������
�z�������� Ȇ��&Q[��:Y��	Jc-m9I�Z<�⾖i"t3������[ӃYv��-x��P{�׸&��li}�mj�k�������{]���lc�~�sWj1��v�"��ИC5��I�`8�Ӝ w���kO;X^�믃@j��|������{QǄC	$S8\��E�l�!��l/,��Ufa������� ���-\M�L�s�M�����IU�4���=F���[^(ǵ��V��~���#Z�H�'��=��@��!n pQ�݊��"J���Y�{1�DL��{�QLdQԃ���3�
�� �J�Z_�6�+�4Th������_��In����2a|�b�xnJHQ|��C��l�VMDpr+�����/�Z4�)k;�xV���,��v�|�LqM�v��^%2VWބ�"A��">�<�W��|Y>_�*�S-p�eB0��Qf��\�^{������eG1U^�xN	�I���Q`����Qf�[v�e�j��8ӫ|,it��M1�i�[�����w�*'����X��jei(F�N��K�MӚ��i���3�a�S�pvmm)=nz~٭Ӽ��F^�B��@/�{dk���j�+�����O�P'bǖ3�٤�r��	�D���G�B p7�Ơs��B�mV#$��^M�V�?��xS�GL䶿J�oc�T���kk��7)�V�d�-����[[� �Ș��x0�/#ͪ��+��YaN�-[��hNn�`!U"�ô��+'�\�W���-���� ��2mWZ��6�P�-˴�	5�pW�{�ĕ�c���sg����I�KT,"ro΢��|U;�}G�p��/���-CW�c��2�ͤ�":'����9�H��n˲��G	`O��y�Ua/��\��}bҪ�V���k���BEe����U�3M鸴.n�t��asʸ�ﶂ:�U�wH~����F��n���o3d���s��3[��& =?��i�ߨGm���p���vN��"���\�o���꾷�ַ��@�"n p��ezs58�'Y���JX��	�d�7�L���x�|��f�6@quۭ���YT�C.�+�HP���g��t�L��w��K���ث�J�@n��,��k�8
)�J���k��?*��o��1�lۥ�j�ݠ�w\#��0��V�k�߲��6Ia�~���d
d��P�㵔4�V̤Jx�����i{#U��Eli;:=��֕qD��l�<����b��ĉ]EE�P���y�T~��[+����bEkz�N^\�ĤB���*F��������1_e�4ic�I	TYm�_�^�g��Z���kEK�Hr%��&l��\W{+�9�F"n+P{?���D���8�i�����V<�B�9&c����C�@�Zc$㺨�����Ή�W�������z�%4�k� �&��mݪ
����D"&�ݘ׶[m�KU��{��VF�� �L\&nd2����AQm-붂�va����P#�K�XJ�֝væ��vu�x*�l"_����/k$�
�H�I^v�ҿP�����l��60�̫�O���Z�Br���җ��|�>}fݖ�3_MQL��������b�á�+Ԯ*Vy�X���߉ǳm)��m���wެ`�<Ox��h�����Զ��s��Yy[�"}��������ޚa6Vm4�Nb=�?;�b���%�2h�(}��Qx�l�B
� *3&��c�"T^٩�Y�-���?��5B�@��cTF}]_�1��9CP�V+�=�	D$ĺ�a{�.��4ãk�^Pq���Ā�ౄ:��D�ڕL��*�����,�;�� �X�&�NW�>!�

\,M��r|��}6���啬�{w�a�k��>y*Uk[KdXx����ն��gUnv��*ǡz]�ЋxBB�Ĺs5��!g����yF�z��=99q�ݸi�Db�Q`��
��m��A��(z�M�Ǎ�?���)�J��i	����Qv[�����[{�ƒ)���U[��k[�o�+t|[fK����)ky���R����0�̋�z�X�qs�2㻨J��e₟�;!��X�[Y�b�"�l� �/)�\U$���c���|��$\��#H�� q��@շ�Z#��F��B_�V�`��U,���'��_�R�Z��*�X*�.���^\���*�?�T��Y�U��=GA�`m�o�~6��d>Wr���M}���$Q�l9����km� ;C���Z<�W���n[/��L����.=��8!���;VA
5�ߗ�I��G`QEk�4m&keM=?'��9<:��ï���}�'*�H���Q�7��~R�g�bǦ�yp<o}��d]篝) f	�e���1F�TC��3L��ƧV��>�M�˲�u���E���=w�m2�NŹT��N<�X<F���D]E�B���#�/I0*���q_���b>k��z��'�6��~�,�M&]�E�����C�@�B;1�{�h&%/$���}�2JH������kg#	5�a�e��ߪ��˴��b��/��f"? ��5<�����ok���'��m��r)WWWJ�dq���P|����N�[%@˜�<����ƨ�|T�su���&��CT٩x��܊7U�dP�>)C�ct7=�C.x�W��������1�h��i�_�x�U`��ɷ����gk��l{��/�	��%D�z��R7f�*��2�4������C"�Ei�i�����2IW�;だn��'��Y���@U�=�ھ�c�X�V����*g�j�;x�䢁�0���#�XD�|��VSy�uc��\�#���/�a���ZI/��H �~�\C0A4g�j��F��+�����X���SU��J�[���Gz<+d�t�ʃ�6�I���#���}�kt/����
~؋+�BqUz���J�˕��� ����⫗r�e�t>�����WKY&b�����:{���������9��#�*\zQZ��F�Ǩ!&^Q_�#+W��rϨ�}\'��5��(�e�V�B�r�o�t�\f{���}O_�H��i����.K��W��U��\g�iNvr҆g�j����jў�2��y�}T�Er,#�r���/]鱚:����ZE�N���l`i\I�����g�g"�%�?�*��n���L�2��,���:0��$QK�6�����v.yR�l�L�K��c�C�i^�����KjOƨk���b\G��%@$����w�	"��g�����Zhd�T��̮��^	�*[��B�Κ/���[���%B��Z�r���K4�����Z-HF�L�2��e6��t:K�v-o@dӦ�i3��Y�,���(�%o�moqn�\�jHB@�1X���b�k��Ϭ �i�kڎ�	"�@�Z�R}sE�N��_�N�S��
�}B+ڪ��m[P����"/�P�݃����{��C>�G_�ԙT�ȵZ����G���QѧD<�rI���럡�<�`���!˛�:�O�Rs�sݛ���Y-�L�M߈�Zp=��
�*��U�|��K�@�cn��	N�mx73- �x�5s���uxL['[��F_/s�{Zq�zƝ�ۿ��5�![5��V~�������	�f$���ퟦs�.f��5D�@�BVg�\&���UU��i�"��-V��[P�E�t�^�j�Ѹ�5�����P���E|-�kެVrѭ�2�U�ϬЃ�TXQu��h�n��Peg�,l)�M�3M�h��&r�ZU�:}jMm�M5��� ��<�K�/�b��>�D]�3�̶�-Tٯ�J���z��W���nW�w�G7�C%m?j�+���V��� ~���RQ��4�Ƚ����z_|�2��R��絎��
�zQAZ�s}ݕM"�恗l\����{�3�cG�X���H�7�t�yH"��u�6��^[%�b�YQp`'��z!�v� �����v{W��R������W�q�j#�T��(l,��%�;y��{�W������i"���''D�@�"n p��f�*��3n݆0Z
#��$7%P�r���P_/���VJTApW��(�EC��´m���H���JiP�y%����SUa�ނ�N!�E��D��>�Dd�W�Mg�����3?.^;�̬��o(tW�K%���:s>[�r��v��꠸� �=�~F�ܷ��^�'t�VƆ#9���V��2¨�M�1d��Ec�ښn��Pr�h1*�ًZ�ϸ>*�:R=$�-}���-k��6s�Kƃ���⺯��sƮ�Q�8�m
�+�=�|�j����qhm�qm�hܵL=YB).����q����=�����:�;TU}�$X�B���ok�y]u`�����/�����3�`��V�0�����V�k��P�ê�$M���$Bp�k� ���5D���Ϊ�Y]Nre?�\g��� ((k+�K��yZ��Z7%�k�j5�	�\Ӡ�+��u��E���b!��d����&�0��e�H�����J`-mk�,`�� ��F��)V�5L���|��,v���s�,e��_��5�k4k�qy�S����z,%����֡�}���Ո5��� ޝw�kF2��s{ϡ�S<�Q!$�oHX�N-���I����dÙ'c,!� �禮>�L(�-h�7�@�/K�p_keJq�
��Щ����e{LU��V@�U�Ez<�^������]�w۹�֢ͬI������`Jp�-%�eo�iW��W��,x#�Zr�]�7X�א�'��q�Hp��hF�Mҵ���@�"�u�%�Fr氊��k���w�W�[��޳a{U�V�+Y���Z���D���m.
��
�%?-��Z�m��*���d�J���Qe���c[�1���5�T������lj��-��U#'-	+�Ŗ��I�)S�v��TNA��5�G5��.?2�`�kB=v��2�&�����9�@�	�xl#�bY��/�{�B�[.�}�aT����l/'*d��{�-v�c��To��?�c٦���M�{#���'3���t�`�>�z�V[����M&��
��F��FS>0Y�k��V�Z@����J��Ak�?�'i��~����;c��1Ͳ�}�8��jZ3�iRo�?a�=���!_�|�9f+nä��?�@ p-7���zd�^]I[md:�+mڀ��ծc��^X�Gnh��g붕)H�+���p��L���И��A}U_��o�;��,-k��*���~��L��^�U�EF)��B���%yg��9.w��.>Vy!�\>֐	��#11�7��V��o�̒��S;q�-��PG�g�,Z+�ӫ����ڪ��o�)*�.����zW}�ʨ7Ƙ��eo/mSa�8f[^'?���k�/%wCa�֦P�DT�s*�%xt�v���O#�-�omr����q����n`z���m�[1�Sǋ� I����7� Y�k��u���~;�®]��\]ں���+O��N��"�k� ���5��z٥m�ցzb�K��a�YsG]����d�)l[ka�*���a�b�o����Py�U�fh�H��2?'	�n��i�J)"��l��6�����l�K1���Z�2eL��7�!���b�i9��:E^����\�#�x9}�*>WEnփ��W�;Hi?p1W�]�$�<^�Ӑ�OH���<��ZL&&U�RU���>M*6���A2;wE��J|M�f�W>>�o�F��DF�F!angl�	�zT�Yx�Q��1{x�s�ǐ>���;�3+&�ښ:['4iV��hS���q�ڎ�ٽ��w��E罶�����#���~Z�m$(�Ap�k��Fk,+�?\��0,�^o�ٸ����T����_���^)��&�sXu��&�4ϳ��.��n�<��<��F,��gk�}�2�lܶ ��h��X���PQi�b�\�30���c�v'�&)CA�4� ���c�ڭ��ޛ'$�&	wrVUclօG�T��}�9H��s���	�����5%�Ϫ����1�W�'Ο$�2�Ƹ�!+خvW%��W�[�.�ףD;����Xu�θ�_����'Kf�RMk�����K��j����鴘l�����`�&�L�e���b��u�u��l�<�ڶ]��x߭Xd�d���x��n��we(o�b3�����u�'��=��@��"n p�\^�jy!����mΥ�`�$r����[�@([S�Z�S26�
}zbś:�r|}q��[�v�
W�7s�J�+�$��:#�z�*�-o7�K��+HR�G�$u������˜�Uoe}�x����w��}ٚ��c��2zm��U�S���,X��bQ�ρ���Tx�Zr��/�3�$-��z0��?�V�<�-Pս��a���܆�1�;?0ȸCV���^������p����_c�����Sr��ޒ������Q:[,�غΉwD'��w֛n礱�л%E|xA�]���͘��U�*@k�����^@(^�6X�]��sM$(�Ap�k��BպH��|-r��⠱�-w�N�j����$^��w����q�ʊ��������iuI�U�F(p��~��fղ�8)��VFD6V�D��d�N��Չ/�dh�d�d�V. f�>��ީM�]��^�ɡ�Y�4\<��-IOާ�� Z X�E��}�o�ȣ"��w@����r�>_�ډf�UO[�2_�*��-��]bB"�.���5L/��U&@��ڤ�أ� ��;��*�����cܐ_lߴ����je��Ш*��T��q=��I�T���bKt�Z˰��č<!s����\�h�:Kc0{Aퟝ�^��Y��vj����[ӕ~���"�ߍ�R���\gĿ�@���N��"@�[.e���U�kVH'�H�y��X��eվ�1��~�A�g���f]E!h��������r�J�x�P��&<x`�`�Ъs��v�,'�Z+�V�jL(�e&'��!+��M�\=-��R�n�K�e��`�X(�,��3��a���x'֣��P�q���?+�M9ʏkd���Ö���I�_
�R���Lm�jTo���)H�%�?c�����$�-;8�6�h���+�����H��w��y~�j~q�׵�.h��_v�[�_^���R�}�'B��|�m��O�,At9vjksG�V��'-�m�[���x��VD0�L�����f�M�Ӂ@��"����2=I�����Y��]�݈�a9w�V����hU�H&��ʗ�e�0,O����㎢4(S�ݪ2�?��>�m��km�K�ha�z%"P��ʕ��ϾѲ0k� H^��&�N���2R2�z�Na�k�*�B4�M�e�}_��8vl��uK��1k���AշF$�s$Fu�	���/��j>�k���9g�X��WWe���ڴWI`6�y�dwt�H�|�q���u��}iO�cU&���b���R|�������R�yтB/���f�:!v[A]!���U�G70&�_�N���Me2C�Z��wq�D�o����=(�Q�z,uyi}��$��H=_k���R�ME`c��N�Ӝ,�'�_h p�x���_�����û��(�Y��+��6"&1L�f���=�R��lU��T�Pzg�P7b�Zf�`ǩZ3\-��CE<�Sݯ�N��h2�.E��Vy@�ܜɫ'bK����`$MN����ebQI%�*i|�$Ū��8�ԦP�����	�S��2R{_ʦ��$Hɴ%*0��O�S���%z,���(��z;�!��)Y�{W����da��Q�3���{�R@�<d��
nOŸ ��_ߐ	������Rf�rRcפ�'"�㤱3A$]��t��X�4+�켨PwMϡ���$M�������M6��!�@��I���-^���B��j����}�!���}�l��.�4���C�@��bzp��D����x��s��z-��F� +dꔠ!`�ID��I�k��4�i����+��̵�aC���&����LU��ŵ�}}]�Z.�r�\	���S�e�O�$p�����^�y�N�*�+�FZ�(V��ܸXY��5�WG���U�S����������$�Ml�%���v��mkG���Y�̈́�(Z�C>r�eɠ����*;)}��0��N
�w|�֣��QI��]��^9YtoK�T~}�hZ���K�Q�n����N7ml�mp���[8)�&FP-�W2
����i�Ej�����WOx�pv��~��/H���6�3����&���q�ގ�6:��B�Aǩ�������2M��Wn[ݚj"��ct�������1����}���7��I5��7�F~�~.����h%P���^��~����ʬGmPi�Z���\]��Ol��Qb\��Օ,2'������<�\���r)K�m��jc�F���6�h���J��X�U��Y^n�NT�{gI�ؔ`�$�&�^_��R�I�gSHL���>��5�_�%��9��.ZZ>��}+��$��q���$���Gk'9��v�A5��G� \�<�\Fw��$�w��sN�0��$��v��$�eFp>�A��hPk8XC��9��G�U}6��8��f��J�5\�K���=ƹ��Zǡ�|`�ca��ba\���Vt�$w�K����I��7=�X�Fp���Z0����c'�������,��>],�?m�|*�@��"n p�1�O/�����;��?\���e�����+��u5��Zi���D��+ɗQ�P�-
�z0�Nd~����%?��>��fobz���Z�6�Z�
H�3����G�#T5�V3v�l�	ս)�/fM����v�\&��a�[{���J(Fb�z$1��֮>�d�l�\����,�Yi�F3qr+���~'�C�"�W���A��)�+��ܖ��-�i��0�y��5��l�U�՟�s=��,��N��V�J��#�l���bE{�����f3,�ܢ3�fue~��}W�Y���t��v��N�]�?�:��S��Z<����F�LͰ��V�������b�4y���Z�kD�A���|�$�m p�7��X<�����~��v:{\���Z�w������e}�&�+���ke|���j׉���و@	#��{p��$�(�J$���5��������ĩm��8�b�<K��%gS��=�ޗ~��t��I�	�Nrsq��{��ֳ�*���2oCU�Gl�d�j[��X,�P�E3��*���
��73I)����!+��;)��?���[�,�:�ݑk��6����2Tm%�,@����k�����ٶ��������u�����)�,w���8���sTgM��d��Zmr����K�4a4��d�8�6��\֫���>��]�:���ˢ(�/l ՠ�a����,>���=�^h�/�q��{ڤ�L�ve�h�0��"�6� n ����G蘤]�^}�O�XV�_��G��[go^}%W�Y^H�Y)��vy�����J��َ�˺���/��������&��\���2��j��fХ���@$[Wmu9w�*�տq;��p;�j�#y�YaW) ���")%����!㪊[��U5�.�u2*�L�(	�h| ׭ܷ�}���:��I�]��K�t&]��3��EY�?�sr[l�י�����K�K˖Oܮ�|ſk�V�_��3��Ib���L,��⢳!��^^�n0�m���U]��'@H�L�
��N�f���۴!5����3�-��T��zK����ߞg�b�S�v��N�3=n�i<dh+�`�YԲ8�%''2?:��@�;� ���w'���������j�7�����\�z���+�\]&"��%ܫ�:��Dz�yl�X��iX-�����zb~�A%���&7IP�+�E���1���V �@B͝��2�O���V���:�P���q�Mu���jo�:*��	�'���������8�dH˄����[M
? }¬���ٺK��c��*�GR����0�߻�<�a붌{+m�3R�S,�9����쾖�+�Hߍ�������z�To�F7܊�y-bbTsQ�V�5��A�( =a9[�q3�7���z�FW�̂�N��$�ȽŸ]�����M�8�T٘� ��$2 �a0�W፧lTunz2�Z�� k�A��M�rz��,NN>��gQ\|7������}��տ�d6����t��>��^������%�k�is�΋�l���Ϲ�C��M�b��v���.��D����g�S��,��x6f�b���4JTf�U
��п�����is��̎�4wh��� �I�v����i�_��P�ba������Lk��X�|�Z��-L����X*�}e��rWE�T�QlF��W�Ĳ�$�c�ָoIlwI/+Iq���2�n�o�*lN�	w_�[������6��W0��K�o���ц{e��e�o��-V`�Y��j0I�c$HY�Ma��-l0Ec�/T%��ݭ�jb�z������@N�m��1`��np�k���k����䄩v�[������Ӧ��d��{���|�1���|����~:��:l�U�g�t&�/����ϔ�tM�[��5�ѭw{�,��Os��M;H����[q�'��_P�<�t�M#t��H�
Pp��2�'����)m�TC��m�Ժ�Y��`��M;���Tl�`��J���t��_17u�ϗ�Q�!���U�_u7� 7��+g�$�|�׳���ѻ>d�1���'�x���Nf�.�XW�m_ln�@���[�D����	���VK�u�(k��'B�Ѯb
'��"-$S���J..^��ŹzhAr�˫��RǓ���5p�����u\y�����	Ќ�������z�	��۾��|.��,�~���Ę�����2?<�&��!��ĸe~���O���'G�������8��C�,���g?���&�ɏ�9{������ �)�F*4�@8�H&����<��~���t�P"�%r/$
զ�%�^�6,�����KÓ��a��P����~��F.�rq����CY�6���n�4*��J0L��ͻ�:���nU����lla��� `d��ʏ,�,�2g�,�r��Hps4U�����jG��F��:�J�3Z��¥�z�-��R�
��p�6ZF�aM�ͩ�h_�9�^[W���4��-�U��# 	A�蠶�	��*߫��n���ez�J��e����Ky��Dtϕ�9T�v����n�`2U?7�+�����T�JW�!g!RC�� ߖ���AS���\�����8��-k&�p�I��P�sGǲHl	�t�i:��5��Ϗ���)�nn}`Dw�՗O���_��<��g��H�WROj�eK�u%S"�(�h���2.6�����#0�-<C�gbﭝ�pL��q�N.�Hb��ҋ�Db浪���B�r�8Tb=Q�d�}��
r��_k�騤U.�"�V�Ka9���U���ӒH�G���c�zʹ����ܾܷ��V�f~c�!Nr3�}��V^�fg?O��F�k�4��<���y��D����[�v�l����(h�qk�Y�i1a�q]�a-˫���:�W/�J$����}��z�B���\^�+�Gj�&<i����D2U�?:9�E"��uS&R�̡�"ȕ��8[BB�j1��p�����A�M�������ID� M��7i;���S9�}'M��d����ѩ��M�i7k6�M~r����s��0Lo���������dr��d���/es�Z	�4��De5	�lR�5j",���������U��u���Z� �6U�<���f��e����\���e��0c����*q9:>��t;KS����+���V��F��#���.��y�\F�J��E^�0�"�].���$q��f+�p�~�YYe������??1�����}=��aT]� �J������1hV�s-�Q
���Q����Nf�&�o�ӊ]��E^�4ʋDpA&/���JS=���e������M�&]�rrz,�oߖ��#%���"6���#Wv���[����<QR�b��gh��Nv�ȼ5V!Xt'j�8s)���oߗ�����}�}���[SsgO�v���m~�ѣ ���wAp���ӓ�4�4�{�-��M�>��?����ҬEfU+([��霶�D6���X	��������B"%æWB�
sm��9��&�Y,k;�lz��R�C��JT��=��N��֭�^G��A����*Y��4C��	f��Ɗ���l�j25���*���c���JV�	d$t�[�W�P$���z A%��(���;8iF����t��}%�Gi���a��h!?o9� vu]�x|U��|�_38�~ۡ������P����x	�;�D��1$c�I�e"���Wҟ7r�ԃ��4F�J��4F�or�����ܹc�b��Gz�u��*@l[/L��@+�Vfz<<��Ŕ�o��|b������j�T-
����|���i,ށj�4��'�@M�>9~�Q�@� n p��}���_��=I?�ݝ��}������Pm�ĘT�m<b��,�/x��D	����
�c�>wDS"B��ɨ�O�p2�[w��i�N��UE�U	�v6K���Υ6v��2��Ԯ��`/Ƃ�f��ds���i��:bpBZ��\�Ŏt����nZ�X�W��.�q�����h�u.垃���2J����
�Ϊ����_=���n^����z���9[[�
xv�V�D�gm�g�$�:�'�98���~su%/ߜ���R��{:������r��-9X,�8�ãC���-̢6kKg���7汭8���?��X�=r���f�Ԭ6P����Z�W�T%�}�y��#�}����[��,�O'�������7Ap��{?��O����l�Z�����Ldc���L�u��S"W�%�D�R�X��jmEb�ܶNv�Jr�vu�-S;�����xT�'R19<��i�J��[����9�}j���2.�[��n�*N��i,0���T���G���D�TO4x�eԕ���lW���dP�����S~����U>�?�Q��?���g�y,{���Ɔ������C�F[�5װ�<Z3z�Yh"�O&���`�mE�@�>fm���24�DpY���I
�Ĵ���i�sGNNNd�Ԗ��L���v�K�A.2;�5�䖗��̪�FJ��Mn��q���Y#}��X�ޒ������h}�&i?��/��(n0��7����/./~t��gˋs�|�B���!,���t��~��ܖ���hc#Zׅ��ZIN��]N�� 
d���%�4��C9J��$[�bix�>ߙzk��I����]�Z�M�V*��z��vmc����Wk�Z6����y|��f>\5�Y.���ރ-����$�ފ����������%��������,��v�>��W�3��g�W�������m����*M������,�vv ���ߤ����y~OS���׭w���}��Ź��F�����|�㳣]u=]�ѭ[r����O��?���ã���<x�6����p,n��W�����Σ��勯���v�����F���x�z�"��/w��t*�t�h/|U�J&Z�^Y��ƺB!�	U�k�<�����ܑ����?M$�I=��P��\b6/����:����=��-��Cyp����2��W�~��cQ������W��ߧ�}&��\�&�GE��)�ŻY��Hp��Λ}�oƟ�7���m{���U[*ɥ�jv�{�.x*�}�i"��O���n �/��\�n��@��qÕ�2��Z�m�����ҭE��:�U��6���8�����i,/u�����I։���{��~ �w�~zpr���{An�}@�@`px|���r�����=�⹼|�Lm�H����B�],����BVo.d��p0�
�5
�z����4hg)��Ea��fӓr�{���?F���������?���n��@�?��W_<�E"�����C�fx��9y�� �N���i��"�֫Ux��������~���z��,�i2UuRo�2K�u�[��UB�bv~~���Ak~qUg�q#�k#���hqy�m)�4n����壿�K9}���u����އAn�=A�@`0=���7��ߟ̏n�ՋS���tiq랜)I9]��ԥ�~�R^?�J��FfӉ���C#��F��2��*o���t|�c����DNnߖ��ٟ˽?���]�������T|G0���G�/_>�ٗ/^����������7����ݬ���N�6i�����5��qs�*L�����x�^D��1�Z]e��v�˵���D�|��}���ɽ;?����q���{�����t!��C9�}O��:�}$�OO�n��٫�y���/>����Z�;zuy��ʫޚ8\AY[w"���y���=9�����[����?9��(HE@�8���o~�o?�{���$��}��N������J'S=��"��EW�Df'��c���6��I���$~Ti,vJ��(_$�ܶs�z[�4�M�$�m ���	��A���@��(�>x(=���#�4�V�X�"��2�g"3��NgV���\MZ� �X-�]/,���9E$؃��������An�x���>�������𯏏�����Յ�)��i�t$���4F���{��`�����4ޚ4^']z.M�&˕4i�^-������2?<��J{��4'�&�Ap�=A3i�TM����;g���O>����.���/_ɛ����y��\PKu2?����]H}rK6���t.�ׯ�_wRO7����]�����=GO����5�m୸��{�������ܾ���_����:m�099��݇� �ѭ�i�͵�
"�ǽJ�u@�ֲt���V./.�u"�k/v|��e"ʇ�������i�X<�@ �w��	n߹�����������mrO��Ӧ�/���^���>��|��<��y"��8�K?;��i+���L"���Z%Z4說g2=���������	�,�q|��d�����]��U�=��#y�������H{{\�sq.닥|��+��;F����r�����������(�v:�7��N��~�=Y������@ �v���dR���vwB�>"��Dr�Rɛ�J��:��}�\$Rqr�DNo���c׽5E���l��8�w+���/U�}�����lq�Y���N�4�ŏ�~��?���+mr��ݏ�Tn�(��F^}�L^&�z��/^˯~�;Y�����C���m��qb�i,�&w��B3�u�/��O~1[�����D�@`���_�F�
�Wo�!8��|!'���������E"�ϥ�� �V�m��Zi�2��w�b�(�z�I=���[r��}9Z>y��A(f�?�������?��O�'�}����.�Wr���r��L������˿�Z^�x��	/t��w���\�4~�(�`踷\�����{M%����ɇ�	{� ���^� f	$��[�=:9�mqx ��\�q'�7�D%���^x�.�ҭ��m����<����Hf���٤�@�������_���=9�s�l�Z�|~�c��չ��7�����7�E�������Y4r@<��c¬�[���������|�g���l{� ���a@�D����L7m�ZW�Sx0���M+��L�@l-=a#}:�d�0R��I�V����vZOg�ӉԲ�qv��\�6,WFbCw��m%���N&:A�E�	��6�+����iguU������@��#n �G��kⲉ�֪u��F;Cq�6i�0Z�&� R�X,�H�|�R�H��Ve��h�?�z��y�H�����Ass�h��N�si5�L���X�\��l�`ʭ��h �I�b>���~���?�$7�C��	` �Pm�&�1���m��PgApA@"@r�n����Hk�����@��q�q��e���[��ч:�z��>�[Ko�W���-
� ���j�Ǔj8�l֏%T�@`/7�#�����C+☨̒H8a����s�@��8��f�4�	
�?g?$���޽�d�`ȸ�}����"�cb�J��Z���b��$�%��{-ȁj�u�܂8��K�$���܇U���H�Ǿ%)I�ɃHP�҄��آ�d����T����:>��b���@n�/A?96�����D�@`�@K H*��6�]���d�I.�0������Qb���o��ogi{�0X_���c��0�Ul�_N��&l mDi�	�� ������,�$�X�y(��$�$Tذ�}����DJ'2{�1��S�b0/�/|��Tu9V99��ˉ���/��{��H���`�<P��$�\&&�(	II��w'KTaIHIpAn�q���_�i
 ����O7�o�/R �G(�� �Xέ� }`�����m�X(��H��I{��1xF���'No��7|��]�􁱌1�K�������!n ������ �J_-P�����TqIHh�]J�dX�G�=�����'�)�葊+WX�q�D�Cm��c�m
-��Pp��F�@`��}*^�D�-X.c��]�dLY���(�|>�c��^�6�,-0�`AZ��}Ks�@`�7�3��[�&'�P��%دT٨�R��B�]AK�K+=p?-n1.9�ʤ�Ǡ��'<�o��{�Ӓ�҆@b Pc�^��y�C�[�;�Ғ�Kp�r��	
�Ҕ���^�O�h���"n �GH�/U/n�"�dLP��9n܇>����$��$�e&3����V>�D��iD��@`7�|���g��珡�Q��V�2��[���ģ܂L��o̐�r�IL��8,�1���������� ���� �/���.X�-��覲p�$�2����c6ll� �-�c�,�j�聅�xm9!�"�@ 7�#�R�X�G�:�DƢ��_����x'��b<���EJ�[Zev���Y6��,n ����	���t�I"�g�K�$� �B���,��}�i�/���~�@��l1�`��t�ru�l ��*���+,HiN��N���"n �'x����_��W�[*�@F�K��.R�wW;??���O%x@��x"��ĩ�L�-|��1��4u"�[\��Dx?{����ߏ����{�_���g���K�h�PV����1v��5�E?%� <",��w���eOb{��m}��ٷ{؏��2A�E�x�*�{v1�{�v������ǉ( I!/S-+�� .�{Ko$��o,�>�/������}������7��-*�=P��ؤo|7��r��]���v�Ap��������$e��{H(���]��(�	�+}<_̱��ōe�-@e���S����1u��v7��-��$�X�%�$�l�
�?��	�Xt���*S�-��x���|\vЋ�e�@`Ap�=�ۋ��.22��<WƉю�[���,HJ����Ν;r��-9<<�ׯ_o?�$���r��1��hW��!T�@`�J�������
. �
�
���͛V*ex���Am0�@n�����mi=(�-@;7�Qznw_�́��"~��=��AJk;EAE+� ��`��2/���4�4������ )e�c��LŶ,�,m7ǌYN?Mǈ|�@`7�#��˺,.c�(��px䖤�V�h�x_ ��?�����mz����8��$�Tl�<�����h���{��EDX ����	��j���ނD�P��`\fL���Kr��@�]��Z8LL���;2���
er=�,��&�3�S��%�%)e{^<R���_���%�ߕlG���/8�8�0i�a�����4@�[F��96*��Ap�==��.�ņ��ǃ��=��E�7=�z�J��� `,bL���>r�n7jϗMJ��~"n �'(�/��Ò�%a�XF����b��2*�j��l�@��]�c	�_}��\���h�y�3ܖ���U<���@ ����@�n�~��a��XDV�Z*c$�ZɾZ綨A$��0����0&"p������� >��\?�'��{�Ӳ�n�1J��.fTf�D��t���p��	XĈ�Ʈy%���AUڪފc�I2�1��8�� ���� Qe�$\��V��eu��c$�\2����IQ�+zm�g�]�`$��<n9���� � �h�U�@ ���_�@`��矟%�J $	eӆR�%Jr(iZ�N�Q�xo<{��,m�QPV����#Tg����;�ͳ�K;-���b�	�Ap�=@���~��H��n��|���0���J[��ҴM&����+�X�qgl:�����@���nݒ������D%����v��>n�y��et1�Ap�=@"�]�΂8���Tj����96x(rp���	i���r�<��]�H`a18::�$�6��Vu�e�a�3 �7�'�&�@`/7�p�e���薪-�]�B!���4݆Rx'��n4~Π�j��Ы��9�e!�Nf���P}�BH_����@`�7�3�, �	���Y�%�_#�e�+� ���i��L��-W��pߖ��.g��2���}���"n �h
B�۞B�}��.���$�V���֫��f/�Y�I�e��.�����K��w��m�M~-�.��@ �����wL7g��~¢Z�/��R�?�ĀE:@�<��F5��K�-x�;�MC<�#�&W̳�������w��2�i�n�����
�@`7��Y�\��e;}�$�,�a)���v=���7A�'6�@RAlvܣ5A�5C���x�6� b���{�D~�n>a�S�U.���~G�S�ą@��B�,��0��-��0&x��1w��Pd;��D�@`��B��X%�U�Y�A$�u���ǡ�����.�����1H�8�hW`~3�/'i���^��@`�7�Ђ@�A���͌$�M H@�O�C���F�f���+g � � �x�͛7jY�$��]��2F�l?�Ap�= 	-�-U1,�R�r/}�$e�3�1N��7Ů��>�m1N���WWW9u��x�r|���@ ������O ��& ��K�ܗ�.ޚ��8�b�^�M��"G�S�(p�ƍc�jD��@`�7�$���dK�X��jFKڤ�\@��kM�B���li��x�'��̴�`��������Д�m�@`�7��x���ً/��H"�|A���-[����TyA8v�q���	��J � �Fj/���޾}[NNN2���$��gƸ�q�@ ����p$��8��3�g:�v+λM'���@fY�F�6�aQ|[`2UZ��AVAf�ؽ{�te�����^�������Ap����Tɘ�@K�t����6�eQIn�?��A$�%Y1�c ����b��x�c��%H1�n �_�� $��@��.H]�	�!Y�Îg|�G�Pq�; �\1 42�ի-�[��U-mc� �.�b�ь�0:,�'��{�ݶ�ѧ�^G*ie���_Sk���-P����6�LT`$����~���2�M��`�b�x����E�@`@�"-����@��y���^4���m����[� ̓���}��ܺuK>���<9c$`Z�"�/��{����[T�@0��}�����䆂�&���J���@VaU ��ЏK�̋/r�^���#%Á@`7�P%c�(	*�,	/Il�����\ P��tttqL���1�x������ft��ظ"Qa�����K �o�n8HVIh���[���V����ˌ\�� � � �Ap��T�&�$�q_ �6f�¶�q˘�������B ����pp�?�jGh���1a%��}�|��|��1�^(��q� ������,ԍN����eF.'mxc��N�7�n8�|B�"2-2�a���2+�$����do.������D*�H �H�-W(b�ю ��Ne�i���1���^�1��	|zz�σ ����7,S�be�^`.�Ҿ���V�O��ܞϧ�=���S	�h!�����o޼�� �Pp1�q�L\�ѲcY�B��`��8^�@ 7�� `�ަmT�������Lp���-�2-�٬����{�Z-��{ ���i������c[�=L�@Z1Ni�a�$WX�{���� ���~�Y���	}g����SԮڵKnw�nI.���]�=�MF�ؑ�	�)��r�g�_�Ap���� \'�e��n.n�q��`Ц7��p��
S]�I�V��R�M#o�B�	�\� ���~#n pÑH��N�ӳ���	�f`~م�d�l�[�X�� �o(NLd��t{VN�@Pa���c�&���0�ͳU�ܲЌ��aQ�Ap��+��[��o��k�$�el�E���'������&R{�F$Th�ֻ�#����>��"Vc$�6�X]�Ap��D~�~�?�.�Q`�����{YY�NB�&$Ł�7�g�}v��_�䔖�$px��I0ǸFC�2�9n ����p�V���;�:����y� 
$e�@�BY�SZ��Sv=�%��ǖ��ܸI��ݵ���D�@�����nAʎd$oS�HHH�Y��'����qvi�
.-5e��}��L;�y�߲`-�/��7%i�p��2j�\
.�JBO$n=e!XDཐ�YC�Ǥ*�u�5FATY�1��3���U/?�8^
n ������q�� �����P��O��(_tt��w���/>|���4&�$��Ikg�:q��q�񊱇qʉ�\�Y�1����� ����W��FpI`�<�����w7��DO����� ��w�����_� ��
�1��c�[� ��(2�Ap�=B��wcn�eL���jX�-� �o��-յ��fTi��ݦ��#E���P�.���~"�_ ��Hġ��[W53eW��B����䣌h�'��j	O�/��;�ٳgg_|���2& q%�����*��Jp�D�nL����~#n p��H�'�^��1H��.�Xa��oC�U�ۖ�V�˔�?���xg &,�ҳ�/�����Ҡ>ݶɄ㜏��B ����l@�J��C�� z	�-��7ښ�i�d[�3�k�t���?��˗/�y6|��{��~#n p����-�]�f�~G�0HwvIox���b҄1��4��H^��,�d.��C�@`��N��F���q����)	�
���2�Da6����G���T�����.zm9&K�7���a��n����Uν�e�ٹ@X��F�@�c��t�	-+�IJ����/RA뽗C�B�$"T����m�t�fE�z�(����Ǐ��t+�8�@`7��`�-�.n��N��m�z�;e�BYݎSTʂ���P_U(�%���$������8G�E��@`�7��(�ڲ-on��-"����y��n����ܲ���/Ъ�\9(�Gs��1V�e�����@ ����`0 Y(�
%	(�l�@�d�-R˦��� �z���'���1ö�DF�J.'V�G(����@ ����`��@���+�>�.P�7��߿������U/�ݥϛ��er�������E�@��DAsoӏ>	.1�o��R�%��ߑĖK��f��7�y��(�0�>�,�(�������~�X� ��@ n p�ABJQ*b��;�����v2{۱�4?�2����\9�x--
�$���ʀ�|.�/��7e�X�|Q	�s�����>Rme�z��'Xf�@�=Q��r��R��׶��D��c�-'�'��7T��B�����a�1�̶|�8�w<+�K���F`Qb����M��!�1��������2�@`�7��(#�X@�%�2G�,�!� rL� ���u��b<�S���@�Z�pyy�5�I.�In���[c�D7�/��7��1L$�&��R��E������tUqA<�25D���I	��ru�􁗖�]���&�]c�8n����{� ��������(d\�b�~�I	�:/#��B�[���h�|��G0��/�yL�q��(H��]���t:}���������Ap��U�J��@TIb��U���K�1�Uo�� �8�v]�re�WJ�L��[ƌ+g���6n ����P<{��/^��Ʋ@�j��ÈR!��hu���P��$���ҏ��{���6C����T�r���o�5�Ap��R�*q`S�m�K[ƄQ�-+��-�&([�"5d��$�$�e�خW`3�ҿ�Ap����������6���	nUW��@�������1'7n��BiA�B��Pv��=�e�2��ܖ��@`�7���%���`����^K�+����o�@NAjAtqvF��(`?�͢4�n�nf$���#��~"n pC��ٳ��/_>&Qx��,0{[3��:����7��+#�@TAnaW�:K/n��2�.ǂu�$7�$����~#n pC�~���3.�������
N��5*=�|�K�A �0��]�LF@�����G�3���$���f�l�a �h ����\t\��U��-��JҺU�V� l��!�M����Y�LL���p8��-[J�VW[��L�@ ���`�$h�Rm�~�2G����.	nY�C�Ky|SpҎ�qZ>��;(��p�.c� ܂�r�F�C��Ap�
�ASի��wW�e�:��Ą�8��Za��y��2A��0f��t2�Vzx����BS����C�@�����LP(;�1��K�����=&7�m��LK�Ĥ���Tqy�^e�-W( �o�8��F�@��b�����vF(C�D�Q���ݷ%.�f�r�@�4AhA\����2$,��/@�.m$�����D�@���˾[�e��c 
��2/�Lb����('O,f�$������6��\�>&a��~#n pCQܲx�$��6<����Z0\���[!�C��@c����LI ��Cc��$�,�,n#�@`/7��(-���.��e�Ӓ��e[��B���g�}v��ŋǘ`�s�,\�EW<���<���U����$��
���4ΟH �K�n(����ײ�:�^�{74��m0�������K�8����H��J����F�?� GV: ��Hd+'v�8v�����6������g�����ѣj�\km{�ӽ��^kΚ5k���Q�FyNP�۷��;��==�2���ؾ�㫣cU2��A�vK8}��e>fO���"�
C�0�7l-3�q��;�8����8�����"����������n۷���9}��ce���A�v�3�Ξ�a��,��v��q�e�7ވ�e���o���8����㐂���B�����ކ]�����ߎ�!����o�����xÍc�櫗��i����	��u����H�܎�#��g�%� /��%�D����g���>�۱2^}�՝w�y�KCl��rQ#��dU>�L���1Yz�o1T�;ާ_���{�BG��D'�G�X��͎<F�w7�)6|ק;����k��aH*i��}��Ѱ�B4B$�Z�&��ݐwgx�5:���8����㈀�龀���'��-~;:��R�b��y�Xrf�M#��x]ϡ�����8Z����"����`N�;����-R�VD���7�����7{�w"�z�i�::::���8�p�������%������Gm����"Q˭��1Z�8�ԓ!�!����K�����fl�K9sRvttNt���q�ᱴ�n�Ȳ�� ���[o���9sfy�/D�`@�Yh�ѱ��s��/�rV���;�x���"{Đ���;l���AJ�Nn;::�Np;:) �U�QbEl�]�$@Z��%A�ߘ.�܎M`��-7� �,2\� ����E�7�|������;yt��vtmt���qH��܊���q��<�aA�V��M�U��7vtl�CɣH�>{l7�ÈÕ���.,�*��[o�uq�m�-N�:5o���O5ttQt���q��S�S�i!L�jT�����\���m�[�vld吼��F�[ye�yK�n���7�t!�,6^}3���#�Np;:)<���9�E�|[���^",��gߦ��::օ��"_?�����o-~t��o�cd�ӊ�����G�9p;:�(:���8�`����ia<�lq
���i�����~;:J�늑5�K{�1N�xr9� ���w�k�bgė�:u��������YG��D'������λﾫ]��ۍ�XG�0��yq��%\�щm�&!�LApB�SK��AZ�c<$���n#͌C�ɬ���܎�C���;�Z�����u��E��ɏ�4r�����Ժ��)� ��<�܉���7�ɰ�r�s��}ߑ��㈢܎�Éq`=���H��Bj��e���߾/5��%<B�$�����Y�Bl�ȩ<�[��,7�tu�ulk>C�;ɪB�q�ܹG��vtB���^]��f"ˢO�=��8�WG�:x�7v^~���|�ͥ�U <F��Dn%��N���V{:1��܎���Np;:!|u�o�ˋ����7҂yNܘ���ut��ќ<yr���\Ȫ2*\�ru��gWX�I|���ێ��Np;:!|�'L@b��R��H!�ej$	�{۱A\��)L9��-̘Z�yi�;DW�IcG;�A���vtmt���q�`ܻ�4��`�A�i��W�2::��n���EX�U��=�u��8��ȭ�!���܎���>JutB�6�W._#��Z�d������$��3�B'���M�/���0�������eHr��7]��B�������R��豵loJ���r�KYNx;���<N���U�/���ܰ����	� "��ێ��>JutBh�W�AdV�x�D"DN�:�̞�V��j�������ݎ�u�e,
��!A��wɱ��ʓ{��^�Y���/.���:���8� <��bm���"�"�ϟ�#s�$/kk /�V��"�`��qio�{}��Ɲ���܎���Np;:!D`=q~\���ۨE<�<c�J LNt;:V��X\ 	y%t�C���e�_fvуq;:�(:���8��B2�z�
Q`x$����'2  ��ۡvt���<�G�\�~�gP ��_�����.:::�$:���8��K+8y��J�Q�i!L;��E?Lwt�ȭ���o\�<yr|���E1f#d�I5CA���s���ἳ�>��EGGǑD'�������<��i_��z8�Ʌ�+�;�P�Y:�r%y�,�%��;��oɳdQ��;�"4��y���EGGǑE�::! �L�B^EȜ �i ��1ziz�ݥ�E�K���cm��7)��3�0Ɛ[N�̐���8������ �eQ�An�HpE�I+&¡2N^>9�>���p�k` �K#��e�JF��NW߳E/���,�Nn;::�Np;:! ����Ā�[��N ��?��K��@^�����q�p�HF��;�B�7��
,<C�c~܎����Np;:)���LYv$�K�F�#&8Y��̞�����EGǊ������?�÷yډ�l[��;�,Cd|�i2�O�o���Ȏ����Np;:!Xd&�h���I�!�,�9�}b�-J�;����ϙyq{"܎���o�����x��7��`��彍|id�	�o��	nG��F'����Bx��<b{�޲:ݿt.��P��M` �Or���̒����KK�ypc,���`���!t���q�������W�zZ^\M�
�KY�q˻�Ŵ��.���ǎ�U1��e��u����1�dS;�uttt�����A��'N�q���*g�b}���mz}J�����l��I�.)錢c-�<�.��@�x]��༎���Np;:�zY�<��!��
L���^�1hU� ����9��_tt��ƺ,
d �S�ŭ�1�����vttt���q���'���z������?�Y�����������?��j�F��Z��	nS�C�g=nGGG'���/�� �'�����
u'���q��c[K1���W^y�ܽ���In��pb;��.����r�-�Kq�鱡'��#�����܎�C�W����t�Ҙ&L 3����Ap����;*�8+1���v�۱2bZ/H����ɓ��.�����-�*�fG��vt2�HlI��eI���(��"@( ʜ�����V��"���gy_e��,�ŀ/cl=�-�B'���r� l�/�(�[�Bu��	\����;�cp;�E-NVr�<��b�n���l7^<��hq1ZGG��E'���������矎7�@'Q���"���)^��>5��1�K�;�2)9�,�c�0��%Lf���r��\,�ϙKV������Np;:�����m��P�|�����nY�C�p�&!2����۞\A�	�O�}���ͻF$}a��yGG��F'�����'\���̲�S�=�;�c��
�ށlt�б6 ��)yoEro���}6�6Ѿ}4�
��;��!�݋��q��	nG�!B�A���f��l���k���ɓ�x����y��/::Vr&B*���lq�^]��f�X�[��
w�䶣��܎�C<����
s�(�Y�馛�v�
a
q�����/��ߎ�@2%���YȤ�U�CZ}���8#�������8������/�l/�yȈ[�T��ӧ�1�������b�;������k@�U/�"�9$�ȞdT�q��q� �=D����܎�Cz߸�I���{�8��
�r��;=�B�� vV�V�U�
,2��\f<�s̚@��@r;::�.:���8D�T`����'A����
B��lwa�r�O�ֱ	 c"�\��[�Bp��gxgG��ty��Nǹ�y���8�����!��Bb�[�g�v�bz��G�b���Mwt�
�e�bv���3��e�̕�˝����2���qt�	nG�!aNN�K�%��Ҵ0���H�F9�k�qP ��	�2~|�8�kK&��	Ƕ�-�O�Kv�y���Ȏ����Np;: xp�e�ݝ� �������	�0)N�M!:q�8h F�����Y�K��m�a������8�����b�0���O-!
"�丅Ă���=���s4;Y���` �}o�ɽ|-|��[o���iG�G'�����rKӫ�V��K�U�"
�~�w�:�ܵ,n��4Bz�B�&�q��Β�N2���E��}�c���E�=N����܎�C����ص�l�IA�������ˠ�"��':��� ��]8���y��a�Ab%�o�����M'oZf^@Y�F|9�:::�6:���8dȦfI��w��\�t�����^#Y����������X,t��L� �Tt�͐Ia$×..CX�F���;�utt��vt"������"�w�{wIz=9>/�b���O�vl�����8�-�+�+,�Kf%��}���
��Y���	nG��F'���;���)�߂�\���^���ܘ���cS D����	�~��;�ˉ�wWǰ�o�y���8��������g�pE ,�qr���wtl�%S�s�5��[�� �����p���}'���vt"0���I��žmN����#7�D��ܾȬcS@�DXo��1w-�H� ��[�`������V��vC���h�܎�C��	��+��0V���B��4���,�(߳���P���)�����s�\a#���
�qd�@:::�.:���8D��c��ֱ}aHӽ��/BX`�sn�馑 wtlȕ��^�Gf�dD2'��3<�xy9�F�;::�.:���8D����'�-�!�<^��S&B!��)��ܲ���x�[����u������E�����	�]}ֻ~�l��K:::�6:���8$x���w~���?�A%ؾ6����q�٥�ץcE;��x{c�m_�ӱ)xHA/��v�cG>Bl<F|����b�X���8�����` �Oooo�x�S�"\�~����0�w�5�)�:
#���E�8���S[��a�嶣��܎�C���^�T_��/_����B��!�8\B�6�o��q(�Do���S�yo���l�x��j�َ�#�Np;:	JS��  ��q�"�"��!��ѱ.|s�,��/&�g�,�E�Y�2`�����h�܎�C����/��:z�[�F��3<���c�m�B9�<�fb��B�{����Np;:	��ƘZ*yGG�{q?�uB�q��+�.����#�������>����Ep����q��	nG�!S��I�mN� h�'����l	Ƿ�-�q�-i�������.::ք�E`�I����I����~=����h�܎�Cyl��R�0�ٸJ��zE�����˭N��Bxuq�������{n�ѱ&�1n��V�"����
�)2�2Ho��::::���8$%%�ӄ��P����._�._skް�`�c��GFNW�s_,���fq�G��vt8�e��{�^�0v�"=�ǘ݈>�۱)d2vu����uy%�+���Ov���q��	nG�!�щ�s�.�-C|\�+�"o�����t>1������Ӌ��M������0x|����i���d�8]�:������܎�C�S�q�<�BI���*\��F�qqo�3/Ϙ^*��c�9�\a�	xf��Ev��w�'ױ�۾9IGGG'��q�^H�ow��DlY�C<�v6�T1$���\��c]��]䡽�[W._Y�{���#w���J~��r������Xt���qh�����]���;��v��f��$����8��w��j���o^|������K��,�`�e�7�l!e����q��	nG�!�0�_a�� b*"�ߊ�e;^BD$D���i,�1tn�F0��(KĀ��3�,l���4{~g��d\xv|o�2�e??���G#�}��W�|뭷���������^�F���:;>�E���}kƩ�j�W��R=k��m,Al�R��]�����a�����[��ٽn��)�[n�����WE��}�W����E
�~���%� ��^:�<,≹Hi;�>+�q _������V��Bܥ�tL�޵�]4u�_�//��fr�}ߊZ�^���<��L��?�>B�q�xZ��a��^y��7�.C�cb~[�E��%��SH�Xg��ruY��|ϗO�>��������Ud�bd��J݄̭�'�Λ��U�7w�.����U�_q��Z�-���mE��ˮ�	�Ye�/q�u�ϫUJ���|?>��F��������������7c��;�r3S�S���p���d��E|؋��5qT	n�rj!���u�(�w9]�ne�S�䁾΢3V��P���_�Z��{��c�)��o΀�� 	nVn$s����U���ӎF�T��}^����zk��o,N�:����X2"Đ�N�;�1ȯH�/F;��S�!�1�\6�\�����MrW%����;~�ʯ�_���:�S�A��5�q}�����u[ϛ�K�gju�\_�	���������~��Q�`�����\6xD_�S恩��a>P��h"�+��ޗ�@T��*ؔ����uJ�N,��w������]�����"�gΜY<���c �z����Ř�{'�ͯ^
ux��/��b:��i�<?��2M�Y���z�r[�A�܌�����E#�^�á&��M�%c��[�xm'��1w↥1&����YP���//���?�^h�Ȯ�Λ��o'�m����:���u�_�k��{��;㘞�3��8Ʈ�M�+�-򟒼em ���[n�<�_��W^ye��`IpIO!mQ�*�}����?n��:���jA˱�*���������S�OMp�@� 廐�?�z뭋������}��\�\�	�''.�r��;��B�	�bsg!3t��Z���7%/�<����g׬S�~SXǫ5u_%���7���?�x���� YDJeTIn}L�1�iO�U�An���� �����X���Kcz�;�S�?�u�7wZd�k���bk����+���a�6���T��_+�-�bU��[M�N�q`���ђ>�x�,,#�E���E0��;^�V�Un��88U�m"���4U~�VT`�6-��=`��9��l��PSnS^�V���ј�t"Z�d/�m��6��8E�_rr�ҟ��B�����g'���?�q���n�,r���ڽM=_��c[Ik�\`9.��*F�A��98Hcu���n��[4�d0Ie�y�"��G�9}V�#�|i�΅wƐC$��o[]G�:_�Jh�:�	�}��YE�@�Z�/S$�V��0e�O��!�^�X^ú���V%�S��{o5�Kרq�x�X�XN��%]��܌����[��e�)���?� ⓰��[	n�[~���8Uv�`��u��i�ց&b�mB�RF+*)x?f|�rk
��k疞-Z.�%� ������-y���A�3����Q���{��˾�Rx�������m1pKV6s�I�1�m��VxKSv<&�{\,V�e߹��A�4�Aʷ���Βy}G\}����Yֵ��B�[d��9cWv�-2:����T*;��V���5W�[�ɺ�r�j%dܣ�g��=l҈���������i˖�Z"���S�6^���E�e�C_ŚUb���Xa�k2GVUl-�� S׮4�/	��Ar7q^&�S�k˳n!8��砅���K�Z�O��9!p䀘U�0�۷@]zn/�y�(ӧp�*�;^:����*��*
j�~p�Ϗy$	Y{�{��T9j���v\Dk�9.�-�tQ����d��#��;vCm��^��$�ġ�8�by}ٝ�e�_�H�6MpK��Qv����Z���zO��5"R#F��KO��ʎ�^sQӻ5���]�����{7�=�t񙖌�R�L��)��Rr0�ʈ��/	��e!�v$�V�V+��a[ʚ*��U��?ȹ��}�X��J���1U�g2u�܁-32Z�W*+��������~�0��n���D  A1��su|��,�W�w��X�x/�����1S���ܨj�ر�rnAM?�ͬ�c�����N�#�D6%�:�Cd��􃋋�[c��Qv��H��o�!
.7�'�����G�8����>�YlҠ)�u�5Vu� �S�%�׌2�ں��Ι��xCk�q��ʜ;&��[볨�﬎Q���gi���,�){���5 �:��2����X���_+����AM��Q|���A���O�^�|�͞�*���cK��]�m�5�罌�t����U���9gK�:�~=���b��'t<fܖ�����qW����dbйx�j�ƿϦ���{��F�#�"�+/��ϙC�c��:��b=Z�Cm��"�������賏9���^c���k���c��q�H�2	Yؾ�.�ǀ���W�)�c�x�Vѥ-zk
s��2J�j��"���5�us�ϣ66��_�[�(��K��t�%}���xLVNl��}L���v��I6.��1����zAY��������q�e������Z�em�	�*ʏ� �k�s���;�Q��ux�[�o�Ϊ�C�Zˋ��ӄv��+ʉs$>Q2_�+�Y�\��t�~�E�L1ƶ��nb뿭�JFcKx�:�\��lBֲ�3�%���O�l�qa0�.�v�u=�,q��X�m�eg��ﭨ�ܖ2[�A�}�d?>��1����yS��T�)�u��o���B�]\F[p\�D��Sj����utd�qW"��:�b9�����U���$� �b!�TM�W�V�o�j���[��+���h ��E�Z��*�s~VO>KA�>Iq�z�WB@Ȃ�%���e
�$ǥ��2�⹥�n%�5����u��+l��-���^�9�V�i�2:��qa{{�[bˑK���s҄����q��S��2=T�G-�ɍ׬��.5���nK���*z5֡�{�>�>-��01Վ��'�s�k�'��^��x�1�+���)x�j�o�X�%DA�s����U��\"R;o�U�r�M*�����NK��'��ͪ��;q��&E��H%B+b�Ͼ0�C��]�|ײ�=qEX"�.�~�T۵7E�"�!r�u�>���U�����W.�A�D^2"枰�3��2vw#eϳ��]�QP�4x9q�!^k���~ϰ	�*GS��fp�r�s�ƨL�[���k���\"���/]w����/?��~6y_%�mèT�}i�Z+���]E	�f�X`dVfힳ���d�u�>�1N>J�y$֕�)��B��"��=��� O�0�Ȕ�cQ�+� �(� Y�bI��}fD�48��{�9J���J�שêFqv��<���������񒹷�~{i�������g���~�ZJu�oJ������A�]�k���P��A8��H^K�����Z�M�O+65vN�Z�־�s�)B[kߖ�	�B|��R\�@�A�n���Ʃy
q����B�)㱵�<%$5K8+/�SV���s<-|��S��yJ�J^J��E�d
Z/��� $-��f�wqu������O)V�^v�x_���d�VF,g��fK���7�Ĕ.(}��V��u-ʨէ�$������[J3+�1�^'�-ׯ-�*jcB�)�AF��y�t�_3��taVVv-�K��j�f�)W#�S�Y��5�5lW�Z�9s���Hˎ��x/-mq�w���yx�6��n�̌��`F���1Z�qn����k��F|/]�2�HK�����6@���ܱ�u�h��^�]Z�#��v8�M"�J������������)�(����*h�S���R���*�g$����k1*K�q���bil��,J��R�:Z�=�:���!�:>��W��uƓV�^�����A�<��^v_��߲���ݲ������R"�N03Yly�n�L�{V�)P���a9k��ʭ-e���A��3��W�>n�sFv�R�~~+��*��[�A3B�ΰ��ρw<�M���q�r�~nd��WTH�מּ�{�u�r[:a&�5ci�8EZ�5G���*F�{YEV���E
�%�=r�߆���%���dJ�LI&��,SJ��*+��֔f�}�Z;f���ch'��&���1�����d%"3�DBP5��Xo҄I&F�<��g��{�Z,�[�[��x�ƥ�wNH2Af�Z���E�V�S����Y���UIҦ�|fHŅ�|.�9���d6n���3!,��M�^�کd�d�m�Ɍƨ[k���y��ѲsjKK��k͑�lL K.�S��E��k�V�9/���]���J�TB��:̔���r]W�-q��S�O�������[�����\���jr<W��:�x&2��ǣ��ψ����/���n
�@ ?�����l%#-F]v��I�������\yh틵��>3�P+�۳6�e�#WĈ�{����d"���S�N�/�V\b�EV��AFy���>�|�X�r��+��xnԱY����&���3B���3d�r��O�I9%]�=n�L�1�
��?�@��S��nt�kg���0��V���nY�2������K����k��Jd"k�����Luʃ .5��+e�2c�4`�#�J�搘�^��J�i)�4����ZG�)�x�A�HK�[t}޷��K �v����[��Y�O-
&��fi\�ؖg���GY\W'�R���ߟ_����<(�Ck�7�V����V�b̻��㜬�^^'63�a-�J�O�x���ڕ����?J}���W	wYC���D]ǛH[�e�:���$�T�Y���5Ԟ_V�W�^^�:-��{,�1Eҽ%�Z��>ni���Q�fb�K�TN�P�k�~/��&�b{���-��{m@�zF��R�x�J�6S�~S�k�}��Ĕ��(<�uТ ڌ8ZH.Ӿz��w�Њ�f���}��O����?��B�k�Ҫd-����������,��b_l�_�Vb]k��0�Ώ�ݗ�񻫋�n4��x�Z]j����m��������P���y�ԙsxQ�[�_�n�Fo:����xMY�������n���#��j�f�T�6;(�Hc�9-������m�R����k�-i\�BVQ�-�����5��[���ʇA����s�j�~+@~n�1�IT�5AA����G���gn'��aAk-/�&yM�j�W�5��ߵЌx�lש}8�w�l��z��-����{�[��D`�>"�)^�T�.�c�>1L��[8��LO�{�{(�M6@�с�:��r$"����m��[��ϖ����sAn(��B9�Zߞҿ�L�玉-��s�E��u�����;���r�Uq�r~cqa|�N�����a���]}S���D�7�Fv���d�|U�i���P&�S��"3s���rK�b�6��̚�
����^;?
�L�U��j�-K���5�P�z#Q�)���9��y��-�80�ܛ���=q{$#�ar؄�eEm�ς��ߊi$fQ�ɻ˖�<�Z}������D㥤�����ʚ�oJ$���.��yg�����,��=\q{��e�Ό��s3��Z���u��c<�B|�޶�h^f1/o4�{�ϱ[�;;nJw��W|�%R��I��c"���������'��%rtc�Hޙ��z8��B�|�P��>zy;�+��D��W22b{��WZQ��X/����vv���-�l�~Z�y'���>ETce��l�4[;�r>G���RɎ�<WYys��b���׭sV0k��+��W�����t�3�ih���,�����X�^s� >�U;o,��*�s|M�c�Q;�,�(�������  ��IDAT{8��/r�_|eӂ��3R�ow��3Ѣ�KP���J����ey��3`˫�l^�H�K�#g�ܿ��6��\0:�_c}�.z��� &�{j�a��]�'~���k|f�=��x��V{f���oQ�J}"��x}�G�����F\��ܨ�jFe��}݁�;1z�9�uA�$${~^�,�*{���-�sZ��dϨd ��U�(-�)�K��S����9�_�^4�i���N�C��)���.�J�#��B�,�	/)))&H/,�1��b���ڿр��A�D� ��H ��}���������M��Xv�9ך��(W\ߙϠ���/������+W�p��bhJ�\�/ef��}`�8E�q������ൿ3R�ɕ˳�J�=;�����V�2�x�|Ҷ��)L��(;��g:�Q���c{�{~����D�1��	��E��3�2U��9����9���x�Q�� d�>�[n\F�����`�ĕ���$��6�r���ł>��m�ݣ��;��%o���k�4�E����N%��s|��S��{/3K5��dH��i�9SN�T�GpK�z�x�Xf��V�Bټ�N�Mig唂�7�c�4;G=��j����oV�+�(�nM�v�mcnJȭ+4�A\���!N�3 �� ��,��ֱxxE�'�,�|�R��)��F�}��Z.�^F��7'��."Q�>1}ǖ�xw	YF��ա�/]\��޻��n%�������!��H��-�:�Y��������)Y�Z��?7��U���~�=�,x����w�=�w�qjo������~���/~���D�:e�J��F���S�]�ܲk������r�!�-$��.x[�G��1���I�70�OL������d���瀺L����ˌ4�w�����y:A�ލռ0����[�_��z��^O�o̝M�=VW�>����vn7U�?��g�<�y�#����8Tҥ~�g���Z���fm��:!k���d��qGoaIp��>�R�K�ծ3Uv�k�^� ���f�[��:*�L�� y{B�4(c�K9��;b�<~3*D��ɨ���"D�/��Gu��[o��8��2�{��l��B���9q.u�8�O!�S�y3��-dJ��~W��s�-�����c���J�)�G͛���)y��m|�*y�by%"P:������0S�S�Z<��#����.Ƈ���&b�g�g�ꫯ.�]��ֈ{MƐ�sI7e�ϋ���8��B���=y�Y_�	Y���1���b�>�{���R9^׈�����k��Q��<�b��x�U���ܢO|���Ջ�BgQ|!+�؝'���6��r!˪��3����}o����;��˭˭}#q.�Z���Ȍ��Hfh�t~L�K�%�V�S�s�������P͢0�Zce��3��V��P�eQk�Z�k��&���2��+�өkGE��:�^R(�ӧO/I�O��B�=����;&
*n��e���c�:2�+R ��OQ�9\s�8��<�r����<�91�����QfmJI�x�Y?�z�ȼ�*�	��}�/)�~2�'O9^����|�+��~���;�c��8i��O|��������O��������>��)���5[�:5h��!#a���q��Y�Wݷ{g��Q;�v�B���ov�n�oJ/�W�]_d�?g����c����	�i<P�{<�~��zA�=U�����d�l��sFG���@�	u��,f��b�������n�"�u�E������3�Yۯ��1��p�~�}�ƥZe�f���l-;�[F���>�Kn#���֛��**j��˼�� �)VPRd���C<ǉ�����C*%  ��Ƴ�_��\�ʊ����`�N�&�S��8+MEɫ��b�׹�XCk9ɍ�����)����+�?�ѳ{5�z�u,�V�Թ������Z<ǽT���2��#m��J�;��{ｋ/�ˋ���_.���/��/�yzW#.�~����G?`?~�>Qw���y��eiN��w���
�C���7j��=P��$[-3%�5j�����F�\d}�������2�R#ټr���»�c,�Ɗ�3��x|��������!^��]��e��oxe��%�p_p(�$a�'anzi6P�n��z����Ug��u�[	%.�2źgcoK���+镬�UxN��ؿ�i�j��Bi��*P��Rg�R�뒖x�u�?~�n}@$1�rt��I���:��3gFEFH��(�\�XX����������u=����g��c���K�"�+��9_K1��ҳ.��S
r�b�����hx�}�
�������;�/"�6w�?U��{$��v��&���.�E�zN)^���.����${�O�܊�>��C�ߪ�x��A}���?�4&�6��O~����\ǌ$Y��z�~�Ϣ�Z[�!r�9�t�\�)��=&�I���\�гx������d�e��ư�>� ^?�]%������rL��a�}�{B�����!�^�}�k˻Jߠ\�yV�g�`k��z�уLJD�W��Q���q��7�|�`��Y�g��x_��R?o�/3:���u�ob��#rB�>n�d�撼X�7�܎[S������9D�t~V���1�wi`ά���@),y�n����ͷ�<*2r�
[���\�J�8������q\�%�Y�M��=1]�$�@X��FQ�����҂�s+=����t�Zb�/�i� ��"g|�W�S�euʌ��vh�s'�%��1�S�\?/��ڵ��e2B��_����c��w޹����x�3�,N�>5[�#I�_�;���oR���+�7�|s_���K$����E"�
6�[i�R��RB�._�3���Kc��]�b�?��9�F��7Y�V]ñ�@U/�͈�a,�8�uv4�0�x>~���p㈎ոDH����,�����#t}����g�ո��ɵ����D]����fz%�����3͌���LWO��ҹ�����O-ǔ���>�����lsP�o�H� d�꺊5|�^�&BZzs-�쁖�Y��{\X������Q��Sw,n<ym:�r��QV�Du+*POV�bbqַ�qQ^�a�Cq��D?'�s�����R̚���dc�$��4g����+�Mb;��]s�[aW�i�H�}!G��5B꿯k���F2��]` ��k��|p��C-����l$��[DWe�x�{��S�zV�M2��c�-	�H�K/���r����c�A���ԏ�|S�jqܸ��n�ڋ�S�x��.1��u�(�� �%@��P;�Q�#�^�=��G�pBe��Bn�{�m|mۅ��p]�A�k��R7�fܽ��\�1�\�4B�Xl�39����WY��.�aH:A����U�Ci,Ȏ��y�\���I��J��Ǵ�e����|�k�����<~�V%���U��,��͉��$�i���?��ɏ!�U�]
�p�*Ҕ��S�����wȭ���t^>�8�ձ��E���Z����Ԕ��O�	�&^f՝�d��V��!#LY��o񺙡S�f�82'�7+-c��nq<g�⢊x_��5�܏�2�琨ɝ"��>8�I��c8�s��c,&�%fP�,r��:1�>�{L<F����(M�|}/���I���9z9��([��Uɡ�����b�냫Bj|��	���J�Z�f\kS:!�ەk�:cJ}}����Y$�ҥ"�
�2������|��R�u���f�˵?��"������e<�8�1Nw�~ǥq�S�Չ=�����aQ������w�|�PzV�\�:	K�G��T��q�O���'�=3��u[�CM�d�ಜb/��Ջq&�`T4���򀻤���˿�qB���HK���)=�߽,����w~�bҹ��j�W�E(�AX�4,�C�8��I�,�<�(9A�x�u��ul|�x�|����i`)=@DOɿ}ӈ,&�e���HINP&S�gi ��<��3f����L��w��M��h��齁_�M�Dĭ�������=�J.2��T_������$�Y�"r�Є?��?_<����v"�VmK��{c;���w��Y��~��/^��}F�S�[{n%X�=k�H�b]�j��͋����Q��rmQ��5d�˭��G��*����;{/U|�Hw�~n��K&5�'9�(�x���Q�#<<ġg�s�zG���~B�A8�L�oKc&��}��q=���c�,IWB^E�ɾ�쨎d<�q���8Oa�����gk�!>g�˞��o���u��~<7++�ya�o�8K�l��k��҃�v�R u� �Y�o���T����:�����+������C����.��R`&��� ���ņ�R��dO��b�i'O �9N*���1Hy��+��u�l�� x ��BaIY�띙�DE3�`e�Wpr����9U'D��A�B���8F�ډ����� ����	��1,�/�t�;�,��*�����E�=�Sm�6W�}��7fIP���Y�%�!y@1��le�ǈ#�*[`�V�V���t,us=�Bfk��2��p���$�T��b_;�BI��b������i��S���wOj�]�K{}JcP��{oOB�d�����V���3y�p�4��p��	����3q�e����� ��u��x �`L��ꟐV��s���cFܼ��Kߋ��3En���������V��2Q#��:��Z������fQK����c����ۚ%1%��)����3�W+/"��m0E`K;�L���[Vu�$|�s�p��P�.�#���Nt]��g�kR�@|���>J+����m�!�>х<c�볔�^�8.n�����$"i�Y�s@;B��y�{�e���r�>�*�Y���;��<��1�i�����_id���~��D�~�]w�ƅ�-+��y[8��Ȑ�#qz~*_q��Nh׳7�xc�G��Pl���)��|V��1�������/���N�_�7[�_�8Ab��ˈ�'ȥ��d�=��d�!������X���238QE�z�a��Š��p��P�Gc ܸ.�нs��p���܇^x�!���B�kϱFH}J�_-<�E_N3W�#I�t=��9S�m�:g׊�#�v�:n��K��b)������W@��9��֩������\2�:����XQ�[ud<��i��WFr{�Kk֧`O��AI"�(OC����B�E��,>_����W}�[K�-bLV,y��}�د��6�(o�]N����X�G]�^�%#�S}#�c�wT�>��9Ȧ��)�<���h����*�]�?���w��<�X��s1�}����&\�=OB���#���jEI�|�������)��EL�o4��	_��l
����k9�T/�9��������"���B���ɘ��xU2#d��~N�~����;f�����3�/��C�;$��,��"$�vȔ@8$��Ce����_���,#i�璑�Uen� {}VE�3b8's���if���R���~�"�Z��&]�cG޴��J����+���u-��/)��|?>�Bbٙ��S�"�Rb$D'�I����;���vQ���б=�����e�^X��CvH]���s_�%����$��7�ӻ3���0(n/GeKz�'���skߚL���Q�x�����d�fHf
:�k�}6�:��!����ʔ𔒜��>]*ِ1%ȓ#o�r�*ޖ�$�57|��zy�O$T����V��п�����$�.�v����ȑ z�fXE�K:qIr��O��c�]!b^��͐L�U�%kG��f �ޒ��6���r}\Pۈ�I��b�8O�F.���2�9�]�����m>��T`�|�����L-:b�=e��X��c��=qq#T^w��N���8��k�J�Ǭe���HW�:�+�Lo�"�S}:ʥ�U�[�o�>�1�\��#�)��l�8�F�����Anc�~�lI���� "j�~�zʎo�XJ^I�"8(16o���NK�'^�+uZ\��&F5��2MY�@���e0��<Q ^P�@��<.ѷc�>Q��S�xi�@b�=�= Ѵ\ �K��,s��b�ܬ���賓x��D0N<ϴ�8������������z������n-�x[f	�����?0�%hQ�B<�Ǎ���)3��![��Ŕ���g�;7�:L-����K���*@MJ��$��uJ䔗��L�,��_/�ol�O����4Er�瓕c�K�x2=,����O��V�j��#Ɩ��j3�?�Sَ��£�y'���y�/xA������7ό��.2�m��p�g,0��m�Äxa^d6A&��(�����W�}%���B��JeM���<վ�e�X�N��S$7���{��\�U�_4+�t̺�b
S�LX2oFD�`�9� �!�d��!.�i�(�"�t\�;�gQ�;�{b��o�;ʉ-~=7��J�nUc�S/�+H�2J�'o-d�).��	�vW�
k����D�ሟ�A�h�X����;�?�Ue<3�]ɕ�@f���K�'��0���X�<��"<��G_��<�������o�n\�����+kC>3�"ϛ�Y�T�VוwY^\�N_���wq@��Q��0�)��L'g|&k�q�W�׎�;��Kw�qAK��
2=�UezUx8�����w�"�g�|��<��'dU�Xd?�4b*�w#��d�v�g����<[w̨^��t�;�Eft>�>^�>dE�s�1��WK�E�����yֱ/��66�1�3��u�n�p<D$^����̒��}-��,��9��[�2%��/�<ώ��4�fe��v/�߲zg�N��Z�:O�÷��y2����x>}��:5����D�05�ט���H�}�a:o1�WM�Xe�N\(f(�R�-��z�]�P����u����Jp��q!#���_�6�l(<Cϡ�����e���u3�>�6��z����)=�
dA2���9UnZyo� ��׍��	wFRR�B�O<'v\z���!526��_.g2b�z$�^~M���|f�D�&�K���>�-�!.�ջ��/�螌p��Ϲ1�5��mP#�r�m�o�ڟ2�K�%�y��k�s��ƽ6���=�ﾷ����NddG� 2��X��	{�<�v�y�,3.1���0tt����C�<���)��2�=�_٦��Q?t�2���e2�uf$����wO�2J���m<'�6���>5��q�L�d�MGA�$��ja�Y��s��e�tL)�M �dߗ�#S������#�A� �ģ��s��G3`�ҙ����Ӊ��K�2ȍ� ����
X�#g.�4p}�2�Dݾ���H�M@�vAzO�$0}'��|/��&�\ce.<;#xCx��w�8��&���F���	3��r�"��%0#�%"N���J����s�$���~�k_7r���vd�W�;�Ż�q�L�:��x�e��^>���mxu��������/�WW}�8s��x����v�Ȉ��-��ǻl���$?����u�2nŷ�(@�b��$GR���Zߎ�`7j���嵎m^n� �ȁ@�K�Ǒ�3d����ǐG]���؋\���F���NU���t�t6���T!f�I���gO����B`}�����pg&È�F��^�	�[�@�)��G9���<��[<.���6�^"�Il�ј�r���d��x�,+#�Q��2�HpYY���h�|l�����[	�_RHY}J�[�g�^-D;�H ��?v��(�,h�-�.Uǲ��W��]�ۧ걠Q8:2Jgv�Kl�Ok�x\i@� Ӿɀ�W�U?)Cr""�C]"�G9�����>J�վN�ݲ�U� ��-)�U�>����O��1$^7$|`s2�툖�^�컩�keez�֧�~Tk{~�yC\��������>��q0c��d�V�i�୿����^[n�~'����)/���u��$4���67�\\�tq����_���˸K���,k'�{*,,��V�>�I���X�T����Z\O.]w����*�/��g��=��r\#��{�ՙ�16��ս�G����}�t����A\��~s|{_b��pd]��x֪�dv�H<7\��p��nyW�c��w�k�9"��lF�+��E]�1�̽�ԑ�`�x$P�s��m#�����5c՟o|�%>R�Kq�0s�֣S����~�$�T���J}�cK�|;V�6M�5��]̽V��R�-���h�����_�䝘��=�����E@:.ܽ)��K����a �SK!�;��<Y�ǀ���50K1�*����)�HF\P�g�>�+�"R�Y����q1U���Dm���|�>A�hѾ?�qs?��TdQ��K�}Ji�rK�j��r�*$A^R�T��}@����{a d��z�W?�������(��E��%�;�FH�n�;��{������u��U_�Ϣ3���u@��dm[2ޅZr<dO�@���e*���d���LfϮDF�{��/N�7{���`,������5����Ƿ��e��uiof��[��ݿ=��/T��7}boٍ]?7|��`ܽ��4��q��ø��` ����l�
���dD���l"���{�m�Wx`ݘ� C�}pg�����9�`gz">ù����}|oՓY_mѳ^�x���y�kԈ��^�¶�Z�܇���G��j
�E9ε��
��]:;�c�a��W�:yqR��#���]l����"��4+ԋ����4���Y^2]C�o~�,�6c�c5���s FA�ث^�XR}� K=b�cW!2/���SϳE�<�2#�x�d�I�@������d}n���lQU�\W�ęGr��y{j7�LɻH�<�"�����s[#��Er�������9�^"�"�:G�R�r�"&��g#)�#]�3��(#�z�����%��ߤX���)���9rԵ����]"���t2����Y�9�7��NK\��:��m�����p���ѫ=����Ó|M�2x\+c�\Bܩ���E�9���Hn��s�۹���Af���������>�����Z�����9����)t%ceL�Ƣ6������N[e<�x�;��8b��!�-��tE��U�K�����Ld7R�K��(!>��:��0k]t����P$�tX^]��BƳ*���%�MO�M��ƒ��Q�H���ӷ�^�v�m」Jp���g;ĨNԅ�X�x\!"�����C��ź��V9���C�uMyv/~pq�jp>��By��u<���׬Ϛ������t�l,���{BAJJ�e�m�:��d�F8�9y�p��lj!�[axg�0ʈ�+<D�^a	?��ǜ�"��(HE�����:O�N��Tf5���]u&ސ�:�3u�����r�qnTԞ�_+R��i��({fB$�q��Nߘ��}<��_7�$�.�����{��ۀ�Z�D��z�������Y��hy���xMtG����x(���8I�"��{o�������w��y���_�C�gϜ9���g�dz�� �<R:q��iFp遶l�G���?s�w��g�]���Ŏ���-�c6����=���`k�q�U\����o��1���e:1�G3�-Y�;p���
�<ع�/=���5a�]�X4���"f��O'~x= 9()���,����ۊg���O~��x&�I6WP:�����XX o���@-E���{,xBPd��ж޾���=a��J���֟�?�ճ���w�Il!�-��=�``�a� 
�w���*u�
,�%?��.*�h�Ĳ��c|&C�9ڿ���X|��_?�VI2���`�}�dI�R����s����d�_�j<��g�@K�$3&Nb��}��L�M1���Mb͌�m���������F���^Ƕ�}���φ�2����i����ӂ(���l�ˈ$�%�	g�	Ļ2���I�'C�]�/�أ,_`�w��9	�N�|��n^�'���c��?�[,�����w������tq(���;�VB2/rI؛���5]K��lbm��FO7�j'ʄqѶ�KRO���h,��ŉ����v�|K�5�'��l!���ή�]+3����sc�:6�)�=­�,?.~�M)�Z=j�׼��VJ��Z�����q�ɽ����{Z�q��Y $�C\�D�=�
hk)��I��.����Jǋ0���;�_�)G�d�^Aϣ�g��uo$����9z@�o�����(6�f�:h|�SV�7�E�����=7�+[_icĦ�+?��j��S"	(��T=�ZT��=���Ua	V�٠lod�l!"�����������Ǚ�xp������/��^�4h	�2u����1�$��J�������3�q+��2j��x\$�"�s�wR⤁�J��"�@���ˌ�2%�Yy^�Ͻ
�7K��w�s�)�o�.ɠX��l�rp�L��׍��ł.7��]v�D��;��ߟ�}v��{��׻������,���9O׻�7w8����p���En����
'�O,�>�~�r��0���P���,
��#_������mM��*�Fzv�Rߞ��m���˿��q��f�(�4,(5��8�X���S�+��K�F������W{��}� �B��鴔G���^^���+f��5�ϖ�"�(::8� , ��X�Y�@��J��{��������{� ��E��!�<)}R�~��-�2/K��)9)�&�I�k�WP��;�8Qs����ed{��ʋ�^#��u�X2�8p�$hQ���5�c�ީ���fd���*A[yo��ߍƛ��������!yZ_|��e���6��YF�obB��w���V��\DB�)��ˉ���H&�=kM�/��WB���,NЉ�>�Z䄲T�M�E,{Y���b�8��BlJe��9�q�L�\n��H�.�ã.\\߇ѯ���|X#��E�߿;Fiq��ᵵKp�pv�Kb�a�����O��P�H��>W�z�YH���ƍ�N޴`aݻ�Ǫ�^X����>���>*�Th8Ohw'�5DC�DJ#[�(�l�p���b=k|n���1sU��cp[1�SU�M��bMdǖ��oKCr�+^oJ`2�vA ��O�x�;�,J�W|��X�z�#k��"�9�e�(C���*�������L�CN^�"Ȫ�j����<�jx	h��� ��qEY����N<�[��;��g=��b8e��H]#��z<k��G|����/
����0|�9�-~�ڡ��eJ�ύ���B׽h��c�=6zl���w:ק7�n��ڎ�Ȕ��?��?/����}�k�R�ӽ�Sf+�Ί��я~4����\B!���������{�)to�/�r��!-�D�W�����>=N�\V!!n�{��8(;�����)�%:5���S�]M������kX���C�p��§�{3d@YDp)�87�?�����Ic��DūK�?�b����������*�����#���0����>/�����>�:����Ш3O�8�a�[�p;�����ܻ���(_���$ZƃHn�N(��[vn�9��"��ȸ�T�]nkq�-N���8P��
����T"��hm��2oAF�[�Un>c5�ŪT����?N����p|f2��x� 7#9ȭ�����)j����?=*(u~Mqj58J@��<C�W�)�݌���el9��mM/i0g�W�x�����]�t-��c�;$�ۓ�(�:Pa��L3@rc"rH�?��Aq �5"x�
��;$�~�Y<�s;�>��Y=\�3��i���_�]#*�^>�A<�dV^[m�K>Z2N��!���dRۗ^zi|)D�c�c�;Bjȓ��T/m0��O,c�unLO�{��$��>8�fb�����JmV�皾��dz1�]�r�'��D���b�u��X��)��|�~��89��I���9K|���pI�n8��xC;/u�eW���S�=)�t�fz�qa�163ٝ�;7��g�1�a,��-�,�<�[C�{R�/��~�:�e ���z
>���N��6^zȯ����,ZM�Z9M&�%}<�'3�Z"�S��Ƕk���WS�V���͊����H�<�zٍ���9�sfax:�ZY���>K�լ��7���8�i�����0���K�t3� 6l� Iݖ����:}����Dle���[�V	����哷S�RCY#��݉�Zg~��Ie��_�����Z<pq �O_��V=���^j|Y�"""�z�>P"Y[C�ܚ&�^<�3���e�3s�/ܪ�E^V=?+���TaȰV>��������c<[�[#Q��-��V>��珶��J���� ͬ������\׉.YH��yp�ā�)�Yz�Xz'��/~��*�V���狄b9 G���T�QL�<V�.��~��հ���頋}��ۍ�1Bb|�ۢT�V�I6�jȶ�S�W�����7�D`%�%A��1x,B<�g�9*G�G3򎲈X���1����7�߯K�a` ����?�1��>v��c��������Q���&Z2���E����n\�OJ���Q<����og�J�g����If�r�ܱ�2J�F��+���EW=_�xMIE�r�w�%�2�Q�����uK�2��X���n<��O�q@�N�ե�H�Q=�@�;�S?ꬎ,��UyLU���my�D
��97��Jdkx?>�ós-� /��a�}~POd�⠄�8*�C��բA��xI)��wB%�Ge�=Ӷ(r�[P��*��A��USJ��sO��Y�z�Є�8+� *�8��'�qڹ������ިe���f���p�[n�e��3��-! 1dy�������|(C����JN�g�L3����F�c�=a-RSU?�YL��NDt���^��avb��oɘwB��s��;�_���Yb{�CB�=�)���������o�"p9;�}m�
c '���@pi?fs<�
u��%����� b(�lwc��uyn��?	��������_��P�o��{���^�����ܢbK&
<��3�~\��܋[�L�.����3>��F�1�2BZ�NS��m�����JD=^��k�w`!
SȬ�L�����(`n�gVI�l���)}��I�yo��D�)_�/2��!��GQ��{;����wO�@�!�V�<R��S=���/��v8��a�|�_��Ʀ���$��B=�C;\�ePDO�}G�!�@W���$����ʾM"b`��!�T����o��Lb|��O�E��	J�+�Ky.\1��M���ci�W�?�3,qQ�˧�CFJ�m�=Ʋ�=��A=|��>u�����[\���s#xl�2�������<�"����wG"�|z�P�3��e f���s�<˰��J�E�}D�g캊�W� �}�u"C�X��di������;�؟g�q�c._����e���V�<=�@y�cN���Ht<>�3o�eX��e��iG�6��<L���j�7L���*,A���p�赽�{�d�6b�^x�׾9|���zj��;��P�"%��G�B�h���u�9e3^`L�:H.)}*^�D/��_�g⚄M8��*�ޏ���������H��Jp�⭍�a����q"�ߥϥ�9=��dǁl4�cj�Rִ>yq�R�eJ�-L�o�d�M,�B��,��z��:ߔ�X ���-8w�ܳ����O���'~��/G���O����U��隷�+Z��(����
R��z]�bX����V��$1렭r�
"�uO�o��^[�Rz�Deℰ�x'~7�0��b��&�=z�K���G +^{ڃxn�f��B��+�Zyn�.�(�7�=���=us�<�ڑL3
��V3�w��e��ć��8mɴO9�EiPr��1��J^�H�2B�L#����_e�Ķ�D<�σF?�����֏��1A�,���C�� q,�!cF����N�f��5C/�=�裏~d�- �0>���[C=��X�"k�Y��͇�P���>qy&2/�D��58��dǍn�I�C+���k%�%y��~/�_rP֮�cOv�Z9S�J��U-����8p���S�-Z4�1�x���y~_��mƍN������*}������� ��Hǫsˊ������/�^ہ`>;\㹃&�vvv^�3g>q�[���'��40^e՝{��҆	�*d�˜}�=[�>�v˭��'�{B�N1א��r&�3q�+շ�9���u�3WL�e��\5�+;Yv�=�l�~�_��_cL����c6�Ee��,���g%{"�2���Ȇ�D��3��Q.tą�}=��A�D�&�����b�AA����⿹N�R���G^��S��Z�~�u�I�+�D�fs�H`���1��q��΅ �;��<��c9r�P��0v<3��o����F�]9�0z�F{q7��D�F���+���؂�F���a�����q��fo��%%�A�5����'��N�ɲ䔸W�o0����]ɦ�*�)�Zc�2��(�M��R��	nI�J� ��ֹٖ�L�JѰ�K�˧Q�~xo�%��O�N�X��Bn~���A䛟��g���k �/���߼���>��SC[��L�����gn��DnȺ E$�F��ډ|���F�g$�/D�Vˀ��`�}�=x����ʈq����1��1�q������ܖ�,z�Wz��g�;�$׳Ba${
�Q�<�x�<��=�-dƽ;�ۖ�C�x��v����$�����=�sQXj�����>���Z�9y��,��*��l@_���.�ť�]�!'�ֱ��
dEpcG�)�(�ӯQ�<�zW_PC?R��o>��#ir4���g?{f��o�������H;!Z�B(�Xf�H��3|�9�����nx�9��q}�}n�ĸd0e�>֭T��Z�ǭ��+9`���w�wO������@��f�����~�b%&_�3����];��6����s͊)���a��3���R0w}����w�=*���Y��_X੟���'O�B�o����+�;w�y���#��H�������A)�?��կ��GW�,�G�h������gн���L�-�q��OD�p�fj������!���yۉ�/3^c�u�WC�5���r��~jW7j�[��^�o�y�����jw0�"(����N�<ăxG�(2���dNq��o��>����@���W�� '�,�Q�06{�Z�=��kѧ�L�e��h��㘑u�[��ʰ�!��ҽ�K�Af�y��Ϩw�l��n��ӈuc �G/���qF�(=��we�ُ�������g�~�7�~�Ѭ��Yݏ�k9 �.?��8�t��1┅c��ͺG\�P�9d?C�s�w�=�ϥq�em��z;�F�������Q㕑|װ��@3����:P�*^�h�@K�+��uQ�[����F����`���<�J�r�g���P�xr0X�	��y�G�J^)]�K_��b�����?��->���W�2݁d�ρ�?�O��Oc|����&�8ǫ�����Jb&u��� �7�/�b,��e�՛�X����yre_��e43��{$�LAFd ����)��鋵 ��@~�y��^ZP� 3,�=ƍ20^�?�y�%��;��s�t��/���Hv��x}#�^%���@�u�ܫ�wW��~C�=��y�(��h�oA�j$ �{U��ez$z��g�X�b��r���f�#���,o$딣�c�E��>����_��?�я��uG��H���e�1&_�˘��H-����Xf��⃋�R�Ap}����]�2��b�����65VE����x��'Q�k�p�,daF�|�@�ck��]K�O��!�w�(�s�q��2Z���\��B)�O���2�:ә����+xNWȟ���W��l�=(�s�@�E]�Y|�!��L�������8�!U����]nڠ�Ք�+ڑU�$�祿��U���*z̉Q..�\d
`��-��`���� G1�kTT��ysbW���ףֿ�)}��r�ɱ����+�
~����T��@/� �q���x�L
ςиvD���7yq�e��Q$s8x�4+!���b'�TqsQ���)q�<Kʸz������9	�?{���{�Ga\)!W2b(ݏ������<��I�d�4z��nZ��6�O�.cS��}��A����G�^�ˬ��G��C� ��/�m��aC/(U�Λ3^D#3#��}�옺~4�j�����(ΐ�g�~�e�M<�o4�0����#��#JQ�d��/��"�k�}+q�
/��NuRuP���<��z�@����%�������u�]w����~��r��~�{�[nqʮjlp�w�F�\�%��	� ��Ֆ,Ѓ���0����l�/#��%�=��X��&���y:�u��)��:��e�2$J�B~��f-�2*�-��{�*ɑ�މ�Ӏ��1��_��CN��d��֞��ꔮ�do�\y�dȪ����P��Xr�س؋ǃ��������w��z��ܺ{}�zn�0��Pq���6�ko����Ch�G�"/���߾�q&��`����o~��0�~k�`��n��:��N�\���,�v�؞�����'˄�0~�~�U�RI�j�F]�Ŵ{n�s?�8�ڸ�r�Q�kc�����@�n��
��Nr#ao!���ǂW\�2v)kҶ����@V�H.��F��M7/7_�2���>S*,�� 'o�neJ��_��_~����^~��g>���}kPO���y��G�j�w��$�����U�!��a_8 dƟxuKf�8,ys�l�"�3#O�HA?�dI�1f�}�c~/汭����1S�L'�_�ͨ��QC��dJ��t��7���{=�ωU��-�{�YQ��K^�l�"-b�5!�e%X���s�ȞM�}���~ygJX��􌘭�:�cy���R���P"5�=���B=����/���+��DޘV������j9���ݖ0������=3�H��t?�x�[��Cο=��,a3�J��`r�P"y�$�E3���l!�%'��������x���,��/m�}���_rx�)�h��V����G��������#��m����h��N��wz������k1�����$��H��wJ�򕯌��_��W?�
����AV�@Z�泟��k$~V����N��y�����|�^�}���s��Hn�\"� �[�^yL]̞���&B�3e���~�^�"I�/�%�X�g�<���{<�c���wn��Ĭ�#[��uB�C(<�$z�y�)pM�]����{���"�,��*ϲ�!R�}/cY��������4xL��q���9��{�{��i]dmɠ^N[��x�Ic������F����&���2�}�k/|���=;|ܑ��gmht&�yvb�1É�'��BI�b�)�AM������81EDk��yQ?՜Y�7�m�9����C����YJ��}�Vv���9רYQ K�kq�(pVX�ji��S�6����*���O?X����ޏ��������}�s;E��]A�62"L�����=�^6�sE��d����Ȫ0Er���� KBqJ�A���:�:r����q�rP�L�<��:�bo='*�._�#�Y-�q/�,��Ɣ>��䞎x_N�=g,7�����2Z�d����[�z�`�v�תrn<�܄�H��HZzB�F_K����GQ�����2���+����;ߵ�7�!�3���{vw3�C��N�e;_7*II�/��<S㭇����-4˰I'�*e�ޏ�H� !��JΟ�ker�N�Op��֜��V�V����:$�k��S"��:e��k��ws,�x��Q�_ �����曖�e�%8��L�]/����3�w�]�x�nq(��ݝ^>ָ�۞��x�G���8�p�Bf�'��G�C =um/�w�ș�.�a!3�Z�=zgJr�����?(Y�cϲ�y�,�jF�\�����Ț{�| ��L����A��v�M<c��XѶY��X��`@�3b�B�ׯ�ĕ�y���_���� +g�fv{��AnI�D����S˨�Z�Mz��F���-�t��l%���(�:�s��=��fZXv�-�|��!%������ԅ�@ gd��-�y&q�Ϫ���u���(W�����ا��nvM�I1ˁ��uq�;{o��u�}�x�Ee�5F�������wr]s�g׫�^j����O�nvN�b��i%�NA��1W�boq�he�K��"K��+��c�'�l79�^���[o��;�C -:{饗����w�}cnC�,U��=ɀ�q������P�X�K�A�I=	.X��My}j��
b	�`U�\����*���?j�l�;*�LQ�B���X�/�Q��(d���vc*��N_ThC��H������؞���YE�+�݉	�{���9��4s�NM,���/�-��cf�y���G\ɔ0��1g����	;����t_ꗄ�H�u��Iݔ���)�g��b�SȌ\Σ/XX���lANnt��4�MnذD�)�t�0�>79A��Qɋ�i�}���b����o�v��"R�wa�$tb��C/8)�C��7�:�����R��5N�q�+1{P4ҳ���r�6���`�b��FJ����q�)�R}"�,�9ވ�=�ɉk�RW��M7��	E�����:%尰��w=W6�P��AQ=��/~�-��r��jE��q�%B��!���;��#2����@$���"�[{7P$��� W��켨��Nvf=��2�C IS��T��{���⹘�*Ư�,� S��yb�;ي���*�g�x�5�ڏ��&1�N}�A~|jU:��Ylњ>�2�K~v�q0t"�mK�C�O*7��� yg�~gv�v���Ov_��W��ed��P��~fج�7k���5F�TV��y?t��.��C�������CIn������ߟ�s}J[��`78�Y���p��3@�=tPh�X�A\;7�����}��cY%�,�~f�e�u��.�]��Ec%K�]��5����5�}��^FKc���&���*����JP/�+4��/�az
+��9�;�)6���b -��S��vێ���YAN3�
)0�_���ޥ�hw<�#)\��se�6 �dFȦ�a�Ģ*2H��i�)C�3	x������>���[�ly�y._���@3سp�zV_��Tq�ɐ�<��8��G����dh����Z{d��4g�^�Y�-�=r��/<��/]�7m��>SC͸(����e����>���xB
|᣷��1��c	3A������ü�� #|�S�ڒi����|��g�|a��,BfH��O�:���$�˜�%=R������qb��T)�~J�+
:$7�����[�Z=�Fl!� ���ΗSʋc������7v\����?�gM�A��vPX�A�����>��/>{�]w����?�������E3D�,ƥ�cx��\xgl���L��Hjď����$ӱ���s�z�e�
VRs<r������Hb����)�U�T�`�P�{\$�-m�B.��t�_�oFl��s�^|p���D��43�����KI���R�"Y+=�x]��q1L��j���q"7z�/_Z�ev/�[��_�{)���۬<�UrB�Y���Xp�ԧ�!f������Yz�.�U����?�88s��q"Zǡ�7��8�%���_�֣4xYB��|�W��xS�.����5#��O��qȌ�����jm	�������8��6U�M�W��ׅ���2����}��Ԟ���ݥ��7@�%��������C�>����e%�:u�ᾟ���{w�G��;e���N���jk�eJ�l0l��R �-c0#֎m�y��!�MF@��F�������4�n˼u)��Ŷ��e�D}��c$�L{����xE��gI��'a��h�g�:��V��D���9��1��u� ��W���Ȍ/�I:m�rh��L�;��l��б��bd�����Ku����7|�~��X��zg��������"N�#��<��
����,���:��-6��I� ��������2�픇S@�{*;�b�S	S��U���E#��L�k�~�9J�{��S�����r)�B�<d$8Hr��Hyp�2Vq��`&�~�7.N�tr��,0u��$�y8N��C�h��~��gz�)rx"p�?$�Rm�AQ�	r��P���c�,gF�c]�v�
�˂��>%?�E��1w:%i������L��LY�-��>�^F�>�8���/s�z�`�=$�	d��T�e�?���iJ�i�x�@̙>v��?��s�Y�<�%R8�#����9��XЬl����ڕk�e�"!�T�{��5��Ǐ���QQ�	��=�ɦM9N��B&Ї'p���yvХ��!��b�؞�b��db��%p'�~GߒJ����5�*"ӯ%ː�)=\:��h@{YY��tr�08Hnu W�A0Z���Ŵ71��c�AMi׎��@f�Cr�n�FN5]$�NGܭ��d�)'u2:#��.�;���zeu�w<7��S�=�h��Š�7Kc�.^Z�w�}��w#l�.S�2�+�"?��'���<�"^��;q��1,��'oNȼ�󿧼
x��@�� �,�1���$%�.�Sf���$�§;y��LxV���������,�/Ιұ����ݝ���c�B<&�	���,���m�Y#1���vqlY���dK���W�����{؍�ؠ�5�V<s��rљr��ܑ����� �[��i���]���H���2�'[X�}�%����r���:&eu�Hn�.�����X߬��4�$�-�d�6�G��@��bWQ���|�Ɲ��1Q��ަ���>�_�޽ײ�8�]ݽmcc /81`���K	�(ji�կ�Bʟ��$R�@�d��!���_c0�s	6���>���]�c̹�n_��׼���z�F��s˦"|�`xX6�WS��=�!����������n�o��g�w��=�ǭ.ǁh�����_���vʎ0�L��q��\?Uk��^�ʜU�K�\:p����7Q���V=�R�6�RYò�Іp�c�K +�B�d�R��,\X�!�_�g��~Q�o~ĲL�y���ae����++�1+��3�گJ#�=bE�a��=�<�j}��P��<����$���|y�]����ƕ%��[?2��YV��6�Q,Xҁ8�������E��3�i�mL�XOc��2����.O=*|�q
?���[2 "H��eieT�'��O�ۍ�P��a���+K̑z����:���w��;""��:�uo-EM����G���^�7s뚮�!$��$��]	C��	u��)�L�&�%�����aV�:-�����U�{ @�����=ϑ�b,��(c8�s��q�HFѪ��BH�Xa��&�H_�C\d��r�Y���F���~�^d���E�`q>Ь21��
����/��Q: ���Q�",�[��b�q.J(J
>Ԭ�(?�W�)M�'�	}��PP�?3�F�y_SX�>Q�鋸I&���9|˵ڐ#y��b��9���ԩ�xeLSO��.�2�<Q.2�V�oO����g��hƙ��E�{����le�ոR���/�7�1=wC��B:�����d����)��y��jG�,J��9���.d�a��?Z����c�~�Gb�-�7����wK��|FY%�	����W<��#���m�d��R�҄��{�<�w�� �[>F ���ቯ�l�����{�x�&�7�D��A�T� .�����-B@p:�tP��'�0�8O2�8���+
���@q=� ���9`��[+q���@� ��nk�W@�J�7^J��C�B��@�}��|v[��G�(B� �[��<;�q)������A����	���Ҽ�{6���g-d��������|��ԧ�]L�,�ݲ���(
���(/�Nװ�hg���c`(�\V�Ǹ�d0�[|�?#���g���������ʏ�ƍ���Xc��4�䒠�n�4�A~��9~�4������.m�dQ���(�io��DL���M��㽏���qUmUʘS5��Z��gi��E�� �0?�[!�*�fغ��u��� �Ү�wzi���<��9��	@Ga�|;�;JXώvo7� "\)� ��&�S׬��E��#p&5
,2�J�#���,��%�]��>��Rm�z���?1��C��*"��c<�{�ͳ�>;�0,�1ҁ��a�\�9��}�v�˝� ��Ҡ�+ �Х�\1�L܄
��X�}�5Sq|�Rx��5�3�Y�ķhVS��~B�鱹1W��O�/��N���f�����8U:���KD�x�@@܌�e`�@����ڔ�>}n��Hl"]++�ۨ�1�7��&�
�e�W���ap#���s>7$��lN��%y.�d�M�j2�B��Ѝ;K,D����{~�J���|��ꆦy�m�����#�b�"`�暃�ʙUFj���,Z �;{/�� �9[�D�s��ƍ1��_�n��l-a�Qh�� V�A�?����� ��4��@D��m�}㛯X��P�r}x饗�a{��qѤ�b�������g�%e�ڶ��}��D��M{�f:�坨����<���a/_Űzd�b)������{N��\�K>n"��u�݃����]e��uc��H�[��M��f�0�q�����R7�@#Dko�f���t�������D�k���NQ2 ɵ��m�mQ�:��$ |L�u��!%�4�|��7��ڦ��w#�T�����B��am�;�t���V�u�=a�l�����)��j�8��P�*��#c�e���<�����(��u.g�zk^��k)��s�^|wk=!�<�`�Sa�z���Te�b�0���'Us_��������?�o���K�q�xd�1�J@��#%���XS���<�>����"���_� y}*y�)Y[�|]-����9+�nPu�5*^1�
n#n����G���H�S�P����G�՗/���\�Z4�o3��$�\�ټ�5����E��\�N�A{�����1�Ѽ]C����� \�����"����s#\ER�����z��L������]?)��7�r����X�V[C��Qkn6��k�3 p`�{,s���[�xǏ�u�P���5�>2��v�53[g|`�9:�t�yL�\�"�( #.��&K�qc��7�Z���E����q�%Ht���o�������:���`�⦃��)l"S����js�ǹ���y���v����o	�ʰ��!�*���9�|B�b<qe�F�KG�nq���_�2!r��Ҋ��c�>�)՘�U�f�9�=���q�~��FAn�F��Ҁ[�����m5te�\
:[T�%�TE͢��?�k�����D�+����Ɇ�Z�$ n����S0q`4,or*\���G�Ũ��V˼�'A�n�lp	��]\��l|�<s_[�[$����T֧��a-e�{����"��2���}d	%~(��75A \E#�$���c�'es���,z�b��^�b��&��y�c�ϫ���q���N�}³��Y����uy+�Ϝ��EyG���� =�:ʹ�Z��ֽ�����8{ǟ�o�Е+W@u��7%s�W��P2�Q���ݶn4z��7����WNu�'c2�`y�߰C#cvt\gx����_Q�z���8?\�����8�=!�ݯ&�.`uW`�3�"�6G=Z
z�den������+M��E04,K�������nn@��f�{���nr��7�  ����Q��&�i���s����qQ-g�`���`�G#c�W���^��K�5�"q_i� $d��� �ǣ� �}���S�E~��Xpz�ܬ�n���;�ǣb���rЎ�Oy���5N��ۨ(E�����࢔�4m�~���,��ʆ<�Ĳ,���l�̋�Ķ�{�<�kX\Q�������K�/m#l���}���>��S>�;v���d�=����ð�"$^���Y�̉�B��ܟ�R�+e�)����|�k��h�A$�=v2@ޛ�[��Yh<���U�ʪ��zf�^��#ߙebW�UV���C_� <��I�e'�޽шݬ�}�]=��q�)��v��KX�!���n9�JV<13_������e�����Ϡ�p����Xd܇4�nak-Sf �˶tί!���'@�A&�+*�N������ DXlc�
�B�Pr%�/�7<�������8 �]�NKy\K�O��\�
�p	ъ�����\,�k������`���[�_���1	w)��B�-$�n�V�8��C���w�������&�����es�j�ʥ"O0Q �������+W�OGh��a����a�[�o�eը�o������'���*�����u�#�*֪�Z���z�7$Ki	�핷��� ����##����^�r >U�d�����3%�67Mmp����<D�HH���?�:[��|-� � z��?z��+�IK;n�ϭ��nCA��l�ݒ??;ݓϱ������4�Ȏ\ߕF�sF���ZX9��b)��BiWN�������m�j��Rd�� `'n�,N5$_/*���*rת�-�エ5��x��kG� ��AT	�=�`��U+�0�J	��K7be:K#*�;|E��,�4^������k�+l��~r���IW�tmJ�p�}n�y� �	���?8��c�m�*��X��e@߸,�����"q�ｏ%�����-%��Y�����Ȫt>��*��=ӫWKa�����@D���^��J�
���b���1��ګ��������G`�>�ߟʡꗿ�����?��/��!z�x�x[-7�c����d�}\i���Yw[ڬ���[p�9��8��a1vo\.���<�`������w��|X�$;v�{]�@����խ5����G��c�)@E�o9�OD4 ����X�;��v�#�gK@���uWD{�Y �l�`f���wG��؍�!��^����k�	sw�������8���r���M�7�ܘ�ɹ�]5_�n�ƲZ���J��B�>�r��R��+�3ސQT���"��42^�ĨP���0�C�!λ�wmn����jb��I	�hT�>{f�]{�nܩ�̜��#���y�?7M�=7��!��[� ��,����PCgV�J!����lBf�!c<.�b��p=䍏	�9�@�Z�/M?k�����{��	-�\w3h)���뛢���_�l����C�E!�� ��f��V%d�z܌\��4⽊2>�e�*���F�����P�GI��_sE�呷�GOq~�o(��O ̕\�"®9o��#+�������"�]�}�+�[�f�-e�c
��-����e8*��؋�����e���{21�ㆉhLbGP��}���@\�9�*��2A�4�J3���m��oQ�C�b��o��m���G͊XrB�c��DS\�ECmI`~�);a�\�E` ����]�pK��}�D-km��8S�ɞ)@�wK�3�H	�r�r;`s�W�l~.�������4|~���4;6�xh-7 �|曺z�2���)3㿱ieA.1��y��#@��_��W����~{��5
�S�?2��1i�����5p��\���XFv���� �˦J௑?Nq�s|���g����?<�_#4���{���s�?�������n
?��O_|��s�3j36�b��n7�Mr���B#��Us=K�Jik�F�����Gύ ���hY��(D�bD�Eµ�<���g�Q��D�5���(��m�I'��& ��E�Yw���ú��x��&(��!)R��S�]�_��4x���p�/_c]���h�Qdi�a�D"�
�ͩ��!�j��X��ۿ����z�d^��fٵ}^e �{<�����H?�
�
�:Ճ͎:.X����gw��()[w�h��Q)i�1G���-��^2]ݏ�6������8� ���H�>�[3p8B@Ud�kK凗��k�h�F<��f���\9��A�(x��9�n�S���É_�~�rO��ʡ�?!"٫�>�(��� p�q�&(���'Og�x�)�~���:����.K+Σj^yZ�m� �c.
1��Z�`+�X �ݪh�^�)E��Y��%K>�Ps��?�߼�Ϋ��M����Jc;�pC-5X��)��H�0�-7߲yǭ� �l"�6�xۺK@E#B0�^�Q!�f#m����eH�O�Δ�J���Y1�}ͧ��<X��=C}�2��&̲>����uj���NL�r�7߲�b"d}����Z�X�����2���v�b��ݫ�s��� �wknV�Q��Z�¼jW�����}?UK�!$�@^w����V��[ˋ/��qsC��N���H������u�A/x���D��W2^����O�eLf�e�BV���ѣU�?V��v��R.��2m�)ޯ�}ՐY��X2�2���:�%�c�U�U^Q�qk��	�x8���Pn�u���LN��Q�s/����w�q��^��F��!�)��q�P���A��r���ƚ�ג�Խ1���j\d�c'=˘�����@,��y}��A��`��e)�>h�u���߱h�����w�oee\Z��{VP8<�<?q�\md��ϱ�5�U��8���?�B��%��9��5�J���\{�R:6[�s)��ۘ�H�R�*/�|���r��#%��v�x�Y"p��X�n���o���/��O$��#���Ǡc\�1���f4�T�/�8n��ſG�ʈ�&SP=�5�r�|�mµ��ǂz����~��Ye����ҩ:�˞5L�[��(�G�Zye�a,%nPc�i1����﷖F�1ZJ����m����d=�)��B�L�q�`�j,=lTQ{�[�Gm��85J}A"��DZ�÷Q s67�m)nql�@�o8��v�P�f��+F[��ӧ�a�|���p聉�O�/d�-���r��+�]˳����(	�)&��o�Z��g|+>_�Q�.~��yYE���q.�������l1����o}�[���Y����L 2N}�^��c�Q�`�;�{��H��D���k[(��R
D,�{��x���t0F��	ɦO�g5n���p?����������瞷��x�����W�:'�����g��`�۟���+��K�+�^=PȌq�oc@�n����er���^�ou���Fy~F^���O]��Ăf���\*p��GKB$�L�\u/���D`�iV�������H���3���ؚX���Ġ��&&��7�R�Č�|��sb2�S[��`�=�s��tծ� ��vW��jo�"�
�ZL"RK	�ƜGup��6z©k�WP�V��G\�N�F^Ř���_�JK�,���l�z�o.����M���>��M�q�j�|�Ea�(
�\�X�e�W���׫�f�OcDڎ�͕׍Q��z��Oo�:e:_��[�{�l����
�+��yV�|�3�1�8�ce@�d�=��p��/|e�65����8�d��&�p��%c;��$�Fo��#���Ѭ����g�cD��D2寢5��"�dc4b��X��1�VQl���G���@d/E5����n({��([ZBń[Ϸ�JF�j(-F�'#�3�8|�,�o�,VZj���KM�ħ6<�ʆ��vR��U126^��� }�<C��SQc>FZ� ���C �"#�����O��s�c�
��c��962Wb��&OB���D0��q ���xz��@�b����z��R�[�JK���CE�E�1�=�[$�����w�������F��4�P���E���5�C١ػ\غ������3ȝ��޻�����׿��/��@�K/���[�H�Kd�섐d��ǯ�������nl���R��Ik�">�|3�0?�\�����Ȁ�S��Z�~O�����-�DhzYz�<����E�������Xw?3��g ���|�����XZ��}�{�s�������ێI9=���9�A��[�������;��LVXN��5��1i��� ".#TZ3�#���k�lS n��qp���+�n�$3U���j���_	��w,���� ��0�
�g���;�H��r�4�uf��ݢ�c�0�<������Z=?
�n��GH�߮��|�E�u1>���j��
�J�~�s|{���4m<�9�n��7����1�t�=	�fiuP|�g?�����4o�vV�g�}��瞻��e>�p��I�l��!ڎ����f�0Pv�O��Z6Fv��#<,�7��}`��-�D�� ��\o-	�2�V��t2F@Q��*`Ϭlk:(�˗|0�C���ʡ@�(�_i��)Ix�'(��3SS���rz����~�[�:�ӟ�t۶�\j�V�O ח�����bvz0���8�a:�Ώ��UiEE���=B��s���8��ӎs���y{�d���r�ʥG�8�"Q<< ֏��y��W�X�xiq�yB�>&�o�� ͔/˾ .�c��g����gҗ" <�5��}+Z'���{�$��R�5�8�+}��:����<��\�t�����ǃ_���6G�O`�+??�g�����?K�_��2�3`8��{�V��GQ)��ct�W�o��b��L�0T�������/F��B0V�Ũ�>2���^�C�:���Sh��֠�����r�O 3�Tz�P�G�w����'����}�mr'p{8�үMmsV�"@(�ѫ�P b�ƀ�Y�h�,|�#V[=C�&�w��z㢚o���a��0VxG���?=�?�e0X_f;�����<�VU�,��Jc�c\�!��և��` �6��Ȝc�y^o���x��(����V����?
ʬ�w!w}q ��a�N��ɭ�Բz�>�W=��b�zJiW�Q����.����+ 3��|=v���f2�hs��/�|������'�x������ �{���|n���Qf��ǧo�C�Җl.#t�o�� w_c�<����w��zy��������25]z�d-��<���*�؁�<��6�Q��=,o.�hh�|���W._�[����`�i\ӻ��-�)L`�+/���Y��$���oΏ�q��Ou���/~�/�@ܪ�e��Ї>4/g����|�� @^�4�j�D0�%�!=|�G�
�;� �˥�-7��pe5\:��=o���F'��h���q+����b��Qp���Ɂ\�W֎՘YB1����˄*�P�|)؏"�7A����k�,3p��~/�������m������8�Kw����G�΢o>�Y�b�VDc��/��ɟ�}�����x��|���O?}8Ɂ�M�������l���2(�"c"x��&��LntE8�-�a�����Mh.U�z�y�-�hU�8�T.tP�z�GF�i�4�ٌ1gB!�*�ю�U�I��$ t�D,�t�ȭ/��8X(�����y�q]�6H]ܼ�hbV�/���,�l���߭�DL����@��Νw�9�P"���#���_��|b�|q�l-�X8*����ƾ[#��xjL~6��k��	@R�,��uT[�=b=��G�����r�M!&�q0WRx�-�1�x��9��B��=z�S命W=�j��L��y�[�{暫����~�<�b���¥T��ak�\� �X��׀[�;|Ή��g�BҞ�y)��/�5rSx��G�/�N��-��6��+�8��3�������.="�qQ�v�ad,��?�Oo���X��ሼ��} ���qZ�����aJW��g˓̲yn�q��jL3��3#���iF-���8Z@8�)�����4��6Z�k��Ƨg��@���&�W~�������7i�o���_��+�R8�m����!.�a �-K��s�P����z�]ĺ��L�X���E�U�,~=0H?��(0�����-�ѝ"��O����7�Z���W�5O�~6���݁����q� ��<D���h�hYF���u���YT�H>6,�zی��]��D�A�pbJ:ʙzp�ḩj���y�!Zp��1Pd�X�!��ê�(Y�b_�ʹo���\9����P�qIз l�T��4Q���x� ��?�����������sUP��g�}�~m����WxP�4�<� '���F�xLl�/��#�8��a����d���-�2*��g�4���KZiĹכo����$3gԙPZ�]��X�D�:�b�K�UÏ0��{D$ށ��?�S�ܗ�cIE�R��ʗ'������o��4������/杰,�� j|�������C��,��ޓk��e��[�]1�;#�@�0�� vT?.P����&Z-��Y���]3�3>�k�����[w����z��wJ�E�����=GW���k)��VO� n(P����g��=!�ף�$�/<��5��g��� ���ҝ���֦�̣c*>��'
��l.D�� 2yǤH�/����c�]�}�3���H�0���H�\}�7|��$�y�K�<����{���o~�_���������~p���{��g�9+����t�#�&��E��j?�q*��Vv�M�_��}�p�{���#��z�U�̮G�䒧�q���0���Pk���J8�J=�{_���7�БX08nA �c���}�f�ߕ���;�����~�����-à")j�T��K%����+�H�% jY�Ӈ9R��*�����`��GN��������XnE�8SĈu�h
�9��/�e��'n��L��-F��3�^[,!�;��F	)�\}���$i��eN�,#����-�_���x��������)�\틥Ϻ"B��(���%ujT����*g�>�B��w.�=P[Qlߘ.+�1�?����+؎�N�iLk>\8����'G=�N��������7�zxx���!�B��^z�K��_2�'���,p�L�~�jWNԳ��lWBD���Ǫ�g����yf�Fʳ�z��7�b��#�?����c��--�ߋΞ[C��q������]4��I�.Ŀ��V�K�����0vk�6ZM�p�����>���G�r�T?����N@�	������I���"�~hr?�S�ůV��.���H^�=H!�s�$ȵ���F˂� W���ns��49��r���w��>b���W���ೄT���J��w,��w"�D��[Y�g�i�U��֢��� Ǐ�K�~�|G+o|�RbZ�=�u=���be�x��tݚ�	x�Ј�v�� [�}-��e�t���s�����}/e]��
��t��敋�̿����p~�Ƃ�0� W�E����ٻ������_���>������$��Q�g�&h�Nm�
��Q㛨3�f�����V���k�1��X�������@�U�ϒ�͝��膌���&����F���F W�g�R����h'=� '���F�w�����C���^n�=���Y�ۼ�6(Z¯~���:�}��f�-�+��oJ;4o�F�eO�!����o}��wO��zOiK! V��h����#��=�0c���F$��˘��(x� ����KV-��W5O��A��L12"�p��Ѥy�0K"��L,�ӆYv��?����B{<��`y�c�ΑU&0s�ͷl�n����%��J9��e�1C�=p�q��V 5*iUޮU�}�]2��Z��%�̡슯���
�1��q?�/�>3�/s�#~�Xy�,@۪���B�i%d�����}�ч��ί��}�{�Ȓ'�x��������w��v�-A��#㊀k��ͻlV��O��Xvc�:߸*r �f�� ��#د5�Gx�ϕ�_r(LX�4��kh�l�k�L��^Z�Jh�˺;*�['�tܺ��^�2$�@f%Ц�8i�_z�g�q��M����9U$��M?01��rK4��}�_�[��Y��ec�>� �����+b�b���Ի0~�Ƚ~�,\-r�L���E�+���x)'c�-����e�ˉ ��T�3�ܬ=*�G- ���`ف��&8�ܗ���'m�~sn�� �!�T2 ����t�*!�X�-g�D��2�?S��w���������'�w��!ٚ3��cs M��}x�yQ)a#�5�1{'�!~}	es��_�7�_�A}�����Rc}��|4����;���,���H[�F*x�x���އ�WN�N���&�������~���=��/|M+}���#��rc �����l�V��R�{��x�\u��8�g�T��L��̏����?;p[��2�[(�52!�&�5e��S��v��,��愫�+���V&�����4M�/O���SV�&A�of�+p������_|�B���X�Uv��pNX'�N��d��c�h�ى�郂 ��k�|���%�!�ː�]Qo|d�zB�%s�c�dLy }������{I[ 5�U]��s-e�ʳ�pf���*iI���o�Z�������Z	�HgK�U{��Q�ȰIH�W`U��/(,(������JA��Z����Pg-�:y�3�G�߽�#m1��k��Y�D,��t[��֦ά�"������v�M[c���z�W9�4˪�ƴ�r��r��i��#�1�{���w,��|E�,�;��1���������t�k���������>���*K&0{8���$.N�[�����y�>j�	w,�X�ն��-���� ����(�f@{yܽ�zQţN"��W`wm�\���󠺱kţ6ګ���C�]屔�s��v����� c��gPM�Nk���X%FƁ<�ǭ�	c���zOVP]��g?���7���6L�U���r�4���H��V�Yfb9Z W��*L������,��b�r�ߤ�֢Q�@x��o��~�(6�7>�����R.���-�_^*��_�;~�2p՚s�� ԯ���jhg��5ߤ�h�Iе�m�^��#/�,(p��)�ʠ��7"f��3���LUG�Y�U�	q7C���X���*����Ǵ�y���9���q5���Ƚ��(��F��T���ïG3�t�A�k_�Q	�)���� ��~�xd,��C�ܻ�b�`a<��P���3u�,�H���Gy��}�����)����,'En�� �Nm���c�n&���q�R4��)��9O|e��	Գ��Am�irD��Q��<�(Z��&�#�
?�rx�7��P� {�%>�5J#Bn�A�w%�+A��Y�2ı�l�"�?��"���l�;>l��p<J�hW��<_����������>o�;ڳ�����<�>���33���avǥvڋ9b|"1g���+]\-i)���E�p��#N\Q���&xE�w7�z��Q��6�C _b��H��u��+�3�<�@K^;W�P5�cdڏ�y�4��������m��2��Ӧ-��b�� �����b��,�c�[�������?��
2�/:�isp�U�B�Z�Dh�kl���C�؍����툵�?�T1O�O��}�7W�J��6,�-AY�5��L�U�hD��ʜ��?�t���x���U�eA�u��3F Bd����W�~zF�� ��G?���)�.���O<4���}of����T�s�ؾ8��s��dH	T��&>����˭�n{�63�ޞ�S�5��Dp�%1��]������qYa�]�g�k�R�J~�w��{|~Ѵ����j����їXȲ��g��T~gZ���y �#�&�;��|	^��ey�t�EWQ������Ҕ��'F���ݯ<��SM���w�q�tuB�T��LB�~�'l���,K�h�~8@P~������g���ܦ�����u�EgW [����V0�=ݖ�(�i��|��2Xx�U�����,^G�"yd��.�E����G�D�9L}� |Q5&r��E�& �q���~w��2_ ��ٕ2fN�k\k����?�D���K.�_}��YQ���l4o�'�4ۊ|}��X��I I�/ﳊ�c��#~�ءo����˕�of\�կJ�eUjQl/�������i�����s 7ư��0�uc�JJW/l��я~����y8�U������}�ݷ�L��>��>
�5ɃC�՗=}~��슣:��;�4=T"�%*pI�ҭ1�U������:����@�dl���0�a��-�;�^���y��#`6�������J�$������p�U~�tZ֫��5�ǅ&Z�&����>)V\bL@��D�QE��ĉ8JK鮻��R��~��G���O��o����T��jىS��1��t]L���՛��f���#f(�����Q
xH0����:-����7�P?-E��W�l~�ٲ����"?, @������g��:D�4�cI�F���&�'�H4��������[�x���,��^Xoc��I�Ǹ�N,H X5�J���O@^K��=�Z	�J�o+2ˊ[<c�"p�Ɲ?�DQ�RQf�����B��	鬽���v��"���)%�&�P�?�{t�q��
��� 0��>��S޳L����C=���W��-�fIWH��:�>��^��幩����:����=����9�Qt��r�񕑳20ừ�J�%w���Y��؏�w\%�c��
���>��|�<��w��)��\4���g�0oULu�|�gZ�d	�2�X�`�33�P c9@#�z`�XA .�Q�l8ȣ�*-M�Y�� �׾���?41��5�����Tׯ(���'�H�Kp�2��A�ӏd�r���$>�jc�!c� �YVc+
v((\��4<?@;��zE��@�Mz "��K����>��!Y��#�hs0��K��c�sY�?����婧�������.�I�E1�vc������+����sʕo,���(_l)K���L���K�Y��(O9k��zʸLxg ��1���,�4
��)�2�z�y,>�b������~���6o	��Ґ1aznv] �7�{�?V�P�� k�f� %2 ���2��%�Ud�����"Bo����;(��*��.��X�2�)�S�����->㲧W��~/��A'I��T���rU�f�c�bQ��eɈ��b�q�W�R�����zNڸ&�Z$�Y\"�b��q8 ��ʚ;1�É�����~��	螞�<3=���w޹���/ξTS�.N�������)���ʃ�`��έ�ǘ%LwE��L�!Ƅ �]	�4+�*�6��=��Ǚu�5|�E���\���q�1\���;�����~�1c����rg�ʘy67��1����c��]�1��A���Iŗ�n�Y��2�xA�]�s��# h^4�U�F���#����F���z�*�٪oV����F�?�� �ܺ�s�����[�o�8�w����==���'!�P�<"F w�`�8����7�? J=K��*�}F�[�q�T�w���>uz�!ǅ�ʾ��}��X���7h���+�W7��=�L�P����֣Sx>ߕbApK����T]UZ�P�(��qR�/�໪����6��4ȅ�}��6�|3p���4�P���ߌi�|bb�A%@���,N�&08\ 8��D/�S]�2�Ҟ�v��R�|���3�<4���~�����/��ÉI���vq禺)(�6Z:�O�G��A�|��P��(ąd9�C*�Kj�3���+�q����%���"��@�o�r��q�کc� �+����=�*Kr�l���h��v�GFV����Py'��z[�e��?BZcEV|�s��������1��>��:��Ŀ��[͙��/ ���78 ��)Zʿ�͗�2�fD�y{d}�}?o�e�Cc��N�_�U��Z��z>���ɘj.g�UY���r�8�h��l4d%��8�}���8C�����Hx��Ȓ�O�[u=4�Hi�v��c�)�e`{��Y�ȁ(l.�M��e 7��h)y<�-�NcM��#y��(�SF�����޾�!v��[����Wh��X��#��
O���Z~Lk��6+4��<�
T������.���*ߘn�pb��˛&~�b�\�X���o?2�%@|h��X~W�-mc	�/�����o���~��K���ƃ��?�a�*R�S.���?=7�}����N,+O����Q��F ��&fM�	,ٔ{�r���O�ן�o=���%��[
 6�R��,��w�O�z@>�%&�b ���B��><�Xj��x����(��X���v���}8�S�0vxΗ/{���ʒ�a� �@e�zD%E��ͭu-��J��@�z¼�3>O��@����4��X� ���t� �������Y���*����(�QnI�l���@)"wop ����\��f_6����+>̩��/��P�������"v-�E�2a�p��Ma^ڝ�����wm���A��0ưJq��l�gc��@�{�\=���Uc>�����d�H��g�w����]�7�[��@�(���~W���Њ�A�)0x��MY��	�4��u��f��>D"Nqq_],X1��oP���@@*FFŌ����$��vBZ	d �99�:�̥2�َ�fY�t_����W-m��*������cL��S�y��nüdǱ��2����1�k�����Z6�<��l�<������M^.\���輌B8~3�}I0�]���iG���$�J_�y��k�S�=�|E�?�9R���Z|�� E�����;������kXo}?��E���|��� H+�֦�(O�Wά<�m���*Hy�@�˗���ȁ��
�>�E2���&p��4�_2��Ώ}��%W�
({d p
?d���/�Bʢv�o����ܗp�����.�MF-%x�B�G�n��kV��]���{m����f	>u�e4(�T�0�%�5��5ZPǲT�*�����*�?���Z�?}� ��,C2���#M���z����n�
�y�gb(�%�`C ���o���I��Wˮk�����4����ջ��<�/��M�/Y�U_��X6S:���o�S�`�*�-�  L��C�XY*P[������	|cNL�v#m�?�3c!#�� &�-��"�w�����7�`g�<���G඄b�Z�>�"�\nQ��*�����%o~=>'��EK3V:����K� �f�����V
H��F�B5n+��s�/q�fm��<C{��x�M���Aaa�n^�v�|�b�G�jUH��*R�n�CMз�8p%�}�ql,�Q�]��w��7�uݨ�l�=�К�)J�#�Um�S[��ƆT|!�b�*,����ϙj�����-WL��z����t�?ZƘnV��8�/��/�����y�p �R!�M�V�h+��ջ�gzL��PU�{e�4��n����ה�C���߹�途%W|�<��'�V��)=�7�sD�,))m�	軡];>��nۅ���'B8�\t�<�����2I�n4pe�M��P蕞����h���f�T`�7����q'9���;C����ee�qA9����Yz>'�5�z7�Mu��dK9�^&���h�� �R��%����YW�}�`RcZ=��\��<�|�%�ͷlˏ�>��9�H���-s ���y���eV���8�Ү�~klzy��U��|���u�Q�\	8ȁ͹�s6S����}�Ư�W
�o��@x�[��=�! ������-��}�.�l�q{� X��� r�x�sYE1P�@EW�5��޶���ml�2^)��3�#?��m6nbz�{X�<7�Y{T�=�]>���GA��������2�Q����~K�:pt�Veɮ�M6��[�:-BSg��f+w��)X�b+���A����C�p<(;K��|���P^ _&0q.��u��� ��k��9��x� f��Ʀ<�m��-%�K�hK�sa=�.L����%�1{g����i�|� t��=�*Ϫ��{�Y	��V������k$��7gu�xTڪ���͵�,��l�����*�� �%�ZJ��+Zl��VT]�?���_�6��P���]w�5����}���Ӌ�0��fL��u_ޘ6�| "�X���2�< ��;�o�v��:2����/�O[��lz�k�iŒ�&((c~��H�f�d�Us��]�w,Q��^K��s���j�Eu0u�%�d�l*��H���Q9j%�={vT��_���� ����l �?�[�=��n
�t/r�Sײ�	���?��n�U�h�" ����8���PD��?�Ͱڊ��y�1T�a�4�r�8�c]���R�Z=�q�\� ��\(��{o�nY���%�u����k�<�|��ۢj��2�z�FV�b�TՉk�����Gl�J���u��.ohݟ�����ͷ\])�$��B��?�� [�+?n��Z����>�=ܵ�լRhyW6�s~<2�w\C�����D+8:�a(�.��0] jx4�.�t`�+��y��DD�c(�UA��.V�y��ц2��з�C�
�j��V�0�(o\!�#�O3��S�1����?���i��V��[�[+��<���>�ސ�8!{�e�hiٻY�Gخ����e�V	��,�뷖ߵ���s
��.p_��� $ �x��?VR]�y�К��؛�	s��,�e+�	�;�E䭏��*��F�q�0D_.#�]&c�w��T1�j�g�zy�ߗ�ؒ���t�Z�+�XU{=`}Ҵf�VV����3>;�䳾Z3^�w#pn���g~}$/ȗ9�R+�-i�;��m����eܲ��� �<�ǈ!�'�իU����Q�(3�2���.d,��@�a���D��p�@#�˾���P��f�i����6Hↅ�-���#�x��� ��ƽ����"��&k����vs�=�=$
��q��(Ӫ1����E �K/{Ư� �*�9�aśF�Fo>x:�S���J0�B�wl��i�
��뛁�vZ�0t&)��8��%Cڨ���`�g �02��%�&5+��,��7�H 4��ҨHĒ~y0+���'#\0�&
nQ���P�׎E��nB�t��O��
�ڕk�q�/�6e��GA�Z�1�VYFҮ�Ϙ�+cP\R~�?R�L�]*��;���rVΑ���ː-�����} ߙMc��k�ܰZJ������?�{�R�*%dM�3 �@�ϐU��H��gGԞ��jWY-�3��^�����G�0� oܸ���|������� S6����C$	�c��D��w��S��-A�u+>�>��Jy�?(�7^2~���|G���x�ό(�=L�z��nĠ=b��Ց� ������w���O�dO�z�`M�y��
H$���eN;��?��j ��	���_�����u��`V��8Dʩ�[mE�2�`:0#l�+��n��JSW,�~N8[@������c0�w��O{z�x\~`����O])��S�/KL/�f��9b��+tY�k�u,G�/9�d����U����Oe��Э�E�-Q c;g�Y��c���WpD(��O���k_�ov�l�V�WL'S���.i�ȿb����ō�Z��l�PM@>��� �����`�R=r���W��1�~d. �����R�x��q�.w p�;�?tM"0�L*M��أ|_��3��*!9�w�=.�A;�o����>�k#b�wU�q�]�v�����#�2�lehY���~x_�% z��>h��]�l+m���5Y�<�-B��"m"P1=�g�<})��� ����˖n�e���~ �k̾���������:�`4��[s|1L��ĨpYfʖ ��eo�Z�w3K�2��7hD���V^�R���:d�I��5b��̻�5�˕Y*!���ʒ=�i��hFq,E�D�nYt-����k� ���uB�W�.�vl��[c��տQ�푥��X��Z0�����z�;�$j��O�]A2C��p[�b=a�T�����k�AK.n�C�`�@�!�;a���p&�����	(�EZ�`X�-tO@^\=+P����m~��e��DL����*V�俣U֯e���3q~/W�A!K;��k�
g�ߴ�ì\���f����,�Q�zF���D@����0�z/���=-��j3S��nE�=�v��ϮP-��e�	HS����6J���0@ɭ��M-�
��3DZ`Ӏ�']v�2p���¯��y9��9�?����˿�ۂ�fn��B��q��z2F2Ɩ�uo����f��>m&b��"���Z2P��g���Ϟ�h��J�j��+��uw��y�땡�O#
���e�}Q�o�K�Q�蛕�芏-����*f7<!��S�){�lO	�2x�����l��%� {�c���A:�H%�3���'�����O����-��g�'`���W���!�A*�h,GW�	B=��b�:(&�$�F.r�����cl.#?�/ ��c�m~���Ϲ��������)5��"̞QdF�R�7�T=y�����3b:��uT�F��"�Zp�5��-��KE/�L�.��>(�h�;�v;����D��ݣ,�k�k�I��,����z�+Wګ&���sb6��G �����!�_Lf��h�_=�����a�`$����,)ю,����i/�f��+D� [��x_�1::ޜ���?�cL�0������7މ� c~Y��k#��ӎ�D�͉X�`PY3���\�~�>�\�����6˖تw{�E�����j7xU�J@"|X�����6�4�Y��
��-�W�b�U;y��8�J<�s�v6w��8��+a���x����X_�}��Ƿ+|�C�y��[���G)`5P�	 �zT>�`/���J�G?����@-�9G�S���_�,S���q�2K�`�e�.JG`�vT����#�̖[�gS3uD�����ۥJz�K�F�fc���f
^U��w�,�w�{)6�rcA��Q�k�ߚ���^Ո�{#��R<#�h�2a�A��db�s �; ]������w�=3-�h�kR�t1�l�� !��^���s�-�6K8c�M`�����p`�1�}r��ZM��W�Bנ�c)vk� ��KdJ=�Ϸ�`��Ϸ�7�s�������2ƒ#.#V�5T�ӥs~x�wz�um9�ߞn|?�(db�2A8J�@��oV��ZF=CC��_g)�7Q���\��V}3뛿��3Kg���ӑ�ZrЯg�#���,��8�aB�!{<� a)�$ ��v�Nj}3'�	��{ｳ;�_��_��Z��@�p�W���_���s�=�;�.YYa�����ܥKy+:���@-Y�Y@W�����'扖���m������=Y���;��
0C�8zG�������bܘ�`X��h%c�bZ�,����Iy���N���0"�����p �`��3��
��B8�1́�Z��k�7Z.VW�%�Q��g3q�i�|X��Ԕ���>��J�Z�P��ȽL���	��ۭQ����V|�ϭ⽲��=
�[�n4
l���Vq�_/W��k	�Vz��c��� �Y&L*� e������vY��l��\��O�z�fr"�Ǳ�.�3�\կw��S@z �}݀@[�I�د���=�(7喝�Z,[���1�2~H�(O�T������{�?K��Ū+K.{J0��K�I�/ĭ���"-Ъߺ��UAd��1��\�36��9�������;��*�S�?��"�ʛ�\�������g�D�U�j���b�0���_��G�>�>#�ܣ�f�1 ���A��<�I-ƅ�S�6�R��`�<�P?�Pi��B��6����2v�"��3�>h��ř�>b�~~�'��adX�3?��"#q�4n�rA�s,
��;��(Sq�. ]V�:,a|=ʔ�]�mL3�!/���=�����)4��d����̀��?����^����m�Ӛk-�7���ʃ���e��ٻ-�[��l��KQ��d}����������0a��$����x���+"� T|G��3���얠��n+����V99I���/J��-A��*��pwP���_0J>q�YaD~PG��r��k���%_�>���קk0X+O?Sj]�乌o��@U�^�+����q ���wWj	��ŔN�z����-Д�'c���am��a>L^=�5K�@��)�'ʈ)Ȣ���� 믃T�6�i��$��(!�X��C*�� ؅q�\ �L��@�<����U��d�޸��y��P�1U���� ���7۹/mf|<�c'Zt]�e�'���� �^�K�l��^>Uz��Fh���;�遟�*�*���ѯU��Yip�Z�F��y-�G�ջN�xi���߾�JK�e}�k��F��h�`�hS�MW���H&�\�76c���y��gg�+_�O~�{�ҔK�,��C�U鱉�~|��A|_F�Q�oDױ�*m���O��sYʦ86>W�7b�xx_U�R��RDv�#e�7�Ձe��7F <�+��*����� wD^��S&hz&^�k-�@�d1v~�O�s���ėMĦ#_U�Ǯ�篂K1�� Qv͊��`&ҁGO���w�X��#�/�7�Co�������4tB��9?�b�����,E-{��}���[�yk��k��;*lw�7=�\�Y$FB���Z}����'���xX������"�dJT&8�������]�h�ty�T�г�Umû�a���|>�*� ד���,�6�+�"w��׋��o�-�)�(�.^,���j��� �\t>��:��sp�`s����� =#0��˄�$6.���1|`t�,ӳqS2u!���X�be�����[ǟ�~�;|�8���_����2筿�e��ikf�g�<�׈�D�,��y�$e@wT����@f�×0�,�JI�\(�[����.� <z��~h�l �Ӹ81�W�0�ON��sLn�+��Ra�`@b*l,���|-V`�k�� j��a �@�"?�x�_�M�h���@nEQ�8b�/m�������&��3�����1�������w���E�i��o�����u�f2#yE���bt<8�����\f�6������XW�~��X�{�������zRO����3�9�[s'6�I����c~=N�������'���l��#W.�΍�C ���QN}�V9��<�����]�\� �ׂ[ooVH���yN�㸌����#�y6��{Z�}���b�����ƶq���j*'F,�O��eGwLg���JG������W��9��iV��1�x/�^=Ю��ǦEP j}W,�'/����o~���/�;M~i��󌮋��uחéD��T�<Z��$V`�Ά� f��O���B6�����	��h��Q�.�{�7CP;��]h� ƀ�Q��}RňG5�֜���(2��<�lpߕ�Vp����ZƔ)_��2Z�V��ҕ��S3������@yV�X>��w�EԖL��|�� ��X��F��(U������WsE�q�. �sx�x�#���k��L<���>�sO=���-�+��?+�4$�1�D����[��E�O���A1�`�v��W�ɬ]����S�����sjM~���y@�*q.gc=>���V������%~��zF���;�o���hX�ʼ+UB��[��W��FE�4�A
�!:�ȭ{�����$㏥��I󖶭M�h��#N+`��|���wX^�%/?�ȗ�=���]����3�Q�f�ճ��)#-���H����:L����[yޗ }�-��j��Λj>�߽��kh���A��!� Zf�:9ZϪ�񚃽��S�̧���5/�׳ўWC6��Xޖ`��==���|=��A� �'2�1
^{�:��h~��)��0U���X7���>�e�G!7|\3��uA2D!���@���X��.C���l���W���S21������Zl7_qp���:�X�ۅF�-esG�2N���I|'�%8��W�v�Kwl��Y-fQ��'@]"�3">C��1
�V�^ފ�c�C�e�E�j�/%r�-���{)�NlH�}17���S��1�aP�+G����6<]��J��`\��vɘl��p� ��NL32����_غ+Õ���b�N�A�*	K�[�W�7ޏ����ˬ%n��p��1�N�(�{��7�<�bcط���&.�fi�j���Vy������g�3�Mn��vO�Lı�t,R�4VmТ^�x�� �+���'�܏��/��<���adqL$3p��<��`���5�>_+y�]�+�=����M�rg���a`}^{{��"-�KqT�Sn e|�ߍƆ^y�2����;[p[���1*a��#��>�*f�Q2c9[¯���!ML .'�Ҫ������t��	``�1�XQE  v�R�/�f~vnQ��Jo�J�z�-URK����ڲd�%�}���Y�y��mD���/�{���=
r�{��\B>�#1�c3a�����?��V�[��w�� ����γ��o�%M�~�3�c��3U{e`;#?��p� �G�����]zp�2E%a������{�lX��>��7��QE,{6��8���`?����$nފ���nOT�b�h�{WcW8��>�Hc�Fp���U�Ji�QY����^�~�ג�Ց��p{�:t&�	oo<f fT{h��T�;����e&{ǁ)�����'ST��څ$JG�F��V�lc�z�gJ�l=E���ȭ�[�%�~�5FZy�����`PD،���5Z&o���h��j��k<ﴞ�(������v)�>6��>����4G���s�ʗ��Z���Z�7u�s�`~ci&]σ4�?tK�P����H=��&�����'?���r>�a�����ǡ5ަY^������GFu���Y\z�*3�10]Ǩy<"���ߋ"��X��W���
��2�f)���W��zf ;�U&ח��+���*�j~��#`=��p��>����AO2�î��r�~�,Z���J�'>#Q;�qK�r���ۏ�!N���b$\s_������!n���'
�5¢�3��܈���Rr%�Ä9p�e����W�۪�{u��dM�F�� k,s���ܹ�^,K��V��s䗬<bH!����1<�(��^��+?m����~p����}^d>�~d�泔ZO��?P��,��2��Zl�E^ŵ(��}\����dEv���&Jbj������xm&w�R���[���*ٲ����mڊg�堃���Ŗ��<DK�q����r�r#_���ϴ���e�KVFW���+��L�K1����L��> �g���>N��,Mk�@{���c�Ҩү&������t�����1��2W����P�)��
��F��"Ӫ�^C���*O�}���#?W��i£$���b,�](�<�+�O(k�����'6�����>0+6�d�>Q�o�*m~���:YI�;�_���ZR�X!E�ޖ�������|��������Y}n��f}�9�]Q�*�#�<�݌�sq�HK�f�ľ������֕��S�!���F��71�{y��[�^�}�ϫ��$��w��1Z�8�[�P��O����2;�a�[V}tp�q&ʬ���I��b�_�^YZ#4��8��g�2Wח�܃} �EMM��\O�7�e�[S�
���h�zח ��^d{��"��Y �tpUs�r-}B��PʘV�ٶ n6���\�ݱz�f���h�&5��}O��܋�����xm�����CT8�p�����G�E��f+<�Ň5\A��ǁ$
U��E��בz�d��8ӻ�k���-�I ���h����?���� W���&M���qaѩRX{��o0�}�jU�:���T�c�06̪�8EJ��ATe�y�x�>�m���kK�tj�Ǭ��6e;�EU>����@V�}����w�)�[(�k�A�Re�w|����:�=e/Kc�o��<_ޏ���dfu��y�L$�=�N��c�--#{~� ���W�\R��\��Y�T �bR����X��V	���u��������h���s�qV��|���k��k(뗖2T��l|��������|�In�Y/n��~E�k�7*�@��l1�ּ��*KS�����>6�a/k�α׷�WF(�;����r����S>����A�	�hP'*k.~z-p��"�gs�����=��3���{����|qEa�J�[p3+���ݺy���<����`�TX&Y�u4������y��� �}%��qۜ�j_6�^9�w���U	�C��9}���/u$^i�P��#�?�_����C�i�r���-G|��-���>�+~-��.2̇���z�l��({�a6K���(�s�����Y�z��)a��y�r�i�7�5�ӣ��{�l��e�n��0݌1�@�3�-�ѣ l!�j��^���} �*��~h��X�� A����g��H	�����M��N/�^���W���Z�D�_������d<2�ü�����|�t�r�����,1
J���@n�7�3���%�� p�7�7��|�#3 �T��a�ۡ/ \@��ղ~�C���J�����C'��{�1]�0�����_��_l>��Oo>������O}"&O��.���{������,�'�xb��J��J~=~����Y����2ues�O����M:(v �6���X��N՜]B��if.CU{VryT>�@l���ڠ���vu`�+?�u��w�E^6n��
qn[��k�(�b�ڮ�_˝�5��8��iV��[�x�2~��T�6ˣʿ����v��Z��w%�=�@h��Q�੨�}��(�|F&O���z�| lD,c�ShZ���ۚ=�ݮ
P�*@���An~Z�t�r��pI@qqK_�%
�`�>�~ҙ���-�Z���S�'�'[C}$�|~8Hp#���t�V1�;�S��}@���|�ie�Э�D.P�U�/~�O}�S3��hP�h��v��������:I�+m�S�r���[Ͻ��K��iGo�^���	Vi�D�u��w���r��:/)_&�[��(U
Ո`���zg�v��:��l��ȳ���ir�R "�%���������p<_Qt�Y� -�-G#i��}+?��9Y��Sꖖ9�s�&�e�"�^]�c�f�i�֏��)����Fx~������us��B�0jLK(�jo��7��ɾ3�YZ��x��+ǭy�Ď�bK�f��ߣ�.�K�q�=Zr[T��L��ڃ|U�!YT�dy��6L�1�qo�� ��:�7���q�Y���:c�O���ͧ?���_��_��f��.&"w1@��T���3�'�2r$�||媠<ne�U9Xغ�Y�����ُ��>{*p�ǸΕ�'��,���Z�/>�)뭹�F�+��*Q�r鿹6�U�<R�qr�����)
dT�+� � ���W�ր�P�x$�O����L%C��u���+{�DÄ���:}Wr��)cƌ�X�*fO�/�����V{��"�=�r�����ڜ>sz>B��>���xe�խ�W�ߧr�$t�+Tk�9��)1�j���|��l��I�}E%b��>s��V� ���z;c��Y�:em�y9���/Un�9ǭ�p~s�����O��l�=82T�BN)�X��o�7�\�<���$�����泟��ԥ\jE��I]S�@(r�=�E9|�E���pW^��]����f.�+��+�z@��Ǿp��e��v����SzDO������K��՘���N|%%�כ;�2�p���ϳ�JY�}��\�X�`�0�>��l�ٽ���(V�-�}���ꨘe��Ov=�BQr��}O���H��$��0���7lK�XS׊!diU¼w_�b
�"�KX"}`�Xz}�k�r1���z���1XM�����`"��ڡ�*!�+Z���5�6�dZ�[cH+�M��~������>�\Xj�Д/������{n����}}�\q���qoC�J�U�m&�������>7�[�;|H����/.��2��������[�)�Ɖ6�)m��K�~��_oݙb=3�m��!*`����	ޟ�*V�P�ܽ&_��(�8)���c�O��G�=IZ�{���ϴҌmU=�b�*��� �gռ���겋��hI��ly��蕡z�5N+���R,[�k`�)Yz��i	�yA{mXm�k�w(��f��;b<Ų�@�__
��xq�������-�|˼���t��z�E#�Tu�Z��[��������Nc,\�q.�~Q�� �G��2�V6@�(s]C�?�EQv*^��+�8'Q,���8�Z�!���x�ϫB�}��7�iC���?6P�ȟ���&��;[��-�z�>���H��2�:.W �駟�<���[���Ѣ���xE����]�e
�9.�G޷���*\Ʉ?���'�]+����}�2�HT��'�14n����F�4;�\V�}оArE=���p����s�k�?-*]ve#�vWZB#ef����e�5�� ]Jk �+�!!'=��x�Ҋ0�j�Z���XiYAb����P����D�%���|��	�0�{B� ��tp,�c�mj���}�DK
�K�@�,��Y��6HI{�-�]"��)9�\$oƽ覃���P�~�nE��lX5��AV[m*S�y�ˌ@�0^N�]e�L���e�8�3����q�G���e�\��Չg�����ʰ+L�'���8��&�,Ԕ�d����zٗ�2�h��9���]��Zٞ���m����Z�s�eƙ��C)�29*�1��Uǁ�.�>�7�FpI���g�w��5b�֜��n�� {���4��^�7{e�:7�&z�h�U�\�GK4����9��#;�'��kbQ��ڐ�ׂ�Jඞ��[@;
V>���X���P��بr=�]b��6�+J�7yxYDن�jVc"��[T�8al>����t�M[��V�lŁ���+	����Y��@P��@d)T�e���V�������@�@y?s%`����<�h�1}�0\Aq붏m��((��r���aF7
���y��])QN���"�������)?:�X���d��	�a��20�����.-_�#2�z/�����N%W��;�~0g3E��ŵ�E�ӈ�_B��������+>�[23�]�D�॥���=�,�h���P6)��]�_����%u���s��[�E#�k��2�" �"�ǋ`mٖR5�F�
����]�����F(9��-����q+�/(����Qi�d�m����jȟuEJ���[Yq�V+�-k��� (~ ��Y߀-����
��z�-�K[{; "��V�m嚠�e�"�/���n1F�R�?�O?��cvЫ�ԗ�7�7����V�.T_��",�z\Z���o��v,M�N��v IKI�ƒ��~ã�V����l,���gG�]h�����Kz�� �I��hw���G�">8��4?�H'�iE�ן��;+w�>żb���c�wQ�ZiGW�L�V8)SD�p���I]��Z��K��h��R��R�9����;>�����������5|� M	Y�?���'Gl�:6�ُ1���]������[�fK�����Q�o�o��8�w5�ը%��q �ս�V	�ȗ��T���1���
��t[N��t{7�[��f$�ĕ��ƽ��rjʟ���g�yf�|^>w��@�P|[���V��_��8���JKeQ/Y�_~��m?�ˏ�Ų�z��C��>@.�\I�O�f�r�L�4Y�U|�����m��Џ �vů��&?MNm�h2@�Vi=I�)�#`�(k��(K�s�+#�~�Ƹ>(���d��W1H3򵈕��F0U������z_�
h�׫w�͇6�"�D���g��ՎNK:bW��O�����oj1�0���;�V�2�P�~0D�(��;RG5�X�]&efe�/��TE����l����p�p$�k�F����t �d��t�\���l��J��7�=�>�~]�[>	4N���V���(%��|^~ݗ��Ք>BQ���g�����7�_�{�Z��9;
�7B�<*�����*:��n���k�Ge{�^�p�2+�LK<��3���@/Zp���G�_�V�&uD�׋ ,R�ކ[���_�i6�����Ey\AQ�J�����x���<�����@�˯��']ϧ'oNJQ��!k���n��l�f�z���XG_U�dx���v���K�VK�`�,��hQ��UeqY�J�H�3��0k������4F��RQK)M���%,d�B��h�5ί��Df����G�۪GX�\�ʗi�K�}�\����,]Z��~����������nz��}`Ŭ#9��j1�x�X�'1{@�Om����џ��~��:��;����?��f���>~l,m���$YL�>��������<f9���H�S`T�V��Gyd����sT�{����XoUg����W-�*����De&����!��(��td����{ԂQ!}��5w�lE �+($(z�[���b9�����ԍ ��I=}R`6�����AI���cğhQ�@�G>ŵV��{� ‸R(F�5��e�r�t��6�}�er~�28�������2��T��(vZ� �z6HG����PK�I�,H�I�○� 7n��ʴ�X�]�[���	͓&��ㆊ"ps_N�ӳ0u�eG�n�l#0��7so�)%c��@�5�L5N,e��ڇ/>ڑP]��O>���k+ ����������������G`����Dx}=n�HR�Dp������G?��\7=[�Â�c���ϟ���嫛�T���� ��0g�_e���@�ڕw}�D��Ao����0�<}��$�QQ̫�7�~o�9�3P�0�I���z��
�E0���GYa3�+_��O�2�Tr6�L&�1��rϻ��������!�uk���
�gm_V���DN2[�9��,���Ә�,���q��PO����.�!k$�-����DXE�8��)k�E :�f��O��K?� ���8���{=�s0���֒2A�]�]�.XZ;�L0����KB��k�E�b	�ە`�"'`)+�b-��������@����dk����}�m�N"�p���u4��ʾڂ�ǆ��6��V��"�	%]S�ljt7��~&����Ey8Å���9	M�7�w��7�Q*h>�X� "	�,z&��������JeȈg��kw��	x�=b~=>��H��F)�6�O"NsU���⹽ ��D-�R:	�|=���aN�����=��Ņ��㎭%�-��m+��M��o��z�R�����]��3��:`����/ VCʼ���F���������h��%?d��J;������t��Z��y d��!$�W�&�m�5��n���ra�*R÷����n	�Oo�ڋX�JWu{�W/m6?�ICs�h��u�>mE�	�d���
��J�`�[��=~�u���<`O�ƿ�/�7g�od|�
�z u�7�Q�c ��ֶ���2��7�+�AVF}�e@����`�~U;V2�'{�4����#|���w���4bzY�e�K֑��V��z�W��X�أe��q�e����:Qi�դEI�hÙo��G;�٘��*О�`�:v���O-AZ6޳�1B��R���l��G{pY^���K�G����3+!e�<q���׽��̄��l�0t�O1�.�(�SF6R��T�R.��u����m��܅�*�>��@����,{��7���9b�ʢ<4������%��o�T:r�P]�.��g��o6k1��s�K��s��Lܧ��3�SD�����7n� ��3[����Ҍ�r�]��X�5���IȻ%�g$-oo�l5fy-!��V9��JR&�P��H�1��V@+e�2yz��n�N��-�|3YX�CL#�Q&�=�Ѱ�#Tͯc=�:�����N�}֣5�3��֢d9�^�*3�IHy�T�(k	�z�T`��d�g;�!צ�܇P ��d�4kO�'{�L�zL=
��~쇸�52+�%<��ᔪS������'�گ1}�#�jk;�_�ds��%�������*홵�׋|�5/� ���3��`N��P���}o����-�d�-�] � ������|������B�i�+H��MH��+u���%��PPVW��:�W�o���w�!�,H%�*�u-��������W���w|7.��x�ּ����v�
��`�>|�8����QT֣b�����#�7v#،���V�[�=R,g�oO^fif��I�^}p3�QM�}T��@�j�zd��&�IP�����{���=��.��<3:~��hB�ʯ�׃�l�r� �7��LX+�9�s�㛵�������+��b;�g<o�7Y`��]8asp�`s�[�ˀ�)� Q���s��}U�Wuk"D{�׋�������
t�<�Zb2b�9�Ae!vW]�wA���w���U�a�PS]c3\f��Z�wY{���e��9�y\�x 7"ށ���I��hH��%���_�2x�e��z
�>�2F"��g`Ȁ��C-��(6�2�GqN��i6�F�Vш2U\zi�����G :�Mf'�Գʼ��E�Pf)XJK�A����5�/%=�ۛo��I�u��
 �4�}��Ȅ[��^o��Ppu�� l�pkF� ,��k�&A�P}��0��!΃C ���p~sp�A)8�]��D���W�?���f��HX . �H%�Ƣ��paaYW�\�#޵,θ#��zG�飈r�xꩧ�߄J�+L� �	�ز�?�4�̩�?�g"��v�������L	����xn=�����w!���_x���A���\��sf������������
��3Z�V�3cev��樁#�c�dЉ��A�cr�$U[��L0���\�Z��[ڎ �L"(�r��bA�hߌIF༤<=��T��u&�@�~�n���?n�p@��C�7��2y% �~i�u&L��,?�>�����:��$OǏ�͖3i!�]	�6sŃ>Ap���r�i�6:ޝ�+/[�l�K�Z�Xe���/W$}p���	f�8�n3�hD� �.Z�l���h n="CN��_�M���|���^�[e���ʟ;�hƴw��-����	e����>��Xƍ����1>�[l�Q��MZJ_��8���J�4zs#�u�.cZcx�:���[�]��(�6�&�(�];Ȱ��}	�*�1H0�;�|t?��	Bo��n�0������ ��n�>m���u�Sޏ�ۜw�8��m���٪CV�������p;}��g�@x�#ۗ���L���~"\�ľy��� � Ym9���#U����q ��(�F'��)����o='P+7�mB��s߀W���G���x���.ކ�K�]��w�O�������%���{���_fT�
��A����b5�s�xF�TO.Tc5���>�.�S�FK~W���7��<*�~=�1N>^ϨL���I��� �:ӈV�MUZ�V���5� &"K��>S�"=�1��^6Q{u���P���x� �Lr��D��N�<|70�Y�_�vt��5��y^qGqV67#��������(U�'����� (�������e,g���oW�uY�}�܁BT6T[-�#�e%Ն36kF?�]�8�1�5�eu �T����lT��*����@YD���(���|�������U��xܗ,�)[К�v�/K��x��~g`tmf���}n��B��,eV�J���} ���+��7�����VzQ�x��@��ǘ�75�zK�y�; +�-�&j��2�LK���/�a	c��O 0ű�-��yU�y�.Uz-Z3&2��\=?�W����Lh_��V�ށo봩��c�q�T�������R�����@~{0���m�:�(��} ��=�
�ec����*��DB��f���'�:NW���Z�Ǫ����IVc\D���GB��KP����+Ƭ(\���t��/�Q�'�������֎�*�xm�����F�}
��ܶ���_V�%m�%��A�RF�q�@7ʅl�e��1��X���^�,"ś܊�4 ��vM3L��FuF�QUe��g�g$/�5�?��>~�������������E�������S6`�ЌW-�,��˭�U�X��~�WK|�~s%���,���y�M�Ɇ�v7��g����쨈�\k�S6Cm�=��+�Ȉ'"##77�xÜ3�eu����-y~��|�]����^�(�*0��E�(�:`݂��Wv�@�ř`����*��ҿ�v�
�%
������$~S���Ǔ�-���_���0>"�&�K�Y���s<������o�|����Yˋ��Xy��\觩����]���}� ��A|l�?��Ћc�W�K1W����YB��Fb�5 �E-p��l���1R��9#FE����Fy�]�F�f�NDJ<"$��!��*��תG� �ds��]
�[���e:�*��7kqNVW��l�tpFK@w�^�o n��"Xk�����	zh���a��c{F�v(��%X;��xӍ�4E�7zbn�9.���w߽e�x���T���=-ES��3UxnO/ˏ�� �pyEDx��3��GY@π�_O���Z����
 G!�Rł����#��HC���k� �8Z�2�&�I�͖>�"�Q��N�ӂ��:^
[�=:��|�����<����3W� I?��>5c�Q��g�k#ȥ_	���w�G�h��R�ɧ5ze�ƹ�q��s6+k��Q&7|U��o��mK�>�o����<�m��GY�s%?����nTd����[�j��t\OW����H�4�Z%�a��(�]R��������,���|��'H|R�ٷ��\���o �m��+�I����i�����^���N 燥�(�f6���\SH���o��N��v# �bUQ8Uϭ(ޓ	����>)Ub��@�<G\�P���� �7���"�y�������2(ہ���#���kL�{%�<����kU�oxat��>��ey�c��zQ�cV�C�b���}˭@S�ܵ:%����{�|fç����خk�(���Xk�I�@���2(3#�U~,{���Kl{&�c}{��w�����d�Wu¾t!�M��d[Գ�+���Uތ�s�2{uv�������N��<��ͬ�}(�C6�#@9�3G�����'�Q����/[; �|� ,SU�3C%���J�9Љu����X���������c�D�K�gR�����"G�+W�, ��{饗�� P�D� �\�p�R$��g�Qd}V�A�8�~���6��[�^��x�D�z�Y��R�ߵ��)�k��YF���x��� u�;ذ�'�Ze��*�#�d�6���㵙����ҥ��9�+#�kU���������-'U�stDb^��7S��B�U��>�(��Qat(�u(��D-��*���gva�l����F�
l`�y<j1�j,��hgŃ'�B�'d[c����X�N)��b��+[ƭ�}�=���}�L��3(�C��xH���7}�w܏����W�U+ʄ����@��s��+���M=}s� �bP��B ����<�ЂG��K����^�(���T)�L�kIl�UٔAօȻ��n�Qn��>��}��������� ̾���k�	ϒ
����p��y�<ʞ����6e�2�"���-r~��,ޟ��k��W�]��1��(ex� ����V���bʉ}�5����U����~˘t�q������3,�J�i#����z,� �|��<��+�&�vh����?bX�o*F�h���LyE�s  ������^�|�1V{/�9+;$@�A����y��l��p�q�/���擟�����i�}�Y,�͗"�?�O��-��M�׏XV~ K�kq���NL��F����7s�qt5����|��}Ü�����E���\w���k惏�I[�W�>'3�>T����H}��kx�WM0tă���G��C��@�ώu���?/ǲ}ZG"��Z�s#���WN��L�Vu�|���\�b�V�
l�9�=c.^َ��U���8X]bq]o�����k'_�<���"��k9ؽ7�d	hX�Yn�^]�+��OG����R��S8��/}�6��\��9��S���L���rcrB�fx�BPb[* �e�5R�?��O7�<��ld��}�s��ɢ�2�#�YBm>Ӝa���"�yf��U�N&���?>�py��z9�-z�3�p�8Ƕe|���:y=ƜWs^��!An�ߧ��2��{�*��#ߏ��Ǟ�u�O���ͩ��9U�Z�%kx�/O��Q]2��*G����M�nf	G�4����r�i�1{�>�M��n�PK��h	x���)�
�c��Û����7�w�R�)ԥFJe�z�#<�w~ͼ�\W\~�|�x�<$!��?��+ڛ{L/��<˔��c���Z!(�S�]�`?�Q$O�%�+��/�0��|����j����*�9z.��rp� .�/Ƙ�$�?��s���<��.�L���/�u&J�X"�k{�ח�yj0���ן�c�{F�!�e0�������ȓ���#c+bS'f�?M�x��z~%7��Z�T�� ݈iDe��5F��m�N#�H��=D��n���x��ߢ�`T��2[�9"�R���*�%��3���kգzvR����XX�,b�KYI������H�T�Ȥ�(���HʯxO�g+�?�b��?'�� ;,�yU��Y�%Fs�*0���b_�tKIy=���J/#=�XoyK[��8u���V2��n|��������*fV�Q\yr�7��Gv<���?p��)"��y�5ޱ��W~� ��6�)�A��g��j?����2v��*�9�yJ�M�?����c�|��FU_R�aD��+�5H�{Z2�WfX������k��'+���̌�(�az����D�#�]�4^�mQ�E=Ta��/�sG���2�����r[���\�-��}e��ӣ���f@��T1��?��+��թա-�S}�*�G=F��(+i>:�G��"����%���2�,v�[)q�L����&��uƃ�	��Q}�ƿ%�F��������}�˴x�ܳ��'�e6w+���u�rz`�5���y}h���U���T=� ��	�*U
7ndj���N��\���U�=�ܳ��;�k(���ϋ��ͳ$l�j�\;�� ���L���0T?�^{����˳#�d��dgF����5>���}�G�	<������vE�J6����6Jq~��-�7��%ƾc���ٺ��	K8��e����⏖�e��U�L'�P��-�4�������X��Qh��x}�(c�ㆈ�8�{)�Ǹ�}��5�LKh���@�*�'\[�J�ؙ����=[����GĮjy�DR`�F�^����xo8{��Q�zU�ϋ�b�-/��Y�4D��­w@E�K���WB������q�L�@ܬȵ�!"�qp�>�#�:�I��j�R|�V/��?��l�Q�O�+�=�@��Ov�Y�'�Fȃ{�]w�q������
�7D:1�칼 ;���?�w窧A�<��`��%C8	+�OO��
���K�;t[b��.i�ύ>7�}u	'F�Ǎ�S�JN�1���g��:D}sc&Ҿ�:ӏs�����/����o�Bxx6����feD�C�z�z_��?�n�`T}����_�[e@��%[�E��ǐ�0)�3�����e�VF�l�~=������ܛQ��z� �p�G���������J�U������'��G=#��xlv�{x+�Zkx�C8�Z W�W6H�ˀ#V M��<L!�	������-����+^Rx§?����,���� K��Lׂܸ)p��lv�V������Uo���������:e�D>w2,��=���2.ČB�l�:gM?U�v�~p9PɲXW_m����C�����U]2���8$H��H�Z؉�V�(x�Y���}|�wgFu��% �j���/����V@��F�B�7����������2�B=@�4��x�g}gFGT�}ːh��'������p ��,U��R cG_�� ���y{��;�}��CBK���X�gCU�ǐ�[,ۓ�6�O��q�����*5��~��m�Η������y=S�q C�e����d���l��\�~ 1�j�<����g�x���s��1���R�K�CjTV4L0H ��4vC�A��������qLM�O�96�F����~��h4������k���C�xݪ^����#����YZ���=�:OҐ���E�碘*��
�V  Q��z����H#�f�_k�r�{�Xҏ����g(3L��[u�֖��x�S( �q����� ֶ��J%X�vf�x��2OAIUv�p����u��S��8`CG<5n�\�����Z�/�Ó�
p"8I�%�l\�;�	�
�z����~p��q�i|(������k<H�$o.K�~�S8�#�`�����Ǯk�,<ɺGuT*2�-pK�j�E�\�!�Z��}�N�&�~x:�5���>�c���P�ۥ:,����FH��# u��-�g0�	+rS��(�����#YY#�9�����5^;R�?��8�y u[��Z�tHrL}���l���oq�J��#��zVf��7R��]k {�ޯe��
[�DY�k�e��Z@��^X��j�O���ڜ9{f�h�V����K�s�R�O@͔���
�_�E�����3���:P�4H-��x=[���>}�|2�pFyύ&&�ج�({pP�Z����jB�tVGK���?�� <�{�s*1Ճ�S��V/��_��7��4���r/�RՁx\\�?��B�������?q,3��E*)@5��X�%&�O������������`������'��F��³���F(�#�����]�A>���9Вo�6dz~�~�ڙ}yVϐ��D�<kL�7�l��L��r*PL���@�'k�{F# w��-&}ơ�Z��c|g��� '��lIQq�� ��\� ��<(����?�_<�s��h�Q�{�T#P�� �g�o�CV�aT�P�����Y]�^q�[1���%� ?���"���9֫�_�g/`(�8W�%) �� �9�������x�c_�\r�~�*0������&o�<ʪ�2*�U�~�V#Z�ͳ�JG��	��� ]���zR`�z���6��K�t����(�lU��8eƦ��%/�}�g�WB��o<'{fl[�2.ⳳ6�C>����A@UP�ߪ�=�w��;#�{�f�>~]�b=�7�b��+sͳ�޽Ȯ�n�DFP_M�
H���U�̞׻�<Q`����M7޴=B���Q��UL���zFC�z�,�S%�F(+�G[�eb�A�>��@��1�ɭ[Tr�������O-���_4�l�ʶ'��2<=Ul�����NR�Z�xT����ys�J�{���i��֠�V{��e<tq؄n����r��_��\?r�
��Gj&��d!$�3����_�s<��_�̮�"׭=c�������Y�s����]����s���ȎŎu\S�LnFy~�X�L���6ʯ��'T��r����=�i������׭{Gǹ��y^K��ێw����5�b[VL�v��y��Ԫo����j	�caD eL��|�����3q2f�̄Z�?(Yٹ��\�����7�|薭R$�ˁK�G�T��ɀ�ߗ�k��C�B�c.����m�+W�wϷ�׋i��`|��s���O�������Q������`����o��]	�%���q/��g��ꫳW9spu@ħ>���4ZVg	��� ��W1�"�ݣ�Z����fϡ��D X�@+�!z�� f��b���~D�F��8q����.>{	���ш��:�#��3R�L���Kx6�o|�L	�B<ӆ{ӽ�=f2k��@e�{4�l���S�e�\gduɞ���׵����b�xM�G�s��lw�x*�'�ݢ��xn+7��_�ۛ-�תt�̵��*p�uv6��L���72�载{A=�Ӣ��λ��������K�����5nb�=Q���A����˄L��ƗnbF�g�ƶ��6��1��>�ꧾe�П�w�^#s�5'[��JL�QN��d.�+ �x]�W}��To����W��!�^�`���o�}�a�� �%���SL��Qy:B��կ~u�®�5�k��zT���:������A�Z��@�G��-Y�^P%���i� �3����'�ם�Z|��.-9ￏ�ǥ�;_g� +�5/c���#e{=�{+�ժ�R����8�;Ty�5�o�X͞Y�wH�V��{=�=�#��,�D9���d���b�R�dm�����(�}�$� >�ty�D�Z_J��"����{�Z��- ����lߠ� �,}���� �jW&Ыk*r~�>%����ڼ���W��	L^YŨ�K�0�m�|�U������@�Y&�o�<F�]�9N���V W�fN��&r�/~0I�����z���!tAV�Q���%}tÄ�!�6�s#��c����d�^ >�؞�V�[Fz|��V �r8����,�L��~�mp��T���W�-�n��1>�Q�NY�XV��R�]}>iK����h3k5����Ъ�������J�X�Yޔ���F�#��O_�xb�^oC�����y{}�i���:�����"��Dlc���z����
~�1�.��ip"�ߍ���/k�_��c��*��� B��������Zr��;��8_�S}/p��s�M7o���{��g�Y���2��	�Mgl��iz|L�1�xU��	�7Ǳ���pn�RW���*���aR=��\��>j8�@C��>K�Dhq�s�'P��>w����^�F����Y��u��χ����KU�O�f�~��H������}��P�]��e�\�
 � ��cr���<&��hĊ�>�Pf���� ����  ��܌z^�%�`�=0҇�98s ϵ�?	�͆,�����1�W�=>��^S1��G�*S��(��RElBT���K�� p���?����[�9���1�~�����+�~�F$+n�c�E��k�� p��7�<�
��㊆?'����:-ޮ�_u}vm���9��W�r��0n`�k3��3[�;	z��늗�ͯ���\��'+�����ˈ|/�S�7���F@���Zm��߷�.��rϔyF-F���k$<��ɕHX��|�Q<!��W&xF��R�¡�n���s�$Zw��̛K=z�pi۲����0|��
xr0�d��cVHO'/���~���G9�.��̘��'���zi��?��?6?�я��Ծ/����c��R4#�2���k�G!��%
���&<&tiF�jT��FuQ��։�|�-�ޫ[U�5�n�{���0x0��H�6/#��z�k���K�u'M�ml9gbV��*cf��P��+���z��A��ތ��*�}^#,I���CO���~j=�U��>�MQR�~4)�\  7�E�M�LPDK�'t"��}Ǩn� �#�Q�z/��u��M��y_Z�4{_����>K��ٵ��} �Y .+�J�-�����F�g��}����;zAZJ-�%�. �� /�BT��r��T��0�xl���:�6fT��'γ�XM�+@��
� �'O�o{��*#����s�����?$U d��/���V�q^�������b�☜�^��������pO�]�ql3�֪���� ��Jpd�m��NΨg�T��+�hu/"��3!�%���~_S�l��o����VZO��4,z��J�W���R�R|Z��u����W�����f%$[}��@�R=�$H*�KT������%g}ǽ�l	���g��{���{{s�6��Q�+e6]�<���f*_��U�Y��*Ϧ�$GC �����[22h�8(u��ct �|�#��m4H�E���P �����w�*��[��D���O6FDy��A?9H�r�+)�b��w+�&���ԣԎ���]KGq�h=ze�膬/"�1�����{�O�G�O�~������=��K�K������3�}=l�=���Ɍ�1e���:IZp+�*����&i�7�}v�n��g��CV~E�Q[�22��0ْ{F���қ��O-�A@�p�?]�{�Z������u��}ճ��Q�Ev,_�|8|':�����λ��|c�?'z�G�%�t��P��Xގ��g��es��E @"���S�O8��p6���M<���u)U��h,�e�����s�=7�C`��ە�9�#��j��s��\�
U�צ1�@>]������m�:x\�_�c%F߱��&���L�v ^eS聥%������V2Pأ5�6R���襏=�pK�S�V�Y�o[�ǹ?"�{s,�I��\��ŏ�:�*#���XW���������(n
��t�Mf�V�ef����F �<'�k�w��ZRm��b���<�W��YF�-��u�䒏Q@O�oV��������,s�Q�� bS�h_�'�©͵�����g 53Rc�c��Q��3Z��o���e`d�㕉���U� )qe	�J��jc�^���/�)�˗��!{���8ks�^��*[�҆�'�xb>��z��Q0�}���y��/N�f�����V���Ó�<�֩�;<6߳����h ��Ȫ(z	���y�w�}(j�#�x�ـ��_Q6���#�=Yf��Q�o�L��X��9^�/��������*���2�z�q_�*3��*�����Z�Ȁ��τq�L� �U#��a���?� S������c&���Z���Jэb�7b��sƃ�{Q܋��/�S�e�X?�̵�bb�Kh���� ݛȒ=sK�	=`�� ����i�\y=u����>;��Pyv�}���S������9ho���mL��E�|���W%�F�
���xOv-|�<ƭ���}����}��5�6�P�k6�m�7��Q��=�S���U��{���h -�q��HL}Eԕ~&܉�8$���N-c�j�U�WS��-C�jo�nU��崉�����3ZZ�+�v��S#�dI6w���J���x����Y��ظ�!�gD:$��&Xֱ�����}��'�<�߼ ��N̖��k�~'���!a����FU����(���?�g���j�]p)�u1�:���K�^�qG��z��4��jy�F����A�&,`�������-�������S:FW�V�U�D������}����
�\�A�@q�����闖��G��<��2"(pc ��r���9�8�GF1u����f0~y2޽W��q�켚q��q�7��24��g5�3ّ��jOEO���)��7z�	���&NBIȁ,�6�.���1�^��[1�6��z��Q�'�qQ�]r>̀�r�F�Ruo�]��.�D{{p�D"�+S�K*}(f��JHe�1j�9��_��lZB��h�����>u�NW$����V�D�3[�cGA.�[ףh"��:WKz�=�E�Z)�b=�>\cȬ�� qʌK^�ޤ��"�$���	�U聀(��"�WV���q��1=�@J2@0����K��'�'��Ejk���@%P+Э�e���;�4f��d�{q3�����=r�N{��=>�S�y���R��~��nɈJ�eϮ�^�[�g@��<�wp���y��S���|p��D~T`~t�p6�[U�8[K=+b�5�/�Y-���2\T��И�ҟ� �+S��{��L��>/v�D�}W1��g�&�Ȕ�k���^;�Zy�����վ�y#�_r���7<�ڐ	�LHg�Ї����J�U�LP�!�P��������׳�Eߢ^_F������"ƫ�]���ܵ FR�����N�3����������o�_��W��~��y<3�M\���^��
�ʛ�L:�W��� ,nT
����JfT ����0�Ł,�D0��h|vkn/�ǙA�3���c�yU:���3+C�卾�8v�F�� e�~_l����?`�Um����_�<S�s  ��IDAT��Hk���u�P�I�S6nq�.ۭ0�JVx�Z��C�=�YJ��q2f ���*%�L��c|G����ٵ��I�k)��g�[�R^k�o)�e�_O9d�A~N�g)8�OK��?k�I �X7Q��+�Y��O;�+�	��/Z�;؈�"��^�02����(^N�?��z�+t� ��'�̊��GV�P���+ ��8@X�;n�c{,.m�$�A$o�V���˱��Ц�l��̗�~!�� ]��/��/7����y�sz==�k	�����=Y֒5�k�>�E&ӂ�4�G����~j����2F��8U�M�f�jˈq=��X���V�U���F�M����7"Ӳ�-:�|��mͣ�8E�h&�����z����Q�P�k���E 7�"�ܓ1|OHTB�u_�o��[u��Wl[���~������1B@���$��7�\� %�̓�d�f�1�QH�}6O"���'(�ɦ0��n����P �!�Ǎj�o+jջ彍}��p�����?,�*N���_�c��-`�/�%���M�SY���r����w�\R�y�����U� 7P�L]�r�����fX�������u��^���j��7���ͽ_�w�숏�����M�?����]B������A)`ʳb0��z�$l�c>D^|�ޣ`�﩮���(U�v�2Y�"��W�2�6Z�
Tf����L����U���q��ؿk�O4
�;��d�v���^����Ⳣ~���zpF�N�YI��G@�����c%�ܺ8��Q}��z,+��U�(>���#�3�U%|2Z"TG���Ϥ��%����~��eK�f�K�L���.�_9�9�[��G����X\�͋��n|�1��\_���!j�bXr��?x=Ârh�r��1 �3�ӳLgp�����Zϑyy}��5j���r�"�����	m�
K��׿����{�@�Ta1���
8�UU��˫,�ArB
"es�珇��{_����+�^��Ĉ��W|3J�\_zM.3�ߢ��k�m\a�����^��T��j�!.g��d<W�۪OZ����r�<iJ�}H��z���[�����mU�*�g8_,��V���F%쪉.ro ��I�խU�Ϋz�N�����g	���|�P�N�_������V��A뻬?z��&]�����������G�z�UQ�E@!ǘӌ�9���Yzo�'�WO+�@�v�2>� Z��"�K9q8h����򗿜��
;�5�����<�������*����GV��S[y���/y�X&p�g:ˁˊ�>�j�g
Ԫ���#l��ec���{��ruq�8�u��+ߌ�˞��'��,)���}�0Y���r�U� ~cP��8},�z�����]s�gun��%T�W�29��3��zN�f�]���S�/���j�-�dVUp��ˌL���{��@s�@�um]�<ս��o�����n�U�tT���k���8^�$��2#��vĨ�c��U;��	o?
"n���ͩ`�@W�|*�s���c���y��VB�jK�e�A"�X�I�1�<�y,n*c�~-��3����sR�Ǎ
�귟���s�+�9�>�Mq�������aA���~m:Ӧ6�K�e����u�@�6��.:IM��,\������[�Q��\m�өk����N����g���i�� �Ӟ���(*C7�Qψ1r�����Z����cQo�kZ@�����~����;���۬:���vecݓe��%�Ɩ��^?W��LF�x<���̵���V�dV	��eD����j�[�V����}��U��}Z���zI}3�j1�>�<4Q�f9G�K���?����Z�l�����U�ᕜ����z� U�1 �lQf\��3�Zڍmh�C˘�������������#�t����8�gV�L-��6���o����W�������I���+� ���s�L��2;P�]m�Sj36��|?�BD��[�M�^^�^xa���/ϧ����,��O�e`��^q3����s~�,!YG TFz��R#7��̖L�3��eͨ�HVvզֲ:�]%+��LǬ� n�q|ˮ�n����j�ިl;�z�܌u����'I� n��}��H˘'����ee��c�P����%���� k���wE���������M�p}�&H�듰֣ ��#` �;{�N����T@�/�	����yI*`�kG%�Z�-P�/�&y)��0Q�q�G��^Vm��W��_�����*�Oxb�I������S�VuQ�J�0$�T3#pԴ�XW;�iM����~��W��W}�g�������x���9V�2mxS�To�r��F��y��[�U��K�Ɓ���v��w稘�2]��_K�*/�P�*=Yo��?Wc��#�>#��}�T�V�ү�׷h->�}N���7ʵ
��'�/��3�����'M�=�#VP�c-)'S���{+%���-���*p��V�	@G�/Uc^��z���:Gz�5#� �D���D�R�1 C�_�9Fc{G��QjK�I�����}sm'[ �0��W��?{�g�g�{v���p��O�1�����^N�8f\���~��3X�(����#�`��8j �bw����>�2h�H��@��?��g��3(3�5^.{yU1��R����nLc�0d�#S�Uz��(�����zed�&|�[/��2���X~r�̃)�r�^U�L&?ZeW׵�u���kV/���������2bz�CHb��xOJw�hu��ӈr� H�yZ�f�>���`d�6���i�d�%��u��y��ڂ"�@ V���г�30��WY���^;��Ur|F5��(�F4?bS�^��G<�F���y�=���O}ؤh����8� �Z��P�޿}o�����[yA16��LNW����xU]'/� *a~:Y�,����gf@��o�3=?�IO�f������V W�\]+���N(C�@�r��;�e�W�+S�n�7w��w��U]S�_c�yj���x?g|S�ج�>/}�"��U]E� �e���e���䘷����k~��bք�7����53�=��=�O.s��!��'����¨[C%�m��J)��BTX�әʿoQ�}�QbZ��&nV�(�ĺ�Z��~�c��y�I^���UFՎ8���X�J�dB5�U[*�ǵ�-52�[���j���rf����:nK�}��MY�]�Um��_��/����d�/�y��W�(NU��$��[��>%�0��*�}��6?���6yq]&%�*��'U��� ,�Q�"�z��a( ���sώ��.�_9> "�Sܭ �3O?3�[��0�y)�N#�xl�Vi������P�>�`yTg|��ln{`�${%w��D�*/��N���	�y�g�yDw�K�l������q�� `�������ȁL>Ƹw��ge�����H"7pE�$���u��T�ek����[���qȃ�#�ʮ�4"FA"�f��w��xUDR\�s��!,!�lbWT�/�=k[UN��p�[��kGx"�W�Q���x3*�Q��W�ӊo[��"��pN"���LƎ�X]Ǧ"��m)�^_�ڜج/��-e\��}���>*^T ��`�U\Fh�����;����Ϳ��n��Ƶh`A�����3�l�ֳ��7�����|�����"�{�K�ܣ�hu"�>����=���L@�?���Ǐ�x�B���1.Kzc���J�'[�Ί���e(� �����4݉����jND�[�a��G)�o��2�3�|ת[����Ⱦ�g��u�ތ�&��K�[�����e��9�e�/_I� �f�7ks�����.�A�%:����ߣ���k���V�U�[Ѫ�j� �V��׶(
ڌ!Db �[�t=6��z��j:��-��o-`��^F�TZuu�k��D|f��:F��������Uu�����
�W��=}��%<��R�
��W�/�W�jc֖��#�so&��𮏁�f��-M�KQ4����2�s��[=�<q�F1<����;�+�H�\m֢]��sϜဍ`�\=��U���k{����� <��JM}��t����h��}o���m����2X�}wy��,����}6W�� y@�����٢��+~��CQ�gc�"xɖ��rZώ��V�&>��Kd�R�תg���V��7��c�y�(�^}#N�����i���"CO�mw9��U<��h���54p[���F��ʬ��3��2cɐ���cLxu�9P�n-{9��BǕ��!.md��ұ�@f|�^"{˨ `Vת����x� �(z�+e����	E҄9X]�dsʯ�xE?��=�KhD9V��ȫ�a�u�lpڈ�u�K{�2r�_���>����V���*O�pn3�E_J�轼�Z��3D�:]L@WeK�����b�co'r'Wр�(KuS�t�R���O=���?���y��l���i��f�&p���2G`6���X��{qc|��d��7n��~�(Cޯѧ������㰳�Y�U�v������"����)�c\�/Ye���"^��V�ɌW[�X�
[q��"���k�	��D�%����{p��2^v_�B�	�j�rq`�ƩB�,��E�q��9�t ጌ`u�KT�z��|o�1���[nd�ZEkr
,.��z>�3*���b��>ˮ��#����=o(���cK�W���Z�5�����f
��/�>����U���y:�����^�^K����?���_��_f����e�8�V S�p&��U\���{�Ce�I�z��A,�%M���e���� p������Ϳ�ۿΛ�T���1b߷6����W.�2%����j�Z4��Y=���.��r�\��&�5 �����F�;�����9����ɍ�h��PĪ>7��w��Je ��?g�&���G�ݚ/Ѩc3�den9������ӕl;�%
o_�� �B�-�Z��T�{r��?��ƅam^ ��7b8S;��8�jCYKFƌ�g}�e���3{މ�"� G��H�=ʔTt���rF<���2ł�D�#I���J�G�������m:�&��X�wk�  �w�s5�U�͠���͛o���xF{��`*�V���X%p��ݫ��Vch������p��0�I���X We�8]}&d�z�P2Q6��l�37�#m�S|�O<�y��'fp+��AȪjSM\���03����p��.W6W��/��郬��>���\�Xu�w�E� 4
�F��L&KF��%���/�����2�N�������C���>���0��9���|3pt\8��e�,�)��{�o����b�,R�[b��1�F��X�����e9C-Ul��q�a��%�7��ޞ���L�����&	fy#�ߥȩB�@z�nig�*}G��b�.a��1>�P�Q���2�T>K(/����sVQK�D��ߙ�9����%�l�Ao����޽t�o���ڕ��X�h�U}1
*����_�bN�%�(A,�J��^	eyV��V�N񶊓U.B�P�����`�~�Ձ���+%��;����n��[���U�L��56���(�B���UH�K/�4���c�R���8g�ĕw�����Y7F����o�_k���7���]�<?������\��ݣQp�DOg����~�=۟ѫw�[u_R���d�̖��޻w4��ga�^IByN�H+����aK��r��(�܃��?۸�1�S4{ԓ{�T�����3n��0�S�e�u��=][ `K�8��+�C~H��郳�Eqy8ƀ)M�2H� �]�z����[bD� ޟ���th:*x�P��
ش���_��v�ß���l<O|�������ww�
A�<����/������`D=��U�ؾ�����5�4�
�l j�0�C*o������GU W ��h�K�����J��w1~��ꤘ\B���O}j��N-��*�����(���[o�c�X`������.�Yl��G��2y������߂���+��>Q�i2��?��S�Y�1�D���{{��w�yw��m�˒�|���H���lQv���Z^���tˉ1R^,�*�Eq^W���f����O�H4>�3��z��mVS� ���F�;ȼ.��D�,w���ƛW��/_�������o���\��q���n���[2��u���^{�[SC/x��j�@��5�\�;���V���1.g&!t�ؕ��G@�7Ê�"��-#H�Ap�Ǔs,-�Ƀ43�Ѧ�'EF�"����|�efR��H[Vu���ֵ�`��ɀ�RE�AX�>��Q�އ^�����oFp�)��8�.��O�r>Syz�+\��{�pUF���"3�mQ4(���%C�M�v��z���Ǟʓ*����>O�G�z]�L({���\Y�=�(�\���@�dϧ?����?��kb�3���mϘ��+�y)�wo̿����Ik�yp�=�v#=�\F�M�{��W����'����6�i�T�G�ƺ��d�{���K�q�1��/��>!lD�@g�>�����d@�s��O�W�8F7,3:���[��h����x*�1+�2Z��-��޽ٜ�������g��1c�s��x�0(}�Y����56��M����^��V9 �+d����o~����S(���|��h�d��W��v�m��o��a .i!2���a��e��_��Mc.�4�l��W63po(�V��%E��D9�N/]�^`��&& Vn��Šx̜���y����AԵRb�R�$�Ǣ� \��`2��� l�_o<3k���XF��
� ��Z���|b��%}�8���d��n���ʁ��=^���{/n���
��;xx1��W��8P�P�X���(���%T��mp�'W^J�o)�گ��Ҝ$��S�e�~Dq�{��:�8��ʕ�XX�S��Y��?�����v="�N��XJN���W}$��"�XEq�{[3���{�t����F�nTy�
�Q��x�Ʒ�s~�|N����4p���Er��Y/��$� ���gw6.��p�K�n���b�H���ǯq��}�@�y��|nO��X=�xf��C���X�9�=�}tLD��O=ēʵ�5��a|�%��9)gݩ�;�+BN�%��\!������A=�,4�;D��,� �c�rP��o��٣F����$h�u���;��3 `�#�}�0��^���yr�D���r���i|��|��7%'-�s���Rn�z����	��/��9�����Z�Y��gWJ0�<T���>1�o��?�Og���V��"���p��<ws�<8oz�O<�-�R�y�W��6 ��G�V�� �U���iu=��@�C�XZ�@���U�Fy'3t2�Fiѷ�}�(��Yll���e�`E{�L�r9��z� �˼�?�u��1���e�Ϙ�O;H \`�I�1�>�"@��<ї����AFă�Yāk���=a�r��ˀ*2�mOVy��8���?BQT<��=q�W�tT���ݘ����|s��p��V��V��_<��g�.n@��rtZT��s%����'�p��K��.b5���'9z�[ �7N����h�ч�C�Z�~w��H��=O���AhE���G<W�^z��]�0����;���ƛ�7lC)�YL%���:��r���_�j~�������ǫ��P�#�B��\�܊*0�	9�f+�����֤��w63�ڍєU?'����-YY<����[W���'��h���F� B� e��;(
��-���Z��!��x�!�/17��'>�=r�D���H&� �v+���Z� % i��K��@W���f�3y26�+��+D���C|���)!���;zA�i�	`�3!b���V9<�Ɗy��z (������E׊�>�)K/�$|��ou~��:?E�r(\P�S9:�z:U`u�Qg��)�>�W�� ��Mc/PK�=q�7�xu�YN��x��q�B����p2���~�|���9�rş��@���}�Yz��튺d()�˖���5�zp#S�V���
8dJ-NB�c!�gو�[�sx�[W��Ӓ�wVg� 8S������z��ъF�a������eW�_6�hc���@������ͯ����Ѿ[�>�;"c����VT�O�?F�(*v'��a��z^�CP��ң�y@�����%��c
�ϧw�&��-�|���80��NBLs�M�,��=���LIz���,����ݣ� 
���{Ϊ1�23㵞u��H���e��#`��F��=G�W;�cZ�fDW���??
4�)ʏ1��C��	��{;��0��N�49��%t O���)�*'�+"�5wX��K�rz� �q�_𩾗�G�{����>�W���@�D�į�t����]_ͣ,�uڑ����)�*��G�!c.��-�)eJ��;���w��9��C�{egn����S��;��IheA�)�p�s0/���ϛ�ݷϼ��;���(s]�s!�ߖv�I�fbD�[	����c�2�q�3 ���p����Jpù6gϝ�dw��:�����Ƹ',N#��Q���`#�f����dͩβ����U,�v5�K̋�� ��s�������iY�^�( ^S��SH]��H��y���u� bY�c��8�˻���ݦ���_o��>7� Y׮�H����}3M�T�E�]�xO���-C��W��\�>{c�����-"(#<�1�)RnS�s40���f���_��7��J�*m�J�y��	@���C��ů�~%s�k�\��s��A���7 �gϯt͙�;^X�s�*zG ��>c3���F|��c��ռ�L�zy�~���
,g���;E�!��S�
��Wd��`��6������ۼ�����j��Q�c�l����������+�>G0 ��H���n����U,&�4���B�2���>���1ݡ(cf����l  q�c:].��-�e��"�
o�<e��b�JT�"���/�q}�5�sܬ�u#Fpa�[�X����]��X��G�h��#�|H^�  us���p��C��� \w�#���#���ͥ�/�(z��l������ww�B��ĲL�R����$/��ó��ZZ�7�O#/W|R)�X^�ٟ�jG�OG��	�\/7�cl�{��r�:��eW4Lz��o�=յ��%�lCJ,��Q��00����6ƈk�B�V�)���@�{lm��|��C+pN��7��<�{Y�y��P:՟P6�`�����8.�C��ּi�%�-!�^��������wV���������������Rdg���B x��#��{)����I����]�1�����~S;�[�M9�?���z��+��l�zX`�ғ���SN���_�>[	)N�!�u�SW7���~��[�-�P����4׉t���H�Aמ������h���.8&�]֝�,����
�'W���d1��%.���z8Ũ0���IP>�x��F�'M�W=��*��X��峌�5
V����u����ďw�<O{]|i��X_�?u�+S��8��gƀw7���~��2�V}�gF��͇���(���(G������^���s�=c�m�����<rΏY�`������7;.�zs;�Y�$��,�R�{h�.8B0�>�����8{n�)a���w�,:z+zx�-�0���e���jH7��w=��{��{e��$��}AGe��὞q׫k�
}U��lt8������;V~ܷd&U��z����3�����/8*h���vϛ�z`�1�9�i�����M�\O7���ɨ��v{��e�R:����%�����/1;�"G'ˢ� ���0��|�"�j|I���x,/,iu(����4W6[����`���LY7�:Ե$uV����=����ݾ07��q��:�e;�]
�G��*�j/ߵ�V%0����Á$�O�k�5>,����nIs?�CL���X-.q}�2���0`�ۃ����/��I����{�{�C�Su����wQ�� �US�y"~�u���-T�w6^�5~�ٌ��doU�h,�R�~�<�Q�Gp�}�92*�z�����o�O��X\ �C� �sM��!���{�>�v�)��j�������o�*h�k��l?:}��;��<�aY��x�(��b�8>����"���e��ϑgɑ��Y:�@?�C�i����g?��Y�{(�d6�5V䯾�����.竘!&z����
��y������l�^<˾�Pi�Y�\�C�u�]+'�x���(���_B����Wz4�Б	��N�H��гw�ܒ�@��X6
�K�A��A`�c���;ٽNx��#}�i݂c��(z,~������\)��|b�E�P;g�߇�|�ڐ�kUG��`uVZ ��=i��R��AK�ʊ���'_�;�	���KxK�X�
�����>(e�	�g��7��;<�2�;גc�ޕ 6m�,�E>A�o�����q�9�����3Ǡ�F��Q>��b	���s�->jՁ{��G��ϋ!S?���ߺ��-ϭ˞� ���φ�P��]�:�2��S���=�E�,e��рa�a b�emv@���೧���xe��\C���w �5jIF ���Gc����/~>�6��qL"x�W��#�����3���]˨�����ͽ�"�6!��"������ W�EV�_ܳ �Ͼ��{�3xl��/�,`�� ��w�J\q���~侕<��O*C6D�?zi�}G�߈�Xͦ�O�嵭7
�5T���K-y���� -�{�ԑr� �y�3�`ݐ^��c�+B���]�"R��	U�>;���}x�7~���he`qy.M�e�c��d�-b�"��厹�WA�/�8{s=#>?�/EK�gth��z��s[�;�f
uD�W�gV>c�$up�'�a� >��VP��%.9h`<��%��g�!��~`�r^��B���51Zj��\KAf�D�E@�l���۴t��6G@�d���W`�F��'3@Gv�gπ�wvr�����{$|C�{��<a�q�3O�ǐ������C�7� ��Y�:��CF/-k+<MN��y��}�n��g�AUD�>�������$�5�!�/Ų"����/�g�lPh��H��G_1�����Dvk��o��v�a-F������ �S�'���/�=Ou���Q�!L�z�~��.q���Lp��R��l3�z)��~ؗ���{�EH������5� [�%��7S �I. �B%ƃݧ~v3V	L ���a��ɸ���5��X��!�L<��A��x�v����@,��و7���bR��D�$��K�K2j��|ߣC�8k����2a�����B���O\�G q�QL�V71PO���(�:q�����Cys/�#�AǪ�xT����k�^�4��YW��Z���[^�^Y���9�����̑%�?z�\��遍�9z�3eU�d��Y�ԗ�b�Ɲ�����^ڂA?�9#仃h���q�~�����v�t��nR&}V8�E�8�&�<��Բ0: ����=�:� ��y��+p4RFv��L��Pq$B@�ab�5�V�ϳ�s��_W�͒���G>�]{q⿇��NG��ܸ�6?^�@��5 ��sGG�#��z�^�%_=�DzV]�^�`V4u}�}H:�YA#������n�t�r�z�<���S�u7�|��Hau�\�m��@j#�'q3jf�Mx�<�{rE����J�ޅ�1�Ð,�y�/@C�����ys�m�ܸ����C��Z���*�YF��T@$
�Q�B�r���t��?�B�wŐ�����?�i1"�i�ܘ"��|s/�Fp^+�QQsaA�|�=���2|,�����h9��#sï� -·�3��͡�Zu��[ %�7�����9�ݟm<�,_M�;���ƙs~�<�0�}�w�T���9��^?�o6b�<�M4ظޟ�;�= ���<��K�0��O�A���o�}{j�6$s�2�t���Y���'-�R�@Ec��-���b��3���B&�/Ğ��9��D���y�25�G��ŉ����I>?|�]w]ܣ�d}wz�S=ޙ�`*�����U�q������^x�ê%��C�8P<,�-�HzF�N��e-��w�/W��������a�Y���@�:����ȟd�,��,;�\�_9!ă��,����ș�uFt��ߕ#`���KQ����g��A���.�2)���wZ���(#�P x!����W����� �� D��"��ߖWܾ) �
�7���r��	h�6|/�h��#���_Ep˽�;;��e@^�faՓ�x��v�K��F�Q�����ɀ�>RFfe@�������+��� w�>*��͝�~�M��zn�w{��Z� T�b "?�Wjsz��BA'e��@�7�R�x�̍q�x��،�䨓�B� �)&	�A/	�Ų�O~�Yw�ww�x�er�
�O�s����l^�<�{7���"d�d��&n��E~@�)x�C$)��<�G���T�Ó>97铇?����j�>��O����	t~w��zg�&>��!�exU2���j'��Y���d���>�j���g8������o�#�%O!!X1�O�V�� .�4yqi�<X���l
*��H��9i�b�xG�� %N���=��g|���P{T��;|f���}g���s���%"6�<�hӟژ�R @�����z�P�IE�ݛ(�B��*B�a�n=<�=E��֟��c�����q���P�#��N�W3݇�Y/W�'�=FW��H���v��\恩@[,�E��*����2�W�j��g��rV��}����ʉ@bp�:�[�%�B�����:���8s�(�ݩ���ЭV�}Î�^��s�:^��݋�`^x�(e��C��� ����K\���H����g���K;��;�����j�O�Q��;��eHV|W��n|�\���Y�[�-`�����>���>���7�y�T�*g��ũ�G����׿~0P[ѭ�޺�/���w'|`��;S=��Z����g��Dn��pȉO5�Q�_�A`�	3I�U��5X��{= �Hbi����dr��j3���1-�#Ј9�p�v�,^>��JX��XF@/��]��~xb�Ӿ$�B���,��08.�x+v��>�[o��5Bߩ}ܧ	��XXGx�9!M�# ���+�����R��g���(U�����#�8#en���uo�+Z�����^�8�c;ؘ� �Ї�!��dޫ�o=o���R=�CJ�n	)%"��~��#U(7$�P�ת�G��K��<�0����7f[�!�?{��Q�Fb)>n�!�b�4/���]:�I����H׆�y���N�3�C(�_e���oB�mp�Z��LƝ�w��u�X�N�\�uz��C�GsPeJ�Ho(�$(�ý�#��I��-_�[�������^�X�p�HA��yJ�!�ϟ�A)� n�U���j=`��`GΑ���L���#�u��=[���+�<2��w&y�:���t8Q��087��;�~b� �yL���r)G�ԡ���҈g�)�(��X�,�
�
��e%[�,��]w͞[Y�*Cʜ��d%��3����u�&;����F�Q�lkO�{x��4yC'�:3��Sy��W������s�(.���<ź\p�KK:06���Wk�M A��6�3�7Ox�� ���g��M~T�o
�%5�j�*���3�p����Q��s\����߲�a�n�bG) �%*�y�3o�^� �G>O_�t�PN��]����{��,���We�J�[�ɆF<�AA��]K�FO����*�t�;�<㵙����K@�0��?�����G@nV�����7F�'Ė�2������.{y)_�+���1�DKV�j�2�|��S9��Dx_�`��CU�:�	��e`�  l}c6퐾`�������F�Ư\�A-�u5�{�V{{�y���U�G����An8��� ��^�A�+�!���pXy�υg�ϕn��A��r�q�8��#�=��}���	��hj�c?�����ၩ]��~{����=/��©�!"}��q��u�@>]�~�'c��_n0���s�CK@E�)�NL5D�R`T��Ӏ��K��c�wMV�;V�Į�,�v���W O�[]��t��mR֏M�=��/}��ij���&K��S��==���}�c������6�2�gn�85D�(�MBq	\ cA�J��9��ovk1��QEk�gT�Q�uH������#�K�s��A���"�g��8w �~���|S!������)^��'�6z���CU�6�5�� ������9��8z��6y<c���wո�7�*c�9=�о�T�f��G��Q!{�V� ����hI_���m�� n�+��C��݁�6f}��N����=szgu����uv��� c"O����yE5�Y�<�φl�1�E���J '�6��"����踨d�����ފ�M#��q�+��r9*��G�Y5�h��~�:<�fp��	�>k��2���/~��!����[<����)�%\!,��G����*�xG��Pɉ���O�#���R����<;��:[�Т�"�F�j�� :'u�R~����UpV3��h0����:O�<��I~56s�{ｺ��t��S��g?<���TS{f&� �S�������>��A9m�q�v��e���v�At���<��g�>Ο?��`{�(��M!;���)߽W4��h	�@.^���Ë�1�xB�ځ�d,(ו'c�@�,V4�%���t<��"܂���]�gG�q*>F`��NetQ��+��p�kxb�h߇FAr&7c9~]ƛ�2����z�����fgUǌ��k�����?1
�8��r��K�Y�h�:9P%^6��Qw(x�C���.��~��V�H��|�с�|���G�q�Y{#o�u���2l2#"ޟ���|cp�X�	kH��A�	��W�8�����a�	�et��㤧��ƣx_��HS{�q��wS���F4�׹Ӎ9���=״�76<�� ,]JHF"|[`-�M��R�Y{��%�Cpx�,N`³���l��|u#����Sװ�����#�|l��!��7��q�;;'��$,���s��mx��'����[v�7gϝ����;�X�䪟 "j3i�Ą\��'[���.��ڻ����89\�W *3� }��Ċu`�g�>*O�)^(�(6�����LA��u/,\���:�u�� \��˲�椟���b�����g^��C�ґ�ߢ���g��A����KKe�ωm9���\VH�Eߔ�+��h R�U��v��嫩�b=b�O�����li�o(�m]O����|��pŁ�g�cx=O<�����,��z�uH�6���6y�ıb�B���ۣ%�6�#|���q�.�|��������o��2�Ň� ���y2述��f,�~��Vt�m�}w���W^y�ѩ�ߞ��?�ռ"�G���	�yJ��y��ͷ�K>tˇ����j��;m��8�Y֒O��Ϲ�t1K�j�:�T�p����*�eZ��U�����g{6��T9��s�.0�������L��0;_|��G'���o��}Aֶ@�@)a�/,F*]C��aG�:�W?i2��tҍ�a9�I�"z�Z������L=a5i���s��-�&[���w� /7(x׊\1c�R�(W�q�y�(;W�-��=>��*�+,���\ݏP�{�J���G����c���LЯ�i�/Q1G�1j���y��^��ݽMl� r�KAjw<�7P|#������p���D��p���[eZ�.1���dƥ������-�݉����5�f�3 B"��D��zU�q�/@��H�2 K/2�(�2.��V�������(:b�"/;o�p(d�MP�
��N%S�Ux�Xh��!�Y��G�������YJw�y�]����k5�;S�ݷ�r�(u!�_E֋�$���~���ߢ�d��
7����_�΃�=	$�I�b\}�s��%���j�k�_�g�WS�v��w��V��b~hz��f����?�����;��>�xy���T/�T�1{���	)"1��'v����J6�a�+?�,N��!�@E
���y��=��+B;ģ�����2�;���qy�7�ļ�ԑ���/+�fQ�򛗝��8��S�%O6��wb�}S��!F*�s�����8񯈘@���@7���u�c��5
��5e�0�_�6:_�{��V���uO���� �9O)7_���#���+T�e��C����Q�����l�P@Y1����cp�7��x�(����!hNmvӍ;YH �xiu�d����1��p$IW�W#�d����=�==���K�s*p�7��Y�|��'�e���l��H!�!�o�����>oʽ8���p�B#O���o<��O>8��L��O�/=����P72B�O�VXt��䲂Ol}�H��:ˏ�~,�-f��KS^HR k����,#MD]K,�cͪ2`iª���3:1�#ӳ����������=���/?4���S���xA���"nS A�N�
8�A��,�މuV��>��n}�F\����IZ�-�)�(�{`�Uv
��
���K��=�U,�����y�.�����c^���A!>Õl��Rg�m��˽����&��3�Ol*)}�[mxl��=I�hiQ���ͅ��9�����:��s���H]��h*��=�U��7��VL�����^t��7��x�`�ʵ�`�m���;s��]�lN?��@��[���=R�,};�ٌ�Ϊ�秖�b�}Y=S�wfDe}X�mf�z��������d�!��%��&���t����Z��^��K�j,�ݤ3.N�>���|�����6���M}����|A{��lp$�	�|Ę��1���%����2�˿�����C����n��j�&�H��l( @�%��ԩ2�������e%/'^ۯ~�����t�(��������������z�ٓ�>%�cFP�Hh�ci�HV���_�����:	O���8C�F�$U^,+�s����l6��d���2�K��<�;�>�m�=�b��"��g"?��s�B[嘤�˼.�=��P ��=�,!�P�~�
;me�G�v�8����
�W���#�ʊF t,7�n����� �@�H=��g���[bpp/;�%u�ɼpe׃��B72�[�������t٩�����܏�v��/>��̎9�v���,7��zX��l8Jo�]=A�{�]�. n�S���������|�dY����U�����{Z<�	���t��J�^���*7�u���-�&a��*�����{�IF��E?������=��%b�YD������]���ޒ)�y�N�����YGAN��LFU^-`@�BN������3�A�
��yygu���HK���9�O����o�M�z��i����7���������^{�����[�@�c����q�N���MJ���D����Sr�0U��z�Z���Z��l�]����w|��m�޶=k|�<g�n',��9a#��幞�H�`�j|Ye�dC`�)��G�� ���a���EĲ1˜�k��^i�#�0��uy���v�o���\	3W��r���`٦��˩^�x����>h�te�e��-ʌI�9�~��~o<����,�`p=���������=�L��f(�:B;�Nϛ�vb§�u��<Gn8�R-Ă2�z�o����x�<�x�!u��K��y+ K�;���"�9��t��oښ�+�ޯ�>�#r�����=~mE����=<�`6�}��1)�?=�1��'��pn'�2gJ�������������~��/��*�g����"|B��i�9�I��Ha9_� \�'���S���1lxo�eqϱ�G��H�!q�60#
�������7W7a��_����Ǧ����������*�я~�w�0��br�x≹���/l�"���:���)��k���8��%e�(.!/���n��� �C��3Wb;HN����7o�$ Y<��ωP, M@��r")�&?	�u'�EpJ�}|�z>��?�!h���.0�0�<�'q�������+��[���gU��9VP��G�xA4�	k`�>�
=�N3P���3r��?�{�g^��W[ϫ��a�����k����!A��j�"�By�� \K�G�˼r���Cm�x� �~�2yk��i_�G������_޾�A3�m=ԧ�w���`ۉ�3O	U�R� ���INyV�|�"/G�A��V<�j^�x�e���<��Y��~G�������ϧ����S���5�V���l��}�s����$#$���G����L's�d=�n�FL�ٿ�-�����s'T��uЇ�ķƒ��G�b��*��9�K�p8�9 �8�Y���|���<�Z&��W�:���?(p�4��G�~x`z{�@�3�<3��׾���b�0�|
��`��O�|�����J$=K}��y��ZE�s����uj����7vV:�;u��ㄲcC���g ^W���#�����usm��6��z�{?~%x��9ޚxn����fyH�B<c�I��Y!p`�%Ԇ�0�$E���`}���Q�+�Uy�2>s�x�R̽�*r �m
m��H-��d�e�ds�����7��?�b^&����z=ܰt0��Ct�xt�W-y�F����Ϡ��U���x|V�cE��F�p��Hs��ΚӞU����A�͍�|�ŵ�c���Kq��䰼����3�1.�1��Ws����[��#^���W��#������o��}�9��M7o~��Ov�@���
ſ`���=�m��xsp�d_Cn����8ł,b )UY:~ڒ ���b:��R��������N���Č������pz���_�{����>�eɠ�;яf奾f����ɏKxC<
�7�Ÿ�Q�'
�C ��C�	�ֽ�~="ƍ�CO8M��Q 8�����#%��a���hxu��%�� ���I��%��. ԃ8[=[ W�R]#��Xw	n�N<j ��&��Wvb~�'��xR�,;�����@��e���z|AO,ϟ�^�+k5�����Pv}�/-�z& �A#� �>>����A����1�K�x�>��eid �C�� �x��#.# �v���\4�n�ͩm=U ��^��G�N�W�T�C
"m��	����tBu_�߭9�Fg��)�MDH�H���	r�I&�����X��O�<u��^�q�?㑯�����G�ϟ����>8���O}u�����?���z8���RV�En���Y�QE���_B�L�`��:#>Q��$�2��*.lR��D�WQ�I��VC���/��vb�'���H�}l�N��;S�ܧ~���'Ҫv�?���f�55,y�h*��@�}ب�7�7K�*�1�`����<�k�=L <��'� 0|9� ���ʊ�cJQ���{zPjz��;ʾ��E3��Q�����Ж��^��W7/���N�>�?�gk)O��r���� \A W���9)�7M�<Ժf���V;�����^FP�e���������"� 6�{��yG�(�����с�{�|���<������E/�x�F��;�n�j쑟�Xv� '��y���&�|�f�����W�ZU�x��ݰ����|��UW�Sgq��|3Jћ�*��x��͏ʫ�����/�X��L����������:��	�=�T`�?rRz֧�~����.��T�&�B(�o�w��jHw�Ky�߸�U��ܵ�,Mī�N:��� g��S��٘���V��jC��D�Rʳ^xa��@�O^\��vi��V���.��sd��ޓ�M���o@J��h-���V޷QZãK��D�8hϽ��� ��Ch�B�x?�Ɗ �"����A�����7ٗp	�g�Teh~�[�"K����$�+��������2�D�����8� �& v��0��2o��+C�|Գ�h����J���G��̑z���VY��.�7�Zz����W���2�PI����9��,.�^��������"\�P/V�TW����e��ef#�ʈ�P��F߹ѽ�J�>����Y9�ֽ�"���hNj��ݓ�Z)%�8��yvf\E�)��*�+74������	+Ǭ����k�
iP�[eq����hpI�&������O�wA�Nn[���M�{�+Vj�t,}Dߋ�\Ь�/����RN���l
`s
���ʴ+�����R���ҳ�D��sک71�tXBE
X��~ `���� ' Y߄!">*"嚎D��g\��j�x�Fxf	e<���i�V�y\4� ��E��D	���UB<6�F��d�hg�g`�#<9`�k䱑� ��1�s�WE�2 �x@�p���%�����R��9 Ͽ�d腗V����~W�9�P���K_&U���ʌ�
�V��<��ʻ��8qM�k���z	-��f4Z�΁��j��8����6{�l�{�3 �H���Q����I��=�f8�t��W0Y���P&�a'e��zy������eu�cLMHH�Z��
�/sV�J���љQ2-yZP>W���]B��e��[B'�78�<'?Y;���͒o�O���=������4�����������	�����;�J	!�����"n�h�G���C��r���'i2�Yߥ���MרMN�/`��d�o�!��b{�|��G����wbMJ�OB<O*B��)������8���>�j�[�ܵ��'t[e/�x�9"�^x#���TD�2�x;��X9�X���Cſ�I�z͞�K�nS��r�٠v�f�)$`�=fz���s"^�9���m��t?˷��������%�]�ǘ[�`=�����xӖ�֊�����^��ť��<�Y[|Z���ڒy�{�L*��:�s���վ����y��,^>��1��,n��E������1!�.�9�.P�sH�t��������;�����H[]G�L~�P2NIS?q(G�j�r�v�5�W�nԢF���>;/��5_�ZB=�]鬸��n�Xq���3F�مS=p�������M��>���o�W�L|��π\�b�3�%8�F��5܊"Cy�tGL0<�ǫ	�^]b�pE��Q%(p��[.N�!��#��Y�q�׿{��W�5�߷�� ��W���u5�Ɓ\�j�����C����|f �h�M,��.�ʫ�%��'K^��;�}��=L�x��������^�KWsm2�5e��%��#^RG�O�W������ /���|c>��|D���Pxn9�]� �H�R�Kt7g����5��0pqP�"�>ʯxe���9ʮ����ֳ���\ē�8z��ު_�����i�2@��@bN[��lؐ�i�Dl�����O��8r����K���������,q��t�d3+1�L ^�Ԟ�m2\o�tÎw9�7r��o����U��M��Г��x�9�[�a>2��#+�o��|�rj������&���%tR}�$��{��G�b]/�{뭷�0���?�M�s��_|p�G?��C�h萙GƚƆ9G�\w�0.=��ܖ��5�ɱsԽXR���$4�h$uX��0!'���뮻t��: a�'R_|w������������yJ<����6y�Yg��+�˸r�T�s���zmG�o����?1jx4�8��s'OƼ��1�8�\�.�i�j<��8B�h0*��Q��<��z{�a�*����#RY���}��3?H��Ѽ�	z��� �P�ʠ����R!V>ȫ��m<�,�r򙞡y�\��f�����2������
�e�Q�������P�$������͋hd��nզ�<ݝ�S�n8f���Ȇ[RU�OSs� �+^W��d���Q��ŉ���4�"5G����(�Ps��_ڼ���g9Kf��dj�a|������v]L;!���v�Xw��j6.9�>�(�P�B�'��=�qS�ڽAQ�g�Y�>&������!��ب��Ʋ	��{� �$?��sJwz�CH0L�y�$sA���ÞE��Aq�c���>�ܺ���� oq�X�,s��lLt�-a��?�����8��0�o��"��'���W��9��P�tW�GlU��Ƭ�˼��F��"��8"��h��I�y�XF��y.\�������on^{��Y�Z�HK����xÊE���أͅ�C��j���G1gߝ�����==�N�S���[�fV]|g8ωF�N�҆ b����?^d<�l&`�ʣ��7v^���գx}ţ=�=�Y���u1�UT� Bxӗ����\;8�! ��Q� ɾsOZ�(���:�<~���J�\�.,q�;���t`�V�Ο??o����	����ܙ�'>:tg1=���ߝt�7�p�;�\~��|�6Kk�B�z�?�1�]>�y�=�>���cl)s���T�.F��F����g�̠��g�+�ۛ{�!��wy����T�㱰"O��q�d�xg��j�DMs�ѩ��f�S�ɨdu��>��eع��/ݸ�]̂s��l=�R��V�hY���(�h�{L ;;�4��tӍ7m��1�4A�����vh�O}z�o�������������@��Cl�ƃ�O��ܥ^PQ˪��t�2P��^U;�#%t�uo+�Y���@ O����|�x_����?:������qy`R�� �ᔒD0 ���p��G+&���_�����/^�������'P{��'�����>�?\)oA�����X1�I��@���s���� [�T�2���W�3��JNƺ�:V����|������h�����y^�-M{z��U�Y֏�L�+�v�S��;�!N1�2���L� �)����&!y��+_����(�^`���_��h��_Щ�:�G�]�K�
�����0)�{�S�Ԋ���U?�G��eՔ1�&cC��(�=b~T���3&s�če>��B� �"V3���ҩ���6QZ�����Нw�y��_~p�Ͽ��!��ȏ�����A��﫤��QzTo�����?�^KB�L��.j݋5���7�����{�SA&���@A�o�i�w,1����������{�1hr%�
ٽ%#������H.��7�ھ������u��I)�k%,�{��cYu��F޸�n�P��Mb��.p���\
U��,�Ώi)�����u����k}�*)�nl�l� _1ƀ���m(C2��g�~v�1�k�#"���[{���2לc����ĚC >��R�r3����c�=v���n�/��E��\�]ЍW"t���
g���0_����駟����=�'ڂ?Xt	W�ZXs]��f���$����p�t�f%�!��mKo��.��ZSw,��=�U��	"<;κ�mg/q�˼W�PV�J� ����̌���p�/���jRV�m���<բ>�*ب�̱��P�U0�Bgb�qz��+�Ϫ�3�p��$��� �l<~_[_�o��Y�����/��x㍧����M@.�������R��9+��vؙ�*oZ>���\@�����e�,�i�Tk�ֹe?�Y\��?���NY�r��s�^h�2��ʃO\�e8��?
��G!i�yA��ZIǏ�:V�*P���+V��q+�8��j���r��� ��Ve\��5q	�xת(3n��o/�.4����a〺D|���_��>\������&� �r��Ʉ����z���ֱ��7��+���̾������b[����μ`�en������9��m��ַ�5���[EֶRD
�P@������>,������3m��n���я~4���R��Y����P��象��(���f��鏽ul2eE���z!�?�T&�	�&P��Ӿ2�K0������3{l�:~	�0�X�YNƍ�oxm��~�77~��o��#�l�}�~��ζ�@�\YP�Ȟ�s�<�cH�U`����T2����rKr+��cw�y�Cd��}�s��������^n
�/���ۘ���Xr�(�f�3�����E��b�%!��ܔ�0�
�����ܥ���<(�A��ٺ<U��j��*�~���oW]}հ��L��%[���������q��dj}|Xh,s��4�(w��bGL�ukn2�{��MJ!ճF(��Ve����p� ���wX�8F�K�	��V{`�_A� ��o� n ��>�j��
��n��iD�S���=a�n�)�/+p��gM�=	`t��EL!�q�I--^;-hj�
V�"��E�������,��ꫯn���K'��h��:e����6��}�˪c����|��a�����zX ��Ղ&�U����E�B��v�=+̴�OYq+O���ŵ͈�r�MԚ����b��l$d?�wZ��
����V����
��c�m�5X�g�ڝ��}��W6~���w����(��!������X��ס��J�c���C/�`z����U-zz�We������%�����k_��?o| D}���@�g����Ӎ/7��O?��� ��%/&��]� �&��Yy� o�����f�P�_�g�X|��|�Th��S�ΐ�\�s��� �2��&�/6�Y�׏9�N�#�r�p]�5$�VTҕ���1�F�{bp{ �w��ZN/���d	+3�k��s]�>�"��v�o7tX���o<�/��/g ����K,t .�WKd��1�������9��U�N]cLٚCc�
��}��H�E$]��t��\P����Ohc�����m���܎�Od��Y��\سΧ�&��>�s���讻�6is�t{m>��#�"l��,A�jJp� �6S�ӝ�x7lC������؂Z����w�q�k��D_�c� �>��).�iU�<_`��!�ʹ�%R~2A"3���IZ/�}�:(D�Zo�1���օEi��Z?Y����j��iuf|y=��3C�ᘥdώƐj,��v2�pq��!�T��g�Le��g��~���>��<���W^9�������M^���=�u�����xfdC�gU�k���8�c��7i��2������,r��̬�����9?e�I�O���_T��)6���9nV����zj4�Tm���ږ��Ye����4��n��Y 7-k=K]���=��D�t��8�\X ,�L�B�g���� �Τ6�����^��LZ7J��V\��I�b���ﱬt�"���m����ǔ��vx�����5���]y. �I�bZ<rn��y�5a����Ŗ����t�M�s�.����l��6�[�	��ȝ�����Sf^�X`H��e�߸N&�M��<��ӧڱ��u�p@��I)��WK���)����B�Z�h�#��ay(@�׾���z�WÄ�Z(<=RPZ�{��I`i)U �5F��B�����+�j5�t��C���?����g��b����(P. ��|~�����SOߡ ���
X{
U����R�������X��U~����c�#�������wn���y�uב��}��Ƈ��ho<����&�nϹIr'c�sflt�~7��ﬠ��2�h�#��9��n,qg�gn�,���vs�</���~�^�����a��v�P�|Q}���{��v�휃��5	~��[�/��E>#wXאKV<�R�U��zwz|����7,�5!�BO���i-�~Ԋ�@���>0��AMH�i��ݭ���o��ks��b|$c�v�dk�u,�)�6fQ�L7������S��Y5Ӆe&��\hM�Ȫ�`��CPw��e��v���/��/����_��W�K���>����;�V��,/Z��o�1�#�rޑ��,7�L���wtr�*���2a�z��N��nϸ��C�h�/�f���B�
#�۲��Z������wʧ����ײ�~ik&�x^�Ƥ��է���̱nG��_+jV�p��a{*ḛm����&�ɱ�s%Ô���� <F]�,�Wn�����r�<��;�o	_�y�h�U$�Bڇn��c�bȸ�z��������i����l�p�����8(�*�n�"XUa�rDv\84(��;V��;�c��)R��0���Tef
���U��Ў���*y��B7�PЂ+ߣX!��Ȕv��&SJ��ڼ=L�ӧ��{@U�WcC}%���Si)�iWYu��aCӲ$@PXj��Q��&���k��fM1����k�	�8�������W�Q�1��{TΥ�X
�\;�ӕ��6y:���l��Pe��`�;rt��;g@pc���H�M����ژۈ�P--|�=}9�0�|!�r�39�>�ۯ(R���-��r���a� ��P9p���h_��:���Iu9V��Jw$���+_��	����/����>S�1O$8�2N����Z$X�<�\T�V){^G>̿뫶߶�K��Vy*i��%�X�Y�YZ �_Ǝ��8'-d��I$\�z��׿��ۜ:��½�naEǒ97���	u��J^���ʝՠ
*���~��\��G�c�<��L�E.��ИޯH����Ӈ�rm��>KK:^�E�����R�эVY�2qi�
0 ;��YP����	C��Z��De��m1����B)�5�Eת�Wצq��@��5`�7_�6E�6�p�:	@�+���c���q��<��U�Pܧ,V��"ѥ)��b2�C���?|�,k��7W׵ $��<���]�����=��#��j�p�]w��o�l�+��EI�O��*�M1�~�}����3�U�x*G�5�����җ�4��i�U%�1E��eC��f|X����R�}k�2I����x�r��y=�,�"Q�h� �����k�h%yBx�}Ry&�5�<�����J�Z��n�
KV����ư�1��7�g(���s���g�I�r9�l ��X�K���*����ߴ
��c�y��b�,6Ȯa��w�Y�'�I��Án����#Yx�����mosڵ.=FU���<���Nfiί�+3��:�%C�̃E��h]JF�4�"��̭��z`�_���������� �P�0P�G_�t���8i�ժTK��9˯�E=�R��P�	��ŗ���T�B��u�Y@���bD�[��������1��'��l���!("�'���R%������,7S�������?>ծ}/1�mAa��XHkȒ2��4��c�^�L��Y_j����Y�i���ti��_i�SvU�e�Rf?ڎT�zʬZݧ�f��!�����w�ڷy�tu��Y�9��]d</�A�kBmS���	z�u6�.΁eH��<ט!�c1����Z�ac��g?���۳�]���%2��>D�d(R���S�s:�޽�=7��I�>yy��q�+�+��v�yL*�~��p�b½PYyd;�J����=��=0���ַw��Q���;x]��7��0�F�|J�=��M\O�qW9	2q�E4�I�	��h����.��ڱ���Z��Mg7$�� .xZ��L�LRf�Vc��\<?(��� S��2V+����Qf�א�q�b�
3�ɊƢx�-�������_�@��wN�Z������g�s�{��Ų>[��Ԟ��
�Wl�@; �&��ϐ��`E7������k�'�.��$�(2�"`��Tc	4m� ���^�%8��
cl��w�5���=�x�}�
A��˱��O�kȘ��짂�c��2��L��ߝ'm,�@e[���C��f��:����j�0S��Z�O�z뭧�뮡r	2�9n�9���=�s;�T.!ׅ�(���R�=�+P�� n^w/ԫ����Y�U!�g�0�֫;6����'��,�h��g?;�d��if�ʰ����|�Uf��0e�Y���TO��Ib&�� �t��։���"ƈ�A��]�1�Z��rB��I�d.l龮�xhl�����f���Za朗��Ji��%V�B��P˗�u-�J��կ�* ͜�ט_�%A�7cYT@�8f��}]�Fu㱿�򗿼�&n�mH�]�r�\��b��m�mڣ��J�<�1&�����ӊ��Z�&�$Y)K:y�5W��) �;�cfU,�̥�,��<k�CX���7��Ȳ��$�:'�s�:�)+�LP��g�%���PD�'m�������y�S7�|�mnm=��K��B4(\��ّ휇�M̾7�1��1�X�7nJ^^j�u!�c���w�yPγw�yw��.����%�]T~9���#��Cn�� W9hNʜ���]%yt27��*�� J���:�'X��*��*����=P�|G�;e�y��w�5W/ǆ�ТWn.$
�1�L����c�uzB�2�ص���\D���i��		nI�qA��|�}t�lT�W�(�L+����B'P����?|�=۽7�x����o���]��	n������EimYgaM٣�1�@Q�f2�@���x�W�[�`fy���w����
B�ٴFJ�nJ�;(��&o�(C,!@J+x�d���>��bL�rB �L�s���j����̜�ϐ<�nx�X�u������ؿ��/�3�°�h��B�n��\8�]W�X+�쿌!O9���7�9n�a��K�Ks��Hol� ��QhHl=��
�)�*�������b?2_��2�qn���
=��(Y�@
�>j�j���&�?f�"�v�u�큰~����?�4Q�?��E������Yg��=И�*)�Ϙ��}_-=c�J��"�`����Ts��Ħ{TkX&�,-�[��[o%>�ډ�w���^�e{��R��p�}��L�SpdZ.�N���7���}��w���o���O���Βf	Fj�f�Yaت;]ﺬz��|��,�Q�N˨�:��Ϻĺ�9ϗ�˞߱v�\sg��_D�ܞKy7�l���V�z���h���_�\ .n��\{�e"G����|'��w��8^#E�*�޷��ST{ʲ�m�l�p�!�g��Z{R9 ���0\���O}��믿����/m�l��� ^o����:�wUNr����,*X�嫰�6G�w��8��q��Թ�ߍ]C���y*�󹃠�Vff�R�#���'0��vx@�#��~�����e"˵�nT��W���p%��1׎� �v�������=-J)�l��u$h}"������p��*	i��=K'i����zBo̚������:�UV�9�_�%���ͅ��] t7C�A�Gz?cg�����qݟ\w�-��2�;�u�]�c!HM��q����,�� %PCyct��7���5,r?c�~�M�a���FXp7.� ��8L��+{h@ �7�#CR��_���=�ؐ('8�&(�w�OO��#G�YWno[>��˛��2W)�Ӳ�%U��/�Z_u8�O�㴍��M1�y���Xy ��&���K{�>s&$iU�-�39��	�[�&��^稵J��-p�K\�]��.7���/�j
ؽ�t�$�W��qx������.�,c�7.�!�ғ��ݹV�*{��h��jLI�X��T�O�eE�{�	J�eռvM@>��QS�����a������.����QK�|�����)@S��iŵ��2�T5��{�F_ݻ9'���uQ� ָ�\i��Qw�*C��s�1�
WP�¸.����J���W'N�-�|��FP�Ţ]�O�ӳ��^?]��y��j�˄-ۓ���`����fc�����w7���� � q?�����^-$zT�k<?�ϕ�S]�c����z��7�5��P�	��gAm�.Hc�j�N�RsN+p����qZ��,�Vu&E���ZrQ��|P ~��\����j�������R٫�Ķ��#)c���i��g�p�1f������o������d2�Vv^��W��d����[�!8)[���m�?Ri��B�WJ����'?��rb(� �*��L����\�R8�����!G���aM�~�A'�L^�k�,�ۣꚪ�Q	��A.�)��y��8������ws�7��U�M*'�_����	1���?�	{�,�iZ�ƀn�*��N>T�2Yǘ�T ���a��U,p�6�{���5�����V+�<��J˕�rim�8�����~��<���g>���ma��l�6�uӂ�<پ�[Z���I �D��w��=g�7����B7c���=��HBU�lw��	�*�J�Z��m������)�y��$0�=Za�
�WgWY��t�.*w`͵2��z��PE�g�YZ�E��$�yJfd��c�����qZu�����B$�6��D��--��-Y�х_d����K��\�$��3��]�[~�����ʭ���[�6�����@߹=���ž]����H�\���|��&���c��&��������P�~�PЪ+�&���Č��0(��M���-ݝY^��1������O�3���d�j��b�^+�������ʯ�ӯ������Wc���+'$ٶ��i��	\��K�D��ֽ�-��Wj�����t <�R-'�d�iyNw��VV��C��r-���X�+�k\j�*����Zw��|'�����l�-)�f
u���*�ӂ)�sB�ǹ�Kf�z���~ T�>t��{�a�GK8<��K//�Ę�
e�4�jAS^���Q�9]3��>k�M �w���������-Co��o�eT��;g�ݕ��\>�d]��z W�\��ǭce�C�0Q�2&����E�,�R�d^��9��@B�����)#3f�Gɟ��N�z��a���	�`���S���%%�LR1N����u��	��n�������W)-�s�g��%��R�6��N0��!��꫆�x\��%n`*�\w�uk��.�
���Qȶ�ϙXA;�1�"g��~P�'��f�M��/h�\��T������_�^�ƪ��9#���gv�:~��`q�26��c���[����X�/� T���Ǘ�cX]r���b� 9�Z��]�Jn��g���� ��'\�u�R�Q	��bƔ��!��Z>l��-�h�z{�\�n8F�JC˻K���a�O7n*=U�����M�K�v��~~���1�"���ޫ��e�!7%��^���S�Z�X�rC׵䷪�&V�ᓊUvm�͘�޻�Km��׽R�_��h���#c����>gᕵp{ҹ4W�@	 z �wm�]u��6��z�ߧЯ�;������KЯ��?���J��ҞE�u3��@�%+ݍ)]�/��h�7�x����p��-@&����H	�fUhJ��� � IJ+-�h rQ�ag�Z�m��\?�)��ej��ؽ���z�tKO-�U�3.�d �n�馁O�Uq�y#�q3�E���ɰbG�}�t����e�WH~�Xg���g�y�@�Q$M�;��+����{�dN��8i����ʹcb�^����(��E��M�;��L��n�m� UůW�)z�)�(�z1��?��m�$r��-c���\2o���|9Y7�{4�!�YMA!��D3u�Z������Z� �]�܉N��G������޹c¨~��3���Im�v����[�c �n�cG��e�h�>��O�
D�1:?d��e(��$���̬��{�gȘj��	����qc����(Nn������Y�A���#�-���_�:��aK^�>��O.�Ct�gX$0�m=�s��*�����κW�Ҙ���?�[^X��K,�ʆ
$��uΨ���iA6~X������#Q��;A��ڒ`Y�R�\&$^�D�����'�sH6�Ǉ-f�k��A�u�RXP�+�R��Ki��Y��)��9�F2�U�b$�R�jY����q���w�2I����ߓ��{���ڪw귴"$@P���j�L��=��M����XrJᆰ���&U9�c�U��ɯr_��������yP
l��Y(?W��I��&㘍�"BrY��j�m�I���/�^z饓\��OΕT
3&תR*,j��݋+�"i��D�0i9u!��H�=�T�1A���&�Nɵ��k�/��/��XnY�V�_�x���H.�(��jX� i�\�?��g�������⮲���_���T�`��s��k�
L�O�a0^�V�k��p�UIy*�֬�{eX�k�\����a����%6kq�q�ӫ��F���y��p��y|˙�V�Լ�@�_�7m��T�3-=�`��;���[�?��I�8w u�����߫
��R����9�X3w�P�E��%`��hlc�ﴇ�7��Ǚ�_wC���k��� 3��tm�ի�CU�U����'m�,�kN���C�^��zS~Z5�:�o��y
oy=�`s���(��3Ǐ_;���w���X��N����8���.�W0���������7����A{I4K���'a ��v�R�|��%�� �Z��_��Wp��y3ZG�0���KZ'�W�<ZSJԔ�2���ru����X{]�y66nh��`��
<+(J0��y}=q�P-d�r7�U�@eD��gK�������9�+�V�q�J$2�9悯�'�����*�ʍ�]�� �޵4p(�RvO���Pܶ��.�����U6���d�}�<������L'��l�Dˣ��{"(���M�C��AU��ɂ;�)��%_9!�E�/�AR.H���~�������z�$V ��UV�1�N�����gѝ��X�e*���i��V%�ܴ�FQ��J�sN`��%��4drI���|��>��r��-��~4	��n�B��ܴ���q,@�[�[�2�:㳴db�;h�����*i�qKNy)z|?����[AE�VZ?��
�>�� ��v�@Ջ�I8�ʂ�D��g���{�o�vl�L�����r:R�u�� �P0^K9��ŭ�!Ƿ�_������}Oh̨���2E�����IK4��l&����q0Ѵ��6s@��Ʒ��٬���\&��W/��hU�ӶS&���Ԇ�y���1ԾY�>��q��\Q^��u* �-�"c��n f]�WQ
�\�j`�Թy�:	��N��n�! H��X׌���Q]��6.�k2kĦu.�3��i�^��K��}%(�� �qZ�{	Sc���V̱O��c���=��/,�Y/�����X�ǔ��y���o=KW^?�>D p�|�ɥ�bO
���X�AZ��\X��@B���D��'Am�����1L'=N��O��G��)YnJr��+���
p�I�U��*[�U�yMyIzc=e1��P��Q�FAH߻�%/e�UG ����;я��Y�઴*ۡT���b�y� 7�"`.�) k"�&ln�^�`��t���%�$�P8	;)���C��
���.Z�PoQ�i�Sm[X{�8�\D��Z���:|d��o�}�=�y�u���&xO��JfL+��HAyow�Ҳ+�|�7h���6�I��Y��Mr�Pc�=n�,��P�;
0��^C�W9��e���wʆ?��O�w���ʤ�l����{ѻ^�;o�>uN�߳�KZd��	!%�S�R�����_��p\��r-�U�!� _�Y��Tpb[���II��d�~��[�B�X_;h�;���G��z ��K��uM��\7���x�p4K1��>z�P$ �A����GC[� �Y;5:d��cf��􎪠��q��(���n(߬���	b����5��{@��&��3�O&�&~�Ls�!��ұ�حj1�Yn���{����
����4f=�T�rᰟ�]ql�C�.�H�[��3.h����eϘ[�D�h���%ȵ���7pw��ɓ{ڦ��_c�������H�;����v�Ҕ��X�x��{�:�$嵽�@(�������?�x��G����:VYP�z����c���c���S9/�eR.���Хte� �i镲�ZU�U>�|k�l��uJ�ڋ��ێqU >��nY�w�k<��k�C_��޾���SiJ���ʚ<elIe(� ��VZ��a�
!�-<ޔ��M!��nj��Ejr��;^���hU7�?�WN�'I��8���P58��1�S oY+��k}ԅ��Im��z��N���K���`����Z��ع�歋G�Uo�r{Ai�������st�y���Mke	]���E��8$�:<ld ���!�b��p}�覝*/޿��J
v������~�$[����R-P�f��7���7k4ç 1�����c���Z9��x���{�L�A�
�sq���s������)�ИR2�
���@d,g��<��P��s����u��=w�P&O֍#�%�@U�-�I�q��L��U��S�T�M��=#�~7��c�&u}�_�Ai��V@�?+	�����۷�a�8 �� <����/O"�M2S�'O���J9Sy8�/�ޮ�����j+�A���GE}P���:��a4�3 ^0En��;�H�N�,��1Bӳ�(��ާ�+�n]��leɯ?�������v�r�0�F&=IUX� Ҵ'��{{}'���~�hg�(���53�k��DAĊ�����4�W��kh�����\�a��l��Ni/A�����������#SA�����Jε
P�B���[&��(�5f0�7s:쫬
�Gp]e�r����aTRZl!�ajΓ�F�� ��e���l�})��U�p�\N�[ۗ �g��L8���[Ȕyu�=Fi
�V&�fu�ydb�x&��\�� p�	�]h��7�����R1jG��ٟ�v)�n㸟�-��;j�pΒ;Nr����-MY ��] � �Kk�1kTo�����>�I)�{I'��q�o�����ǡZL]l���ks\,�k�k��y��7)�e�bw�3�5���WAI-����&0�\�~�}�ʂ[��1���Y�6A��I_��$�<�'�e��w&ָ�y��;B�:�q7<9��'����T��^J�n{LZ��kU0P�j��X�3ηTa͘�{;�����s�]5�ܶ}��̔Ou��sW��
c&�& ���1�Tp�'�RQ���Wt�W�VԀ��d�|���|祻H6�;��_��;������k�믿~OQ�rT���GL���0s����^{m���N����߇�cA��N������X'!L�`���^���E�vO���-&X���f[�����`Xq̀x���1�kO���-��I)Īp���+�Ǝ����
�����s�Ϟ@����%8���O��7�����_?[6����?���b�v�$uQ��ݞ7��~�Ri��~����3��m&��d�����Iw�c�'7������Ë��
�	�HVk�m��j�c�UߏYM����x����R�JU1��"O�ۛw�,�Efz��B�֕i23<��e���ۛ���SD.Gr~�� d�8|h�w��L��Jk�X�b��TȘ�Ԥ�K��udl����#K�����rݟ��YU
4`p��T�����v�A��.��;����<��M�VA� N�NUd��h�mQݪf�1ݳ��^��I�[���8I���>��D��q����7��`&�'�D�-�X��*PXAC��\ �;&�g]�W���B\�� �k��=�,�#�/Z�hz��ͯ���x�v����j�,R(��`��UÚ^�����J�0��Lp��Y�ǁv�A�ra	ҳ<U��J�����[ú��u�J=#A���RY�z��{��]�g��c��e�m�	�,�7 ؍���Kk�������˙2�GZΏ�|���7.,]�zVS!�y1�����ϩ�@c9����X͛����2��]>7v�b�wd��ɠ���5��?���3�<��{�G���kVK��ZZ���Rms�D��<� ��(�,sIZ�h�%��A�<��E}+�e�l�'_~����x��њ��+�l=��'�G�1�h
/�n�$ܨQ՚sc<�o���;��1��ǎ�s��=p��~�ӺB�;s	/��8vxg�`j�rh��z���ZS�D�Aȵ��U>S��Z^K�aC�5�~E��a�[��ʜ�����YP�S�֪㨖߳0����=hN��ԛ�	�*���ws�3f1�s܎ݚ@�
�cm�n格����c�3�����Ƹ �r���p^QtRiN+z��u.~���g�XOA=rG�'���İK�TZ)�G��GO����ֈ{Z?op5��r��$��*�c�K��ڑdV5�1��7�m�\�u%�]��4�B0�B�ū1�=����i�'qk��0�1������%j� ���2a��I������
�u��=�-Ts�G�}���=z�.V��a=��[^�s�K�y �Cpff�\�	R��{BA�op�t��'��=�v��9-��W� F~L�Sc��T�EW�%��}N�c>Fc�6G���N���U�o/�l�*�<ᱫ�֜��u������p�����D���;չ������ֶ�#�"�MA��+��w�����s��{���*��,�ѓ�P�M��^hK�~��|�2[�2tc|t�u���p�e2C �n8�ꫯ~����ZI/�����O?}��l74�5��L����U����V-m]���#�����?l���kC|Kj�&���qQ����/�|��w=j}���b��O|rj��5�+ӂ�9��{Ǜ�X�5M����UV��yc��zn�%_z��;ySahܭ�;��#G��|�4y,~e�Km�>��[oc�[�}��o�]�i���U���Q�=����{[O=��IC]p=і�
��.c�!����gJa��ԥ쪉�^WZg��<9�GWy!ƀn����9��GS���ﵽ����)���1� �5����oV�1�@�N&RM���Hl2`�2�]��dB���zP�5�u���+ː�cG�2OE3����To��Y�/%Uũ*sI�"p�C�L�A���Zs��Kȹv�V�Ƹ��������oY#X��»���0<�i��ۂ��_Eko����\p4c=����@ v�f�y��w��R�� �{z��g���}w�UW.]�Z�r�A7�p|X(�Z�c�BY�ȜK
�j��ݫw��ȅ2��ˬ��<�^�Z8�\L,��s1�ס����[?��N���K����UaYZR.�t���T'��]���'5�:���w����1*tm?��Ng���	`T�2�"���s��[�8�YסU���Et/s�w�U�36Ǧ�����,����f�'�O%Q~�\�d�b� �6Ɓ�G�AC�[_)��.��VO������ۅ����(s2�G��*e0�R�U�"����\7(a�4�RY��3���x߱k_�q'~��_�����2AO?���K/���r��g�-�}���%�0|&���.��U�U����O���4��`4����f:C�q�7@.�Vy����!&��������:skP��{3l1l
`�2as2�eV�LnM�B�Ed�\�W��<7kϒ:�`����zN���	p��\X�U�Q�T��quQf����7� �>��2���2'{Np�c⍖���uq��.�{P���C�	����.�8\l+�M������඗��qc<Yi/ u/�ױ�M[�p���
���,ŗ����Q�z)�Ɩ���(��a�6��;ZG�0=#���9��k賅R@����+��(K�U�y6�� ������!��d��S��[oo{��d,`�{�M7m5<s`�]AXo[o�H�C}x���ʘ����Z��fy�?�x�(�ѷ��.��u){�g�H���dq��7���k��2�m�;�$&�믿~��JWB����O�o
'M��T	�1ʅ�r��s�1��GW�b�~��Yee��ڔ۱2��%AA�|W� �D��^+�Ra��j����lt��G����a/��8�X�5+6d)�\���2�Z ��5���n��c��֋/�8d��渋/Iy
���0������{>���^���
hr�`Uko��=7�_{��. �hK����ӻF������<� ՘�	|�GZ����uF0דWÜ=|h��o��������	�f��z\?��5L*=>α���1�;y���R��2��5d��s�w��דI�"����I��	�7bqٍ���'�������/K޺�����Ϟh�!v��g�"��*MӬ��wz��+Q��U^���f������p!�QO���p�Š��giH&�zLJ���(�M6��Ў�� ij�@3ZI$�5&@ .��V˞qѐ@�f5'�J
T�*p��<�~ף��Te_.z��]�u�	�U���u�9������N�D,�3y�VP��R���A����s8ۣ&���~UQ���/�hJ�H�Ė(�Pi����*S�1�@�Z��x��4���[�v�fq��J�Y�׹�X�y�+���i��o���ulX-�Lo/dz%���l��7�,ʀ��S�]O��}�Lg~���$���YH��qn��Œ����`!�j�'�� �V�۫���^�Z�j;S�h����/곢<��rR/Z�JĚ���ϣ<Q���;B��[��<�b�jp�^�4���6���O���Z�cL�����f�i]2~��(���g|���1��^���)� ��.��D��]�`�-]�F^|Oi0�[�JҘ���@J=%h���S��9 !�k�n־�EA��ɑ�A}�>3�G����'~�����o|c��O���^V癊Ln���K�p]��a�������"a��W�Y���f���~YQ���*��Y��� 7�e�>�̡�����h� ej��yV�wN��Y��:ni=�z>��I�AV1�	[�e[����a�'�ZϹ�g�}�#_��ƲR���\�iO8e[��
X,o=C��o�Yns�*SY/�rc z���eߚ���_L��`�'�x��O|���?�o}���Z�O��͆M�p�K�E&����~w�t[vw�d���=���۰�LY8��cR�	��0�Q�X�ct{����x����3N6 w�m��v�4#D]�� �ܥ`��-�Q�� �P8�w��V��Ť�c�4��'��n.���N);b��`�ȶK��ۄ����xm���c��a������ܩu��U�������׸W����`A�W��.*	D�Q!�jʅj�ME\����>��z�`]Ǯ�|ۻ�~���z���W(�����uL�k.������	�>*��� \�U=m�Sn�o~'����'+Q��n.���G���S�jm�@ʸ��3C�� z�E�~�ڭ�n����~��o_{��܍�Ə���}��W7��_r����:��i��Kɺ��	�>����ic[��Zp�B)�2�,���o~��![��!���t�ث�����ԭ��z rQ���[�N��� v�Zn��=f~^h��8�E�疂�Y�R]��1v�*���/-K��qQ1��[�;����i����NϤ5b�O���߉��~����>��Y77I���Tw����w���vׅ&�`W%��E��	�-��B,�e�!��F�F�|zqx�"���.������7��O�[y�n�TS4w�Ly9>�T�V�	,5��Z��,C6v�!��!�0z衇6	�cM�9O$��O)0�)ii|:|h���v�)Wj�>ǩ*��:���J)�{���&H7�����A�L���'f���i��_=�[n�e����
³�^�e}��]��ĚK�:�:����n��&R�� �Zp�a<�`�Y�qU��µ~���1+LP\�,��R��-α��v��|�iH���+���&�`����O�
�2��0����F�00ǚۣ��z�:���@n�|�{�7�k��r��[	v�:�Jjl�"�X��mܾ}�7��1Թ�<i�b�\��]ợ�X�g�����w�4�u���?��P(�����d�*nD�k��%���92<��IOY�Rr*��Y����qsi��>�`vR�KZ#���ua��&�0�R���o����/�|o��	�[x���7x�x�}v-Ȑ���0µ[p�SW)������Td�%X%��r	�d�1��s�.s�y�'�􉦐��˿�ˏ�A��w�����{�o�}C��x��9$|k�nʣY2���iGe�ENה�-�k��Ä�z'�X2��	p���^B@�0�d�w�+�O�s7�o�QЏ��Mb���
��E_P �`�@��On<��Sˉ��WZ/���`c�����h��@T _���Xt�~X`����<&�����l����,^�	l�a���|ra��3�swK�?��f��@�����m�!�$��nyӬe�L>�2,�.½��U��7�z���u���@z}���������k,y���9�ᇍ�H��}}��UR����I>�9�������L��=/4�ݘ�17�RBֹ�}Y_�`��\��T �N(�V�x���7���ʭ[o����?|������6�������5����֥�1�Wk�ʋ<J_��ǹ���i-��B��Ոգ�Xp�x��S��������7�s��	O|�5�����i� ���ʆ�:l6�9��Վ�G��NW0/@�@�) pL_�1G���uֱ��)^���s�m�5Ӓ�1�f��p�����ed�ھvf��]Z?��O-�)���	O�Iz�)%��g����6��P&�y�^��Mhs�^��t�m��t��eT��Ipk��w�e�����O�g�NZ�}��P���l��r��@�s}����Ͻ7Q�^3���?T��c�=�Iq|{� ��Ia՜S7�K&I�.�XԒb){2x�G+���a���k��d�\�P����dU"xwM�u��s����f'<u�n�ᆏ�}ꩧ6	M��AU��a1�џVXꥫ��Y+��Ȳ�*�W��
h47����!-,iݰD��Jݻ�r�-��+w2�7Z���<hq[��{+n�jp��/b��
��K�>/])|O?�|�̓p�q��&p�e��\P�;�g����Z�z׮��_���=���Z2�r3�V.�
��������S�nY����V;tT�rO-��2	���5a$O���e�Ǫ��h��
�+���_X�w�<��B�,𝝔\x�i+2`r�]d����4&�z�K���uܶ�c�n�Zs�UH�Gs�c�ê���2D�N��`-7�NzS����'Z�.7jk�f����,���Ҕ��o�մtWE0��(/2�ݹ�!K=$7{��?csm�_�:97�ŕ���M E� άP�F�L��������v��MF�jX�crY��h�ih}� �@*N��T����yA�#<ι�g�r̘�GG���{�'{��w��Xi�@�����_�җ��XB��M�A��{�����_��O��?8�W�W��Y�d%6�~�%*� <:�3@��Y�-�?���2��%M���*��+M�D�1k��u���TaZAH�w��IL2���iM��M��;ː�֓��k�*\�k6n8r�� l�w��㷟~��& o�) ۸��|�\x��i������&����ھ�	��?��24E�>R1H����t�zo�a�}y���7����%E�}O{��۹&��Gc�:�+��cU,z�\w��S�V�Xu��U:�^�뀈�k�vT�3�7w�ˋoƖ�2y3NܲW�7��<��~��D�y[��s䅻BȦ������Y��9����4p��p]Oc�\hL�O�����M�mX�m�^��b-�Zu�Rm�<hL��{�G�;��_O?�䓧��Hc�-P��+�5�i��ɑ�0��Ws�OHJ���S����ud��Zii���|��@*c}p��@J����c�X�X�C�(��c���n�੏c�0�n�)��f �2��g
�,� #�����@fq�,�
�

+�Z�{B2�
��Xu�u�h	N�%���ׄ�e��ƶ�4�[��on������
�G�=����ԟ���L���V�Ū�?��q��N�	�Z*��]�vܙ�5�̙3��ݧɌe�0 �	���.�f)��'�L(��X�\��8��h�������8WݧG�.���SD\�ʚ�9�-V�q��s3�J,��W��������+�Rk�J"����I���Z�;�q>�b��َ���8�/wÿ�M=~̪,rg=�H�F������ �u�d4�c�<���\z����m�>u�w~$1�/��!d����0�R��2����Z�ݭ~��ǆ��#�5ٴǋ��h�b
X�Eg�h43�sؕ��<�:��,�nL�%q��{��%c�M�l��XhEIM�A��n�������P��)�:�&$��9 �?��O��t�@�*�I�#�v�e�
��νF��	p	�̒M�[���2��)�D�i��c6���/�n�{�����{�lmڲ̛�y� �����n���\�5ϜisnV�O�+���'?�	�7�3�>���&Y�?_��X
L�D�p�>ã�_�(�r������w|���ݴm�c�Σ8��O�Q�����T�j��L�T���TJk99��������}x%������y�g�У�/VW�rBO��|�!V�^��$2Ø���BUQYW���z����� 7���� ���,8�E[�/�!"Z�b����܀����~��S_��W?R���a�a�&d���dH����b��0"x'<�yx�x�	�}���'�%kD��LY�S��<j��C�\<"���Dv�߀:�7���F ������D�O��^'����n�tة�n��#�0=��8�ۦl�M�0��B0��  �;��F����W~g|j�ɱEH��w+�Ʈ�{͹@$����"(��߻1�*]�-s�:���z�[��]�j��t�0.X��R
�'����9o�
%��I�����\[w�Ɇ���v�Y&�6w��lQH���&��?nB�n-�3k\�y㌡�{���"=f!߭U7Ǩ�=e���^�ʇ������ѩ�u�;�L���҂k<_�탘�7�|�j��w>�V��}�{C#s��`ns�9b)4��؟�|�ϯq��$&��_��*+T�{^�1�:FS���c�Gd����������7K�!��'��?��2�[��,h��Ź�������Xr�#!\�:������~ �RC��Pf�H�`ˋ>�
�U�3��s���[Bu�m|�<�I���a��5��-�X���c� v� ���Qƺ�Q��[�u�����(5@?���NdK@����`��#�x����8���r�l(����V�G��N{�����\�R�C����Z�a�ѷ�g��(h���V�$�����ߺXn����܀��x��&0�1_���՘�R�c��On'�(P�}5��빰���~P;����e���cY��RH��������<�b���sp�����{i���\����������jkkOy��>��&�R2���X۔U����g�����E8�V�[����+��i��-�7ݴ����~��Lx�?u�:g �Aϔv8�2�(�_@���Z|ki>)ﻊ��l�v���W�q?)��߮}��d�2}BL�Z�F 8��SCH �B�a���xp��_���z���\'m<so[���j��>2���3�U7��ì2�y��'&���[��B)��ʳ w�W�g�ο�����a�}v��_,��M�
``���m@����E+j�����Tc�˖a��-�1���H��@�a�	t� a0�P-�I����d��� '� (�yc п��sz4�C=0��f�Є�uk��.�Ӫ
^��Rв����@s ��.^ġ+�'�U�r��_��a"/ۘ��̢�V���Y��:cYis����nY-�cDp;瞦Tｉ ��𝅺!�;���!!(Zۗ��Z��g��cex��`��Bs��- \�z:��:�(hS�ث�d���~P�c2ê;��i��o ��6<%���?�)5n�%��3C����<�3��s(m����K�J;��]�8���S��s�k��zcY���wcs�&�́LŨƺ�������|EN�SD��0lN������f6o���{���������;��C6���I �͘W�������e�Lb���)Ga�F���P;������ͯ̢�CŶ'z�Ez���-f=P�_{������?Y����g?��2Fs?%�0ƪ�g�������7�x�i���|(��~5���` n��}�+�W���J�}n	M�X�;w�����=�У9 �'<��\���ĺ !ˀ���5]��Y�z���]f0m`���e� �b��0c�qh鎱N.Ǩ���H�c�ZFu�y�c��|y����'���Vk�=$26��6�*VkK�s�+-�j�����H۬ s�q4u�]��������N	�����z�aOFV��-�]5oz}1�z���/�?eVϠR�v��u�9P�C��^^xC6o���}�'60"�n����d�U҃�!<Y�<ɿ�B&�p��X�S��X��c ���hE�{U��s>�8J0�����Zr�2�����/��L��E��}�Q��DR��D��������?�@�05Bhx�9 ��/�`7���:+��ك��<��y(s�=�|�O����_�f�_�2�-}�ʛ�Tw�*���) ��n�a2��w�v� ���� ���׾60���2�T@����\��2������_��__� �����i�$����Bi�Ϙ���u�pxȝk���TMú��cV-�=!2v�J{uE������Alfk�L0��v `�m�[rm,�xt��b�*4���<&�����ܑr�˿}NIZL��h�����L(�������,�������vA�
SHp�	c� õ�A����M��El]e�
P�5e��}?զ�T��q?hU��@��n�@̰)G���v��i�"��Z���sU�W,�`l�s��������~��d����|�_l ���[ڮL/e��9��,�"���E�a���)��B����Ei	�z�s�cJ��|�}���Cu>�,�����Z���;~��2�3NCc�d,s�� ��7���n�m�;��jX��>��Dcm5��#�<r���&�2���.��z)�o��+6�������_��6�6����4��O�n�u�֕?�ȇ1p/��zM��h�	g|ǂ�b���}Y;�E��4�S��N���t|;��6�5ƺ�	��FT���![�0q�L�H-p�6���[�*�O��E��"(j�¤P�+��,��)ޙ�~�|�P���O�W�/�X����W�l��ii7����p�����r�v�l���\<"��)~���>�ZH%ݸ�k�m������}�	���!<���a,f_g�\lCZ�l���ܹƅ�~E��
D�����9JS�u���O��`�w�nh���okl��s��$��v��\\�V�-ǔ��X=Dk�q�Y�խ�u(���ԧ������'����kƟ�ٟ]�5cg{���ֺ�m.l�
���=�g�oL�vRerw��-#�>+�*�\s(�t�e�Q ?��~��2�K� ��U
���V-�sU�Tz5�W(�B�u��ֺ6okr�� x���Ț�/��/���`�ַ��%���ݙ믿�X�3m��@��s�:p�^x����־-<��
|�%$�P�$��\'�U����c��| �ɫ�yu�x�o��9ا�>�x���{,�c���YG��E��w�� a�5KK��X8�Mp��cr�F;~0���{_���o���=Х�w{�{ؖA�[8}%�RX����%�����!�kc.���$�9����)��p���"༆�Q'Fm�~�0�-_�p3���/c�̨�m3�>o|��d.(����ih�])��KL%O����i}Q#�"�%w�zO;�d㗻�Z��6!��2-�3�N�Mr��Љ����oG�� � j�rα��ڭ�'y�'D����5k[�
������s ���T���V-Vy�VZyM�R��|�52Άqy@����[��O4�q_����r�-��f��g?�l���F� Wh�]�Z�0C/�>i]Dy0��aAʂ������[oo��ǋ!VAp#Ӵ&2�t�W��:�~o���]o�4��x�$G~��3,��U"/�d�ES@^~��lc��[�Xs��t� �����-^�i[��~�'�k�~������◆�05�# j��a�0�'��ny6���L?Y�*��axvx��A�����<�>I��*�]�M��t��.�u��D:���}&=��j����7�uҴ���t�B- sh�m�������{��gN����[��g�B�R.�@��u�8����5��8n�@�L�߆ypw	��`W�18�Zz��H�b;עV��s S=W˫u��u>�R�<wc|��
@�}j<]&ayΎŭC���w}�6���1v��F'�p��Y֥����i�
����rHp�b��-k�V�#��*�w�̙��[�Ƭ��.����j��h��ϔ㘯�6����j���i�L>4TK�3.H�^ש�
�����v;�O��Og�\8���i�Ĳ�h4ٽ���ɶP�sα+a���\�\�R��|Cn���HBY
��U�-��GJ����R���Ptv	��E��<����+EmmP9�9^SJܔr3g������uy���<I�O�Y�J^�*��y�Z6%��+@k�U�#Ɓ�U�Ck6 �㚲Ex�V�[�?N`�m�k��������.�O6>9�>�ǻ���؁��I�\&h�X���6.��� ��O.K��[�Gτ��-o��y�V���˄ͽaen@ݒ��7���hY[�;���i2K�5o�"dU����=�K`�ߺ���:Ӯq�w�����¢K��6�y��`� �Z��6�	a�X1��3��r�5(%P�b�?��2LZ��K��Y��>��U��Ǽ��ر1�W�zW�&@�/�ܼ�׽@r ��J.��
Y�/�0�z�Y��f�C�$�a<��dm\Z��;��e.��t��VNT�n\�$��!e��V��f\�]��W�r&���M=^�+�]��[�*_�A� �~��^c�r��*�9�c*j�N�|y;�u���_G�0�t���5qk��&C�����E��:�������{�<p����Y^�x�Ϸu�d�{�XD�����������H�k8�0�P�����C,�9�;�_ ��iY,�[��%cϬ��8��#Z�)���㕩��h�e@�[�/��/�iiG��߳f���8S�h��h�����(v?cG�Y��n-��6Y}��]�[���{i��;�<3���{���;�p�����?˲i�e���}����|��֯����9� N1�ּ_�79��XU���&�~ �� ��D��Ә���#N���t�w�.X*E�h�
��t�y���6~���m�߶!���� �K�>��g�����e� �گ �KײL� 7��s�)���r�YƂZ}7�a��ۥ����u�o(��v�,���b!q����tű�+]�,h��ڿ���MZ:-Af���"��p�@�q�
��mLu���SK//�mx�Ϛf�������o,؇��cs�$�������y� D�L���q�-ͱ�����:������kO��}��Z��I ��1�Ѱ�7���w�@C��:Ps����P��-p�N#�s�����C�. $���狋��H��6�;�Y��zh�5�bȿ���a�]�k�Ը� ;�	 n��u��I>[ΑZ�-��KSJ����1���S�m?e�;N��z�|����w(�B˸����ʋs���a��0�~���Mes+ˋx1b]{�[<�a�O]g�n�|����?�{vm�k!����[�l�o��仨�5�V{��9 }�<*�bpX��7�n<1�����M�r��:f=92EݫUS�SLQ���A< �@` mOg�R����f`�OK	),��q1t, ��Z��&!��ig�k�y�Rf��h�y���M{As��3��E5>J��������2���c��v��F&�i��ču�'����qs�ٳ�N-���ν��L��!�I�Z�r���^�ҥ�"�0��W^?�q�şڰ�����fܡ�Ѭ�`[�,�V	����B�-�� 6�`	r�_�wx��;C���~da@�1܁/��	��xf�h����~�~.�cמ{��y0���k�����!ߩ��2�T�Wp�ˣ�c���}jM�u��ok�j���3����t>�s�
&���U��ô��,�)�L 0xnm+@�y�a�`}5�(cv�U��>e�]W��-=Z�cSɭ�)ncF��ڕkO��jٵ����
�)����b=s�!�x�u�j:���N@����.�i�� c��
���ws�t�=6�>����&<#{i��oiI�\�mԋ�kd�L��ZC؅gz��؄��?�9�C��C�P����Sx�; �*��^�6�2x����3���"&m��mI�5����$
��|2a��-4��k��G}�L�{߲�=@�ﴁ�V0)�F�(�a~����(��2����k�"�0�s�N Y����@HK��HSx]�9�[���j��+�Y�|.��S���1Ԕ=�3���7(���.�%���C���;,Z&�T���,���f>sO���z�j��y2Vb6�8����F���j܇9�B��f.d����j����[��n��4ƛs�RZ�<�{��s��s�rZ�Q�fHB�W��3��^������z �U�X������XA��a��w���2쨮_��f5�T �<�ʰ�ü��]�n�e+Ð@�Ƿ��[-�zD��5~4�����1�U>�U����,�uM�;7W)l�\�G@W�A�c�!�>7̀��0�X+�$���;a��:c��#���X:^Z�-�Hq�[��-�s�L�\�$�5�ֈ-H�#̂�^g�9;���"yV~v=�3 \#%�3��2�9�l3�(sP�V�V��.��A]���1�]-�2��g7�x��z�c��w^�+ r��/~��ݺ�x��]�x�m���V1d��\-J_����}�Lc����&`�)��$��o�>�[�$����"S��}h��R�ke\�1����Њy�A����gLn�%��]�/�pKИV=�?��*���lU�KO�	J!�q��P�8����c��k�25z��m0I˘����}�j��:����ɣZ��	k5�����+D԰�Z�Å��
X�떒L��Ci��afR\^{�5���M)bc����;���b����glM�7��1�ɋ�j�1!�q]��"�1�*�ơg̮VSH~�qH�j�Q�.v�bNo\��tf��x�	��ǹ�y�2%�zN�/RƤ������v�4���ߙ� !���Rj��g*�e��c�� c�����͑U�u�z����׎�5ɷ��뮢�3
���}��_0�Jc�A�k����&�|�ӟ����Ro�-©�(e���k�bG|vC'���9�%�	T
�l�Ww��� \w�c>�{�۲��j���=~:�;h74j{�urAv����J�NG ��~x�@.�t�M7ݴ��KW@�Z݁D0�5t٠Y�K&m�-�~j��,C#��ro���Ztm�=s}α�*����b<�
"A �-/��%`��`�l�����M�WDo��٪Pk��"[A�:�k
t�ږ߻ 3�*+Lf�Z�Ұh���}�hp�eSkj�E�#]�7��-���p獕4Ԟ�ؘ=�qƉ�����3�*���6���E�V{HA{����<�'�,	���h����E��� N)���}/4��wKs��\�Y����\��;<cj]@�b����P&;r��Ӱ�Tʪa�&��w��X�$@h�n�TC����,��p�� C��}+`�7�:��d�?�H�Ҭ~3��O��	j�ڐ@{�����^���[�Mk�N�A�;B�T���Ǽ�F�O`K~�~���#�9V�����~f(��:�.��Z+����id�o�!P*p����ՍZ�;�y6��<�4�-�ã�H�d�/����x[�95�c�z���މ�}���Ǭ��U�
*h0Αc�X-�"Wk�;�Ȥf���eMYC�.�t�U2��v(Rk�d��dr�LT�Ze%�Ƣ@&# �,�����q5!� � �{�e��0g�[5�s@c�xaޣ�׳T+a=~��{�����KA���$��E���u�	������g��ڞ�.�Ǔ� ���E}�o��ƿ����p��彳�R�P��x9�v.pi�R���]�.�#4y�iP(i#�m��:@j�q��~�KA���SV׵b�Y�V��n��ւz�g�xzǒT��f���6�c��U��}����z�e���xw�w!�T��Aw��p�����؛���S����	��K����e<��������-�K�x&���;�P�_��:�q�7�]o�3�d�����'e]��� )C����`��k����Ǉʙ��2�(���.�5.7�<����C�+b��O��|-+h��C�h��-�3	�MIX��aZ��&�LF)0��1C��H����� Q�~����������*F�j��Y� ��t �)Ls�w�L��X4$���f
ju26���4�#�R���MB����� �j�;�V	A����0L0�Ɯ�����`hH|�f(h6�W ���56ns�ZVigS��nr�	�
8S��@) ~��o7ξuv�rZ�#oI�{����^7ϭa'k.��sν;��.$�L�W����y%c���aZy�����"����~��!i���\�7K��5s7��B�~�\et��6v�U���~��A/�n츱����e����Jx�0���*�����m�ݩ�{������6�|t�T��Cm\��-C��Vr�,)|6s�a��,�٫P�[�{ w,�z�{|�M��1p���ͻ�5*�q��$B���Ě�����u���@�1���9��h�0�&�2��`�8r1�f��#�	�G����r���-�3�X�RÄ8�Dk��P��,#������9Rz^j�̱1�� S20?̓z��[A?&`{��Qi9u�{�>�΢�KFK)���2��sQVcXL݉�2[|g���JNZ�\�.�O~�V�i���9P
�a����,K]0�`@�CZz� ��"n�M@�K�q9��y�z2e=�_�0I!;Ơc��P4�G=��1��E����W�^Kk����P��ꂞ1��`���.�R�	Y� -�W]yՠU�sG��V��=�b�>��y����/�m)�g.K�\��^
���f{�j^���:wVͩ��[��� �
p�_��5����uC���@!�kjL-�R����y7&����@��o���r��(�dk����� 	��0t0����P*yi�q��zs�%ed��{���H0��ܣ�
e=�6d_ƥ��;����ʆO0�0�Mk�բ���16q�]�A�)=$@��mQyW��2^��h�0L�j!��R�����)C!�)7J��- W�5�Z9B+uV)��ߣ\[�{�
���%��!o��J�T��B V5��L^�c�����
��@���/X�U�i����l�������uM���2��Q-R�N0���Y�o<3��]PT0̮5�Y�1��k���҈����}z�q�T����\iL���UWK�� b,���P"��;��1+�|g,b��ڞ���x?�WzO/� � �����ͫ�Mˀs@���%C��:s�_�x��G�p���b]��A҇�Js��n�Y?Ͻ^���~+$=+��y?s)���k��l_\��
3'�\�(?��؆lG�����BP�IpY�)ۙ�c�c&�����q�{�����Tx9ToY-��i̺�}]��~��U��z�ک��C�׏�V<b���Qnp�_q����\�c�eC��$���X&�gC&T��
0�}e����Ng��F<����kP�b�2{���H��Q�u��3N�����JK���-�7{2�P`�qn�k"�&p�.V$��;�x���F ���uM<C@XF)���VO�@>/m�zO{B���|����Z�y&�"ޙ ���v!�x�m��a��[��\[s�9����,Q�ڢ 3 ��e�ԆUR����c�:�Z�{�v�k=aG���޹(�����m�T�\�6���L���ڊ~�b�$���"�J�<-s�8v]�Z������*]J�X��AX�WQ���������M�$ݞ*o鵐gs����K~������Y=^������	 �j¦���t5�g q��fn��B	�5ai��ћk=�X��~��)cBZo��c��=�E��z��]��ozX�~��!���\º�ڑ<����{� W#Z*B~�X��%{׍�ʓV��F(�z�`0/�<�c��a��i��R^�J�����1�;���f���؞��r 5R�@k��j��n�?>�Gw� �f�q L�����{lM��^w�ȸM�1h\�D��pm��i7�Z�#��qf�.�H�3��n��ߦ�gEYW8�@w�n��Z|{��	Ț�6��	��geE�4j���n��0�4\�¶�(�H.��0�E���҂�ǒ\��l,�G넠\+��:|�k�'>ÿ&�X~F����
��ؼߴ[�0�t���1�u^�ݫڳ�:��B�Q�뺐��V�LN~�j�)�*�ڶqh��+۔�Yy8�i~�xA����� � ���$~p��#?��C��|�ͱ���19^�n��[��Uu�{����9j�1�O���� X��@�
T�º��A�er�f&�����W+�@u�:�,������+���h�|������~W�!�	���d�����C��I+����7�WAl�W!�� 2�0������k�0�!`QƁ����Y��8����A��Z�7Kz�,0��Z�u``�9�H���A��2a��/����.aPx���uh���y~�^���jq�n&��H��w�^[{�:���j�%�2P�a���/X2��բ���{�q^.LW(o�.σ�,�)���W��W�%{(��l��.0c�*`z�܏��`Z��Xd���}ʠu�u������]o��v�"��cƄU}�;fꜩ��:/_Ryw�x=�P5a&]�Χt�.3�7�������~�����_/A�����m�8�p�ܫ1�*�����
7r �ry(�xKx�j����U,�M;���~�͙s��������S�dZ�5LY��oq���c5�H1����S4��5�T�\'h��r�y1�7֕��<^�
�!�`*�ܢ!�����w��*�����^����1�;��k��Z�\(5��T��5Lz���z̈́@cy�0��2C֖���7��&亶	�~Z�`T���	�Ծ��W-�� G�-h��j���h�s���t�*Ȓ����c��kۥ���%o����d����� ˟��B ��n�g�h����#O�H��Y���[�x�H���`@a�e㼆°�nSPf;�X*�w+��φId��E�E}��Q�_G!�C=}
ȍ)Hp��wo�{�z\�Z4r�s����g��ڸ
����;^��1� q��!���v�L���,���6,���ݹ+�X-x�ĵ��f��R�Ʊrn�M�1T!��_��Y��p�N��9�M |�z�S`�7Nc4GٛC���9�zl-�J��:%�~�%1��WO�dMzR>k���Θ�6�܂�M�m۲�dz+���X�A-��	f�N�4�i�� r�����׿����'����*�h��M������c��9.��{jK�KQKr�dc^4��Vw����U{tg`t��ѕ��Y��
D��:xn!,`�}U�J+�}��{�y��~��`�❞���ɍ	��B>�}י<�I
�$c�!����u1Z�gY�`�s�Bo����o&(�nl�֪��N@��u�j̡�i�'�,c�2�a��
ڪRiU��^�AO�JS`wε�oS�sn�*�]eh���V���c��8Q��-���yǶep&Kɇ\-f^���`�	^���ʦ���y��b�E5�&v�K�8�Cub*��0� DO�����)Jc��s*��çc4�4LC����~��[C�S���oe~ ��,<�̪4��jNO���n&��3�3��!�C�b����_�Z���򳊥���6�o��^�V�Vyvɫ(��jU=��J�]��m[U�6l��� ���ki�LWn����ok�-�F�2�p/��fZ�����^���� �e��ZXƯ��~�Գ:�>Ͻ�^ۓ4��~��M:�Tǀ��㎀�җ�4�@�?H���#_՚���;���x��U�� J��X]�WUA������W_u�2��V0+֫y��:ƃV1%��r��X��1��|:�$���X�悔��� z���]5���`γ[�Q����EG���j� 7ݴ*rP��
:�d)�z�\��v��Tv05��y��3IZ�`���W�^��Ϣe���|�Ky*�N�kP��+?���ң��ڒg��<|�����~��e�3e�%(c`yO�q�<��U����VÜ!�&��k��X��9����gwX�� V�
�K�O�圩���:�������qI�3��x
%<'l
��Z����|oi��2����(�r�05&��Z��{R��ݘ���.!���	2�X����k2��e`?��hXWS��ϵ�Ρ)�0%���V�S �����z�&<�l)�Y��Ex��f��hߧ;R^q>�%>hqͤ�e���JK�}�;���\Kw��Q"�]��YT��?����ui�u�u�.�s��zy��Sƀ�h������%w�V��6]��aՃ�U:\��'��u˹�@����3�$x��|��Bf�S�������k��Gp��*�wC����ºg���Ķ��l7�*k�S��xc�ܟ��)���a��ᜪ�8Ch�ܘ�r�S+&��_C���V�r���TK2f�y>��ۥq$��c�ܣ*�o��W]����ܶJG��~/*���q�� �B�jͩ����qZ�&��1N,��J�Y�������ư��,��e*A1���n�Mhk֥� �Z��8��u���cV��^;�����<���RqZ6K�<5,�G�-�"->YuC�ՃPی�	�]iRCυ8]�	P� {w{�6wS�:�m�yL�4��2V���3���3���9��M);�w�"�u^�s�|Q����{���vL�/ϫ`����2���֬9�u	�_&Q)33>PS�O�[�g=�L�J6a��=�醭돞���.��˰$Ꞛ4��k��ԥ񒆶cK���φ�J/���}��<��U��/�~P5|A��r�F�u��fND^�ы+��R�&��s�[��a����9ú3���;af_�^����P�mNR{�K�p��L�<� �k]u�nij�L=��T�gL`ֿ�y��&B1�!I����r1v+D�_c|e��=g�J�+�4/��ք3K�	B������Ρ:>�@�s�1p;6�c �Ǭ��5�m��U�:63+���~����d8��cӝ
	.��s˾Z,Ew�4-F޻Η�bl�$�� �\K^K��^�!��������g+J@��x���w�*�X�'�?+�Q����S�V��U4u�z�x�חZ9��ȹ^�-�醭�5.�:��"��{�i����2')˗��>���I=XxT��J����n2����L��So
$ ��g�L�%-�s߳�!k���r��
�,�8�&Dp��C��돎�?t#& ��(FF���XB�,�ՖYg����_���d�[ow��NM�~�z�%�ɬ�,]���
��g�����5>F@��㺔)d��s�o����S&bF��(j���79��uLL���(x��(����'�G�) ۺ��w��}\к w ��mVN� �@�t���#E�3r���o���a=H��0x0������AhΙ��˸��m
ZF�_�!�I��\�8c�:	U�h�?��`�Y)��`ء��e|�e�+���~�� xS��KGw�;@�]�_	WR��鏻����?�����e�[N6��Be�<�=���"�I��Gs�8�n�Xns���R9�2� )ۺ�waº��!k��p��7.�}���	"V3b�e���v���?�
�J>,7jq ��G�5�E�yDq�Sy���
|Csw7斷ek��5��;��
��%/��E��R4G�ì��;uo���m�؄1�+��	>c�Ҽ^�W�=�gz��"Ĭg	q�̃(7Q02e��d|}��;�� n���{�2!��p��,�:�����wt����#���N�&��-�:�>�b�l[X�4��>iiv�sۦ8����M����;^��`�^��v|����
��P���&c_�̪R�Ŭ�܋���g:X������O�-�hI�z6 Q:"������]K]��){��e)�k����ݗ����o1�Q����ʨ� ���t~�xDl�M)>gt�2du���5Bݕ��b� \�pQ � �`1ƭ��|������(.�Mp}�t_��әK���0��䊠�_�iB������kA短�P�=�}��n�1ت�\���o=;{.�u]��f�z�ʉ8
�D�'Y[\#��@x�Sߤ(��̔1N��z�S��u�7��;���x��R��Ys*�Q�}LQ6Ib�-�����я{F?�ϡ�g�����3<�Ǘ�Z�=ul]�j�H8�:mBs�V6^�xKћz>�>Y�/1-糬�.6�MP���"���:�!��W��c���\K���V���Z�.I/���ⷿ���ͷ��x��`L&���M{K������u!ۻ��\�Ξ��u�d-!x w��v�<�����D�,Zwﻼ����W�U�VV�DXc�D�Ն���gZ�|<zj$�[o�uq˭{Aɬ�����b��߁�[�}wK�5���T@��.�:P�����,�<�Q����=�{���zY9�s �ኩq��b�&F0�%ϝ����z�񸻨x;�
o|���/_-v��A�����V�e�jj<����߽E�؊�o]<E>�Gk0M�le������F���`�&�����ZSKK�T���z4�9Y�ƶ�����R�F�:u��� ����C@���� 4?��O��1
%W�X��z�*p+`]�?"��G%`�3��������1�������#L�E��������xV��62WZ x.�w�>#`�G���j���#s��"��F��ۊߍ.�Hp�0���Y�]8�������[)�4�*f��A���G� dߴ���r7�\W��?��ϫ�:�,��2�nF��es�i�k����4M�k4@iğ���cs���������|k��F�Z�����V�E�k�Gz}��u(*�\���lU �7ey�Y�|2�)+��w�S�|��2h�t�:�v��#�z �����X*�,�'o� �|[%�<�E#�V ��A1����	j��<�?&�'-�>���/���:�2H1�	�@�����2�c�~<�,e p.���S�X�x]d��Ӵy���i�S�7�F��)%!�����g�R����À�p}Y�[�q�I�kyZI�#Jp��8�1�}���h�᐀����c9�I�O�3�����ݦ ���5�{�d�6�}s�?���d�p���޵��� PK�yg#y�1�<�ȭ�뒏�,f(k��v�q4��L���J-�#�n����4�����)����3�i�����ɮ������L]��6�w4����h���,�[��ԊuaY���ci��l9��&�%R���<v�#����i�HG�I�@��%s.s�v����U�n��`�晠�����p4z=
�9m�6����ʏ<0fK��7��4 @�+�Y�-�]ds��rB�f�$�A) ��<�#�1 MF���V�V+!Z!��_�k���ֳ�Dp;ĭK>N�2�)Q>γ8���{�P��+���M`�M�\��8�������gΑ�ν��>�7z�����kȩ{�;������Yj�w6c��ο�:��T�;X�A�4��X�� !N�u)2�E�(��e����JL��G�֠�Z��{ɸ}�0Ϲ�:� ˾�{O���V�u���ٻ��dF�3��3F�rkn�Po,M)��Q��ؔ���{�0�M�:����\�,���5{>s�Szi�G_t���l� ���q���Qc^eh.��K9s�a��"w뱎�c�L	������v���U��2�Zs,GSc2*'����rk��@n��Z�j��Ͱe�QTc�X��,�Ǫ��9��xcp� ө�_���ZG��u�%H"c�&r뽷�q��SB�@�>�������<A���CK������t���U����Kh��m+(���N��t\��]�� G��@Ɨk[V ��TQk)̏{ ����t� �9s.�L��
�� xj������S
aV�V�=������b��� ���\
�7ua쳥:J#�Ey�[ߌB��!�-�O��0~�d�!=��T����12u���:�1&�pT=P��=қ��kMS�<*
�;Uޔ����~�U:Zrv�6Ω�j�B}TxL��l�w��X�"�����ZL%c��jdۦ�>�ҨI�e�����D�oj�,�*І�C�-�v��=t��m�FVY����q�K�i�� KO8��mE����=��g�� e+�Qk����Q�B��e��e.O�{F�m�Ys������^���d�Q�dq%���#2��̟]NV>�b��zp7�zW�Ȩ���{�����t}��L �S�)�1Շ#<1Z��Xu$h#2:�e�>Hy�����`�'���G�cFڷś��#_����#��z��m1�f��Tc�� v~6�ze�:��Tf�rf�wF�%˽�	�9V(��FS�jǌZ�@��M�ko|���֘��D�Y���[��O�,�K7\�[���-��D����������"�'�$���H������̀��5�U,ޖB�SR����
s���u�so(�i���;�sh�����%1��l-�� L�B�KKF��"R��F�.u��Ҿ�M��]n���4\��������� 4}��l�7��x�4�1�~r?��<�sj*�WF��2���[|�����S�"��=�|�i�N)S�����g������s�>sPN���^�>�����F�A ����<�6{e�w�ꨌi�������3`1����H�J��\�ЍQ�1��h=b�M1�)j1�V;b��Xܖq���{H{� �x�
e8aA�bI�w��9�+�ܩ{G���g�90�9�[��r����=�ID{r��|_����D\DX����X
��Xf+�:΅�\����>�*���[�������v����?< ������7ް�f�߬(�?x��-�f���Vf|3�_K)��"��)�y�eG�g�v~�ޛ=;�}=�&��kz�8�WF�n� kā�2��b=��>�(d����\�I��h -�ߣ�g�t�=?
�쾫A>P���Ѳ��%s�+��D���z������e�.�������d�RF�������峥�f�qdL���k��sܭȫݨ 4Q"|���}�s����7Jw�u��c��
����%����(@�V���;��Jʐ[�y_����V��)�B7��xm����&�n����٩z]�Xǋ�V��o��8�"O��)��%�Y�qc	���X����;�s��7�̹�N)'��8de�ݩ{[�i�Gfc�w�&�ί%]�p���\��9`eJ�n��m���|*�]��JFDx}�6yZY.��S�&^���e�|t�ε�x�^���Ҩ+�]LR��O�^��\l��{b}�-&9Uߌgd��2�/;�󜩞�J�ۀV�Y��>�ʘ\�:NZ)����X�0�<�����EW�-� X�f�M�{>c,�X�}�[��ne��~ZG���}�cɮ�ο���5ėv},z��3_w_�ȾG��&����/>k*�e��S�ɏO�܌���}H������G�`���u��^����ӄASi�eZ՚`S d�*6�ᎂ?7G���$�-����zFܶ��y[&�z�����j���[��+���?�%l��GW����	�i�J�"ϝ��N;��m�	a�L�(�-�_�wER J����Q{ T����yQY�V�� \�?淮׮X���_���F��@.Q���I�	�*�*@X�i�>D���˃ ��}g/��@�O�wxS����ǽ@�X-��F�#$�
���6�R>�W�s_��<��3�r�2���L)�-��������{��r��.��?�8�>�i��7�֥����c`�<���ؤ��l1�)�u�Ȅ�i�������n4O��Ϲ�+����2�9�� Lxn�{GvF�6��[�2�Y?�<-��U���=J�S�*��?w�=����I�1�nOI�����i)��/���I}LF���G?��
H�[�hw+~4ᳬ���5˓�oX�9 Ǳ���M�؃�ܿW����{`���z���#��:�=�v����H�D����*A��,.yڈ���(h���b�2G`��߅{[i�zԒs�c- ���k͕�ѪW|V�}b=3ed.��ҔQiJ>��f
'Lɼ^��[�l]������hm)���=��4�Yg��]ӣ9`j��� �#S�.
�)�7:y�&z���V��3�F�ז0����0U/�c���.t�mQ�n*�b�� -��]Zee ޯ�{$O�[��~�������'*����G>R-� Z��V X�m��DOM���i<�z��l���
 ���m���.��q����ڵN[������{h'-�|��6���[훑�s ���DY���W�\�Zb�u�H�W��on�65��8-P٣��o��͑qz{�4��s���2F�OlӬ}3�s5��u1�:�`S �*�p���/�V�� ii�����ѐZ`��Ȭ��e�,�^�ѲF&�p;���u��������}�j+?����*����=Oi��X�m���:��TL�=�*�uk>fǢE �A^��8@���������8긬�d? @yb��E1Z���X] �:� ���z/Hou�ͷԬ X�uM�n�����{�Y���?_��꫋������7 @��\��g�F]Tl�X���-{q7/�[q3�'{���j�{�)�4��`6o[׸$�L��Qޝ㑱�3m�zϘ��z�ų�Z<qʀ7g��UN�ʽV��d<}Ӷ�����Qkl	�)���A�k��{u���HCO��ӨF4�u b �(
�,���٪�6'z�9��u�S�"H�s>?z���&������w�A#h��d9H�A��wd:#m��]�.��j����m�6�u�\��{��P���@ Vnw�}w�����;[Yj	(T�ܽ��}ɛs����S\W��2p���<V̑�mϲ= [�@7�WVܟ��g���ǋ�^{��\���6Vc�e8��}=�VKp��t��<�Ӧq=Y��]M�Q��B/n���0��G��[�&ʖ��#��������Ԛ�#�-���uO���[��C���znB#�o��B&�>�?-8�N��k����:�N�{V��p�d��/֧5O��඀E�Q#`m]j�޵� ���qD�16[�ix�Qzu؄Zu��m�ֶ)��q=֪sk��ǲ[�q�I�d|h������(�I��'�>�#��uj]�	��y��$��S�c5�3�zJ�.�0�f ׃;Ｓ~����{���Z���	��Yu�O5�p�;n������+��<��� 0�Ľ�l��ԍ,����>��rː%W�����ƾ��J��hD�:�G{���<V�),�J�+O��gv�s_c���(�W�o��"�m���;ʧ�ܝ�~��|��gu���we
���M���?w��(�מ��r�c٘����J�\��CSe�d`��Zϝ��\˽w��g�9�;2i�I#��:zJsr��=�a�(Y�[�a0niH����C��:c%�++�uM�.����M1�����%�5��m���b#4�St�$r �����T[���s�l.8����@�K-��#[Yp��+`Vm,`� a�6���+;^����Ņ���D�~�
��)�dQ���c{{0�@�r��r��@��������4��u˰�4p���\��o�A�x
4o������=�����7s院�w��ۡ�S��3<%Z��M��$4w��y��� � �M�'?�cV�m�ɑ�NQ6&{�U�ѱ�	��~˂�s8��l������:� i������g�Ѓǟ'`�������u-��`N���0�3��RZ��1���s�m�佱���Ub%�{�+��F��Ё��Q"���2l�z�=�{e�w��;Cwk"�g�$/k� ���x��
rnu�C�4=]��+@����r�}<��>!�-�����u׭@eU�Gu����o�+q1���p��W��;;;�+�L.
Fӷ��&��a����9`7*7�'�')�<ݛ�7�l��,�j�vp_c����)pڛG����O�|ۜq80GeX�MK��z�l\Gf�h�#���s��8F��p��}��r�'��gf�c�j�㱂���2U�Nuvv����4���l�D�0/?N�^��������ȌGڹ��u���9�pȮ�L8^x���X����˻�D�cI�G���MYp���"_��w�7��l��@0�w�(���,�� �t��2	0�L�|ׯ�=zl7�oY펅u�0 hn����c���!8ʳ(����>r��n*���@������T<2i����9�N��ҭ�4Yv����ӇqE9�t����\����:������|�z����c���<����5����Q��w��8���[
��X��|�@w��9���_��{T��ҔL���i�>GI�C�3|1�}|n����	��Ъ���@�T}z�׏��ۤ��b�Y�L͑߭@�^��0�~F��ۏMi���Q��u����Sz�����7�KG/�K��K����n>���6�l�;e6�:�WD0(��>�� �-�:�������a G�6�u�r)rqa��k����y�.���w���p�;�a���uOS�����]�`W��K�~z�-K��s�uy	vu�1�p�f3@�ʓ� <�*�}AuPYr_�ۂ@0��U"��L��(Sv0jg���&��������o��Α��;��؛>OZ��|�K��#W���1�w�;;��^��X����P�����&���Ӳ����e�9#�%����)ʔ��w��2칍:v]�7�:JsPk L1胤��`DK� pr=�����l���o2����ȅ���E��:�q��KK��˛�tx̀5��AF�@����^Kr��{����,�����`)Yjfe���٩ W �ܵ�7τ@�x>T,�:GnY ���[:���o[��7�Z�[ -׉���Tg��d�������w }u=�����@+y{�VjC�����߲��� Ȧ:'�y�;`k)����\�c �g�]}�'�������X��o�z�S�gql�(�	�@��z�g�\�ߎ(��HqP�v�2���l|�gnz����ڽgN)(���u��^ό��-���^g��7�Uσۚ0~.��hJ�ؑgĲ��N�dL�Es�&��l�[�����%
�HYlɔ�Qƙ�8�1ѫ���g�kz4%��sڙ�.�.��f��{�&�{���֫�10�|�>��glK����|ƬG VB����m�}��'O�\eFГ�S�U�%a!uЏ� ,%�&�S:W�#� ���C�wU�X���@��3��|e�+�z�.���{�W� +@����R �6��tUW@?@�����g)_m*Э����~���OW߸\��6��=���X�igv�� ���򜷀fw���ee�����ϫ�2�  ��IDATm���F>�O�9=Z�X��"x�{���LF�hJ����M�w�\��Mj)�qLE��b1�c�#2*�wn{d
��,9�ze�{J��P�(�G*�#���u�H�S�8^�Mn���Ȟ��06��ޭ	���z9C�~�D���pv?�)��L1�6P��p��P>~���	���I�plϬl?�B<>;R({;��G�����/�ˑ꩕ 0X���
�n]��c�S��yJ����XX�=e���׾����?_���N�a���6Xyv	]�k���?V��_xq�ʫ�� ���7~�4���Ǘ�wp������7q� �o�=ճ|�ˤ@&��o��n���[߲hK�� �8�u���q�6��R(t�@��/�\]'t��4�P�i_�l=u�[T3>�{��k�O��Ñ��ҷy ��7��wd�c�շ������&�����d��3ų���gTP306%��X����Z|����Evm�?6��G��?׳
��DSĲc��6��):=�F�x����&�Jk��'3 �u�6*��X&p{�_&�#���-�����D#�BY="E���&����l_ʍ>�Y=��悈���߾�P��,!��MISc4����#¥E-p;5�d��C�uK����-Xש{���x�п(����J*����~����>��j�H� (AGn��`��,��/��x�?��O�U_S�!��q
0s0���E߽�:y�����s�]q�p"�N�M�bʈ��|�����Nu=���xq+5sT���bѕ�X�Y���V�q���\��7�?�Ca�c��iV=k[��#{���������,���^s�#�� �-4�z�(^�Q�EY���3���9�B�O6��y}�*3ٜ���)�29{^��|�-c�S�*��-j)3S�d���k��mu��6)g
�DГ]ߛL1�;c����F)YG��}kcp���7�ݏ1�3�~z�Y�C�0�$��%�h�q�L3w�m<S�F�r������_tQ�j%�*��ì��ɩ%�����x��YV�@������W�����?]]d�T9���f���&KZn�V�д�� �,��p���ZAۻ���M��[�U�E����	��b���Q�br��OY�[o���cy%ˀg��1�<��^�\]�v��[�Wk�rW1����P82A�O�xi_����A�?q����r����;O��Gp�곃���?7;h��s�wv^�ݭ���)��L�8yY�:e`7��M&z���5�z4z�զS��E��(͝S-�ǯ�<���5Z��w� Z�6#& +K'� ��{8�!� p�y|}���[�F��2A�q`ƒ�o��r.K��p>�.����$� �j�.�	�
�'���� {��6��@nk�9(t�XI}�/��[�e��/y�կ~�Zoe���|��nF�eV��I����
��nj�e���uL���.�1b��e�0ߣ¥h��g�U���U������/W�X�.גּ�,���Ǘ���9˴#��:��
�c���⥋��1����-����զ�y|í�Y� ǶyH�]�"�6����[|f
n�'S@8k�^�����rc[�}��U��(���㖒w���X����c�<�-���#u�gM���N�b~B|1}��'LL�@�*��og��ߐ���]�p�� ��J����xR�n>A���ش/F��i��HW
ő�oGs�S���{��1x��7q�Q��/Qf
fTt�sH�9|@���/U�[Yp�t\�E~V��&���9E��i�^>�*�`22}�(��(��!�=�8�wֆ��>V�bag5D�(WY�t�C+p�ౝ����8�[��r�S[	(�o�@C�ݯ�@�3�!���������s��*NJ�[���kҩ�Nގ�����R\z��M͛Md�Ј|o���pk�3���M�G_k��l�o���]��.S<�#�Q��2�;�fAo٤���`DqX��������Ͻ.��n���C-�?2h�w<��K��LL����$~h�@�!����=bܯ��y@	BE��r�#��I�ە0Ӓ�"��	2-�
�����D�����̨�ʬ��;�{�u�?�����W���`<�{n��nB����J��K� q}�R=���/~���*�L�[w_�߾� ��r~��_/~��ը;��}�lj���D1b0�EOi��=n�n	�)P�f-�,E@J!>ؚ+Jm��=y�dm�Gy��)hk�ʢ]��Hג�@�Yʂ���r��[�����6���� h���o��x��]�Ƽ���nz���Zx�+t�q����������Xκ�+ch�ʰֽY�-0)fdh�W�XD�(r���;۟�[�a%�-y�i��(�[�r�E��-�-c�\���s(��}���yvԺ#�oi�#-�� � 7ӒE2�պՕI�)�|P�~�d�o,Z����0�A0(_�vM=�&$ G]tA�R6e���e�m�Yq6e*=�V�>�D��!H�sfʏ ���m[c<S���`'m^ ��������ۿ���S@��(\\��]e�������3�<S�\�Ā?��	�ҽ�S��Ѿ�Ͽ�z�.{�hiU��?ܲ�"��r�S;˺-��E�p�?��C5���*��	������U�\=S W�������ϻ��W7�kY�{�\o�V{�F�o|�ֺ�Bһn�Y�/�2~�2�
��>�U�dQP��2.�A���E0� �y��S||���\�I�^�ec䠰FO񜺯W�^��)�gr��t�����(��;��5J��Li�칔1��M�/���-�w�K� ��9v:��q�LOM�Kp�Z�k
� �F�_}�Dw��SW	S��%L�,S�"�����l�N1�pɅ[#�í��,��r��@��<Ιף��ǔ2��G����OYl����/��oT�[6  m~�NyO��~q�ܹų�>[��$�t��  �y����ʓ�[O�����ՌO��/��ͣu=��u��/�P�-�q	A�T��:
"��� ���ԦrOP[I9Y�ҥO4�O)l�>�o�y��l��/������*����s%Z�I@j]��Q��������z�_f��?��d}���F&�/�0�q�-�!1��΃�xLD�J6�RÖ�����>����4�m)1��@���R�{�n�G��<wM��f���Q-�%b��;��y�[u��Z"���K6h���`��� ��H$�$�!��-� �D\�R��g%-�,gDh�y��C (C�D�-�ב��]��-k��.���~i����j���f��Li�s��^*�G
���?(F��r*
 �Ayn� ��̌ie�4�A��u�(.�!,��`��XY?���V_[eM���z��ow��Sl���K/-����.��_����2|G0_��7�cY4�ok% 
�ا�6��3^�]%bjŨ��o�-ܞV]�kG6ƅ�>s��x�+Q�G�wW;KA�R��V�,���[YZ:� W����pM?"P�U Ց��|�WG���&~W�2�}�׵�5*�83���uurY<"[Zc�U������Q�� ������Z�/�m���v����^�*��7��F]�ˌ��_@.nK��������m���rs�e|c�j�%o���gn�~#�Nᮩ2�x��yp��S@�u�_�꼹��=m����Xnd��fn] �\���?1.�������h���?+�&����T�u�jet��=k��\	-�(��IB�$�"��k�b6z��Q���T�GeȒ���]<H!�w쫩q�.�c��`2K���G._��-ud�f��#��y.,����Q��y�����M����`�����D��p����J(���[��?X���?���1�@�Ah�#�<г�x�em'��s�El���͗]i���7�ew���]J�@�H��O����@3���,m�����"���P?�\�w+}˻��sK��m	)/�n[�FX��Z�+2e.�Y�Ƕ�����8Ȩ7��NQ��w��;���潍P �ѯjov�ӷ*�Vf��C^�� �o�!�<���iD�?`��H �ȕ�`J��)�2��:o3o/�W��(*��R����L���OY�#rm��s��0hV�V]/�z��b�P�������"�<0�B���Q�Xo`*:-.��o�M��ș�"�?��K/�BBIװ��x�K1	B�$ ���t��K��zG	T	gиk_�I��٨R���9�%
��X�%S�!p�Xqc��(,��z��T�D����K�D}�~�ԧ>U�le�U���S�e�h�hx�� �\����U�Y
��(Xт��?o
z<��Hc�KvMd�=ᑍQ���1�����g� v�|�L����y��a�+��?��"�s}�Y�Y�`}똔Vs�%,�=�kӸ;�y:�eL��(|=��>A�h稔��k��{�ʜ��~f��Ϣ_\�R�㶂RA�s=
�H�Z+~�1�����{c9eL�����(�>�Ɠ�D��i����OJ�����_��+�����_5ؑ\�Χ��iT\��5�e�c?�R���Z��jc��2;5./����У(�3�6e�:�FNK��z�;c�r�[LfLE�V|h����s��}̿T-&^��^_&ԇzb1�����h�
�%�YB�K@ u`y	���EIzg_�"˗�@DEa�F-/=�}�" ���NT�����b���1�Bf��b��ƺa�ӹ�'O�ܶ�`�����D*KBGB��R��f��w�������W<��'��XV��2 �]�ʫ�1}�Y'c}�Fe�WO�&�9���|���'��R�x}!"Yq�������� ױ[��E�W��/:��9�����͍�>��N�{�mJ١S�u<S�"�{{`�������?��yW�_�->��44�]q�׳U���òJNc������~��� ���@�#W~�DD����>�����<���v���
�DX���S�1
r[׬��Z�Y��2�"v�+_��w��o��d���7i��z@�g�ɨ|(Ǘ�"��(R�p+��O,KAb(Z���c3c��ƅ�@.�Ҹt�Dv�����A@�����c����,�(P+�'F��#}ء	�<#8NLU˩��n!K.)�|����r���|�:�s���V�{��|���վ���H�R	���6��F�6w��o(k�XVy�U��RS�#���������_�ە|�*[cF��*�p�� m�\���sT8�%ը�z_��3&},@�bH�j��P��	�?V3�,�j\N�%zHsH����w�*3���N>��<W�Y�_�=p��xc �Ŗkȳ`x|@��fk��6Ƣ�!�=3������:����z�Ӕ��K\7"Z`Á=������T ���P���J[�Z<Ye�n����w�����}+�}l�������q���3P�p��3�Nj���V��zP��3����%S�Ҧ�+�m�[S�;��Q��&-��}?�HSV�(��ʋ ��]��5>�߫�˥"MFMB�ZMD��a�u�[l<`,�h�pf� w�>g���	�c�n��:�?X��XT�=��H�&�M�Wy8a�ZU]q���6��������H=�Ժ�eՉu������e ��2����cFm��}#��$ű��(p�zH��d�s+��?t{�+�+q<�'��՗ʏ+���D��dXŜc�d 7{f�	��;���(8`��Dry�8�����+���YG�%�D�ӳ� �i�h4^>�YX"�f����X�!P���X�w���j�U,�@�#��1���X�x �լ7ߴ�k��/w��(��� �ӭE����xXvMO9����P�+�A|@�R����ɰ����}����m7z�Ϲ{��g,�����> g@1�f�E�x��5V-��p�7�6�l��O`W��ڣ���|Z��X�Q >��+7�f��nC������α�q�:�2��3_���cG���4��aH� ���9C�u�I��[���X�Vf�06��5�4UDt�=r�5�+&#�&L]#�oY�жɮ�g�⑁�)�R��l,��a��\X�2�>�6��V{r?J�n" \]���ZN�!����w7�C�k���-�����* %�*E����F-��F��1/_�&�2��:�
p�~k�֛o5�(*�:ϼ��'��ۉ�c����O\Դ �?�-�S�`2����uc��i�T}}��ֹ�y��x- ׁm���/�0��i���d�KcT�3��;�Vü��Q����7o���*����r30�:�o�)@��J��
+7��x�x(}�6�y�CvɃO��!\ےy��nǊJ{�(
nA�7�#�6c�]��ѻ8��i2�_�/=��z�ƳƋ�R�$Ys�)=����jR�����9�[�LΎ( S�F�&�����Pٔ����( 3����4�8��z4M�^�L�?�&iV t�����RO+��V�k��lV�e4����_az���;�i�0+�	Q�b&���T��B�G�|�$R71�gU�'(��"��ҖX�Z}6g�d )�������+�_K���;my
-��o����Ɖ����Q�HQ�o�Az�Y���-��T��$��L�m���k}�~J������� KA>�oO	t�Xe�,���n�j���X�בq�3�
��2Y��b� u��Z����)���k�~�A.V/�_}����������+76�c^@ ��� +(_s{ry ר����X����D� ��9��	�~�֗��_t^�/��,�.u����ڗ�v��e�' �ٍ^���)A�FAC���HQ��V�H��$5���,��2�����3�����e���#��S��^2�8O�Y�:A�&����@���VY��=��䌮e���>��� A���`6S��F=�R�9�w�\��ܔi�Y�	|[ ��[ִ(ii�= ����oux�c&0��V�P=��}.+LH-�J�Ɖߗ�q@��/�a)R�0��-ם)��h��X)��ɓ'���8[�|�|.��5L�BJ��|.�y�O��O�R(f)@%���v�^1"�k�b:OT���@�6�%�ҹ�)*�uz/-��^i�nY�;0>q���y���A\0<0�,#X|���{�r�:�ߴ�>X�C(,�"�Ob9��Q;���Xx�nUs�c��v��G�[�j�U ��۫��pkN6��}ic��D����QT�"k[ܰg���a�o	|��#q��+���#�O����cT"}F�����������1��7ަQ<�w��ޓ�+��܊4� 6�:���x`p�u����l��(������\��c1�;��8ֳ)[s�n�s��Ň���j�
6 ��|Ȭ��X�|K��c'��g�;��� �d�oȌ���}) ��,9�D�	��a��hC���09�9p���+����R�'������Cb�}��v*O�%Y�^֭�Sm�2\�c�����e�!���g�߮���x�)��zO�CFY{de��x���Yp]�vP�����s[n���x�
�����[ <
�X7�%�ė��\���T���Z�3G���QI�BJ&MP�]&���3�-��v�L�gc;�ku��S�_��ۅ�|����R�SX\�$���|��^�����0��F�c�����f�\���6�?�m�	2����q0���q��xb��MĀ벩�g"d��?ɗ��-�N� ��=� ��6�X�����)b̑{��uL���!�[�%h̪�o��ƾ=z>T�,Q��s��A<(�ϲ�xL���g4����u��G��2*�������^y��S��(x�1�gF�|�1������0�paU:�B�õɭ��k�g��?�]3�r�f._��5��}N��q��`9�M�F���T������
 ^�y�9�E���j��s*���l��r��g�@�b,�� �*��{�\��}�;Vx����Y����v����ϗ�?Q�>�v���3icxJ<O��q�����_]m��#S�.���n.���w�౞r�]�r+>�n{�2R��3�^���Qv�>���*�MjM\��@�	�� �ߑ�� =������[n]�r����Zj"�ޗ���H�TQl��{Ṿ;Z&de$��@^��믿�t���y˳/��>Q�~
��&.p��Zrs�SQ�(���[o��h 1�7�H�_�\�4ym��J��U:1hЂ�}��X�<w-�������.�&�<@&��I�,(JX��ܐqA���˞��{(W�B�sʘ��}�.OKh��]����0V並 th�[�]�p�]l��H�m	����*�����S֒u�YK�v���=��m	&V}4��44���� ��|uw�!O�]��/%����+�����Tc΃�q�߾��������TWV�P4�| V]q����A=*֋sjU�4}$#�W.hERJtL���>�n�1���LJG=S�oe�)��VJ]6��J�W�2ξ]��Dy��R�K�=Q�x
w,ߵ�x\&���i��"Z�I���ϛoY��3� Ţ�{P���m����:�΍�7�������}P��H����QCr��) �5}�!i�m�d��;>Q�&	ڦ��_ڱ��H�g˵O��>��C�mQ��>��Na��, ��"�NI3��R�y��hKF�[diL 
뎘����0.�*��Qf���-�w,���������[|��n�?��O�.R'J���1�M�]�߳�rA
���$�E୾��V9����}����3+пT����@;����%�9����Z_���qa A_��6���x����s �b�n�rn�-���ߣ�9Q ;����B}�1�9�24n������Y� %���<�g��� �����n^�u�[��_�m/���#��ï���� ox���y���s]���Ҳ����x�E2B���	,��%s x�3`����g�b#�tU�v�E�
_9Q�x�<���*Py�>����kU��.�K�e�=�r/7� �1,�E�s�H�UC��c|���K� ʖg��a�mbx�Jϔ��V�{?��놳(d��j�\ @ݛt�T��-�q<SXm�r2 �9m5q4���y`�ׁ�u���r�erJK>!��;����E0�_��WO&�Da����R�'�甶a�o��W"XĀԮN����L���O3 ��	�3�z}˷��9�(���&�n��������,��g���'uf��[Ʒ+Tb���e�R��[�*��,�RB$�R�h��6��$v�����ʯ���v�nMd�ňj�7g~�+���ן��g����u/ �ǃ6>Y��b��A��K`�����S�b�W�E!Ζ�!�6Fj��N[��_�*��?���'&��>�f��˕?~�,듢�!��22����.����r�����i��������N�
c��9���UG��S�������y�Ϗx܁1�a��z+y�/*c �&���/npXŹ���h��Y)�����'�s�_���>W�f���2���E�|�O�uJ
�
V�!~��f5����r��!����@B=L�-C�nyF� 0�2���J�(��[�Ρm��ؠ-���\����x�*n	��˗^fb(�:���u0:,��!hI�0��徧����X�P�Qx�����{�0�oF���  a����:�Dۆ\�I�b��v�2��be��

J�3,��A�b� .?c��n��¢wtϿ�}����������g�4z�v��c���w� �WO Wm��>1y"��e:��������Xj1(��>����=�ў�,a��8vχ�����W�-��C��g�u��nE�?D�`����X���9�Z��<�
ǽ~���L���娏P�<g�x���@����-��=��J���>��ʃ�"�q�`�q����"?O�����<�Y�ڀ� k�S�'`�wĝAo���?���>�-����%�����ˌ:��V]�e�r՟��) �ly��
|��{�ne��2��ۥ�Y>��}N�T�sd/;�H��}(]�3�����>*G�ŬN�����ͩ[[�Xm��$�uK�(r�Բ�����h�Dj���J��G�f��s��a�� �KGX�8ӭp=Q�bVP�-��ۥ��{����/�+���4�Y�����OI�3�c!r�&�"�� �J�%�#���h�쪃��,c�*B�6�yZ[�'�Iw�7���[ �Y��������~�D������~wA�g���\��-�>"����/iv(K;���4eo��x������s��cz�vGv��z��� +�[���ǸγYp��̊b����[ 7���ƫ���1���Y�x?��s(lR�r�c��O�m�z���Qذ&bMܲ�b��e�� ���q���ڕOVc2�ƈ�U�z3���w
��t� ���=*Ql� K�b4qۀ�E�s�zd�'��~W<G�O�r�>y��{JH����L���*m򨶚����ݙ���yk0/p�@A�l�ge�ƿ��({z��Gs��qn�Y$#c5�o
rT��J?�:?�l'gf#�D<�@ǁ�3$@P|��x�9�\LŢc�H���s�kz�G���϶h�v� ����f�<^��_|q��"�w1j��Q����?X]�9<����-3�wJ���3���:	��[��ˏ�8X�H��@܅���D���s�I�Nw���>�{��%=�˂�;\�B�~и(�+���ս�*��=���g:�=q�D��'`�-��Vu��x�� #�b�DπX�� nF��ȃ�؟��Z ���\�o�wV퇯�r���t�M���.׼�Y-�H9��8ߜ���D�c�-�W m:��>>�^?o;��ռY*׼�J	[�Y�����x���q�+�N���;ꖍ\z���or�gƛ�f̛ k�R��b[��S�ܧ~�����t����{��O9���k�;�����7Na�f5V
��R�@���� \��8�k�F�&�6B�\�i�"��z�4MXV�X`��8�z/3U��gu���߽�s(��KU�c��#��~��*�i�dDSD#��n�s�5RZg�ȫ�\~����@���3Ex~�0�G�� �j�1��� ���k��?�W
������8pؒ��eI
��_���t_l�2Z��Y�b�ŌwG	r!�!�@��;�����~��l�l-�ڔ]�T�=���t����W�X�3�s/�����?���?���}�Rgw� hx�Ѧr=�g�|��� �̡9 ��IE�q���V|d�~��[{�0��������/�֪BwÉ�k��OE�w-���vI��x&CJVG�c�زt�5��ė��·�U�� �����P�f@YXSK�g�U�}A���m@��� �' ��'�x&�"�K W�p� ��jYt}oQ�ȡ�M!����y_W�x�\Qҟ,m������;��)�p�Ї�Įo�6R&6'Q�v��n?n؋yB���7e��̸�S���2{�y��Q��� 7�n�+xL���.2��n�=�GK���T"z	&�<(�'����4 ����-�(�r��" ��d\��鮻�:�����I�F-./��0���B�F@�o�hO\	��)��D/�Ss%޲��4nl-�@�|N�Z�-�P�zy�C 0@��2�o�>��;�н��O=vd��L�e����@�������O~�,i�Bڦ����5ۂ�FZi�^xa�����g�y����:6��u1��	?L��(����m)�ٵ�ݳ��s\� ts�|�����)?ڌOM�����}>����}�/o�,����Z�k5�P���L�p��������ǋ���a���Y���%�7�q���~�s��A&�}\0�\��8�\����^���bH��������< ��� 7�����Ύ��}��wG��En��d�Ѕg)���{>*���y��LmI�7�'9ٕE��H�<�O{�U8htϽ�G��u�2^���_���#�yO��漀Wf��u�:�锨eG��BM��W0	3�!(�k���K:��3�%Ƣk���\a����cɈ`�_|��~��=�v�{�%���E|`Ժ^ W�?Y�|��}�< �U �-7��x�L\��BY�E(27އXi	��"��g%([Om��b1 ��>0�)�4�//A�������>"�:1���G7����,)!r[P� c_��|�;�g�}�ZpI��ۈ�'Fb9�s���{���q��V`�@F��ʴxGd�񺞕$�
g����:T�gx��{�6ӻk�I����?Y���]��Ƨw���9+�|�#��10&|�ǹ�Aiq�a�n��v�9���ǚ�dF���d �vvB	�*M�c�e�ET��^,J�NP����HeM�r����[��A�l�A�=[`��ɓ���y���i�>'��߽���e||�������SjbC�.���B��k��R�p�Q�9�m��1�e��s�R ��y�(u}p{�;�2&�N%3���-jYZש��+�څ�/] R�����r$i��i����R����9[��i���>�֩��wJ��Si����)Y�X�Â�i�e�o��[H�$,=��$�-n	,�.% ���}ٱ�y�����ђ���"yhe�Ⴛ ����˭<����)�Z�*��V���#e "��zܟ��g���G������u����,��w�|�,�#s:�s\��Y9-�ۻ7��u��Y?�NYI�Uү���%���yJ��~��:6忨�#�]���U���uO��S ,f��W��`������u�P�(�9˜�zdۭ�>���52 ��Y���J#y��j��wϯ\��������E��D	��`��#R��\��ig�����v���/S�=���J�Y�ķ���WÆ���b@l�bdH�5R��F��ޕ���d��.E��|"*�Q��䙙1`�m�&,>���R�[ڴ���G;����ˁ���V��5]��WD`�4�>�ѵ1bS�!�{y͹�x���g?���PѦ�]�����/�)�\� �˖����x<���?������ �5��m��`n�ܱ7�/���k��+,4��o�G7�Cb{|�'����E���3",�w+����x�����%����z�bY�h8�&��[n@�r��}D-P�Ї��po�W>�?��,�bF�� ��mյ�wZ�@f�i	W�r"�g�de �Im�~���#�U����{,b�3F�7�](���=�YR�����pc�'��Vz�c���sY�we
W�̯�o�eW8pr~���Nc?x�=�����5����YEd�-ҏ�|���9��6Bv��$C�r�+棔��r	�Eܟ+<�bBJT�)t�qD>�F\nvvvV��3�F�rF���u)ә�3^�<#�k�����!�Vn�X�� ���M:p����:��[�t�1�A-n�I��T}�o>Q���e1�bPZF�2���~�����:P�훥�/�}J�3F��\��x�1�8��Zv8z�b}�"(��bu�"B�N�L|�&B�y�5�%E�"��CJ,�o9��X��4Vn)�m�:���fX�*8�|�<B�tl���ԋ�|h�cq~N)ǣ6>7��f�W�]�����s���/��� -O��Uy@V�?�~����s�a���u��+`��|�]q����}+k%`L��3|���+-��q�\"�3x��c�6��m=`ϕM��$�����;Z�x�F��P����e.���Α������d.����f� �Rޓ�~�e�C=t��W_=]ڲZr��ZI��]x����cy�J�(�N#���)㟭����ںv�;����������N��e�S��s3r-_�AE��z������w�y����^��Ɂ� p�ɠ�
�-L��"��?��Ҧ�*̡�tq��'^\�d�O��#�Ѯ��W�I)�ߔ�������k>NbnP���e1n���1�5� �xe������f�V�X�����[[EX���ȕE�7��� �������sZsځf��x�:��0i�y������߳��yWTbG,vca��:���d� N���z�3��@�ϊo+� �<���N��9h�_���{��n�1�p�WO�7�՟�22+�]�g
,��>V���udG���(g�G���%� �����7eP����s���ʓ�]/m����1�\�8���?p]y�rBŔ��� �=�����>H� 7��u�Fh�r,�?��c%v�LKC՜o�e�u�4r����_x��%�RyrK�-ן���p�X��4�>������� W�}����eG�'��>c���Z$� R�)n_�Pψ@Z��.@�{^LƑ<#)8��\[ ��Su?_���Z	�c�p�8.�nC{yo�%�8|�q�И%j�O��j�+�×w'�t�(ޭy:«6- �;��R�[�l�r�#P�����$rw�4��
{Ϲ@�'T�l��c��� �UD�9I=��V�4�B��ݙ��\�d �(��ǰ�A˴�[ǉ� 0w�A�����-`��0�P�i�/Y0JYr�;��/}�P������k���O��vW^o2(��!�H�R��8c{�����}�Y�I���(�zee|l����+���5���
���Q����S)֩�c���<��,	qS��U��a"a����>��o�Znϖ2�<��$�+ߨ������)��˗�o��*����!�&@��������~�,�c����2,�U��X]0��,�-()� �n�����!���c�Q�ֲ0�$��ro,��7�����̸w\1���ݻ����[��7`�s�6�p��#�p�4�G�u�~n|~�W�xq�r���g�[o����~��"�c�#�O(O�3W�D�n#�q���?��1R |>�%�z� �d۠n"�;�sd.S \��9Ȝ�*-}�Չ�`�8`��x6�G}uL|Ne�|��u���c}�Tx�S�}����yT�_�[�`qv|����qw�RЙ+]̑�A����ou��z��!+��e�Q��9��>�*�Q�G�.sȗ�Z��_vG-(�kU�O�����%B�_�V���n|$)W�\L��;�yn���AI��o�3�<s�0�SX:�r(�����7'.�X1y���!J�B.��Zkj��w��|	՟��%�C�����ں���v����O �C���n�=�����V�L!�\�uB��v��w��к�{�Y���;���Gfc�bU#�'Qkn��[2���p��AYY�Z�����@5+o���e�+O�8_�u_X'� ������ )@.�|ɀO,��v�n�EQ%�E�q	 ��C0s�Kns��J+����h0�<M$`޳��nz�ڋLj|p��~��Ǻ�^|vn�P���	���o���EF|뮻�zT�
r��*�� �c�3��(}^��j)ܣح���Za�#{,D�3��z�Z|�c#N��դ)Kq�2KDV攥9;�i�<X�%Z�	��a�P��<e���n�R�ۧ�4�>�� ����-�#���Yq%hHy�ߞa\'��˕���������,Sz��`ׅ���U�����*x�bEB��X���E�&I�U!{y��V�k�Q�.�������S:飱��H����j|�i3�k3>�wzȩ�۔��x����?�aOY�c�E@�|�~��9���5!�D�ZCR&�wna�|��k�?}�����к?��Z�"�y��B��J�ȓ��[ @�,x(��揧��cu�Y����[��[l�͊���1���]�j�e��r����&B�"����gͮp�=�<J����٠>�j+��Ā���k4��u+�7- ;ba�Do��~���)wA��p��Q޴Q��z���&��y���ұฏ�U�r1l-s��S���\����ɓ5cB����qw��&)��/F�XX�a�@�D�%�%@�UM�n�]�|dA��p���JY�DX��"���h�!=��1�M3.�z��ˮ.��0/�\d��\���Xi��~���'n���p�p�̓( v�#mY$�x��X��Y�i��	Ef�AE"�l��*�)�lNݛ	��5��rc�oO� ���i�i��V�{�G�#��W�8H�X@�-�#��>� ⁛��r���\0��DsT)��ĥ��vaQT*Uo��3�#���D
0�g���O�ډL2�|�#9[��dj��gig��}�{���ޚ]Am/�Ʀ����¥�>P����=���Q6�7�s�=\�cu�Z;�C{�}�\��A�wky.ZG8��F\��ۍ�L<���	�m��e���O7q��'���;R�����Ә	~��Q ����.L�-�N%��[DW�����e��9
��t|W0㳅p�s%pt�����_ �`$@�-���'��ƛo��,���=v���f�?�'��vCA㝱iyY�檷��n��3m���9���/�R�
1�݊�����m��-��}��w�4�.�{�Ř�@-��Bc^F �?�9\r�c��g�(\s�����uD+	�,�������Mݭ�)��*S�[��RT� �d,����Y��_�ӓG���Wj"/���	@�5�>Q��)Ğ�ErqH���_����^z��+m_S�i"�\�~R�L>v�Α+Z�b\����\����r�)Ǳ^�7��+3^۲��g��}  �(��uwD0�1(��,��ݭ I09�,�ʡ_Ѫ��vs*���O�?�Ŋ�b���`��W� x<(
�������jY=qC���B�X��,��1pk��CYX|�VT���_�}��cB�
V0�O��]^�kG�[!�N�h��-���3݄���'@Z�El]�}�����������߿�wؖ�5���v�y_�k��P7PYZ�4f4v�e���%���w.cnj�ɝA�H����)��" s�8���'�RD?y����8����<�\�c��J	�b��0�W�wg�����-�1��-ƴ)�T[*��p��=����~�����{�U�ޣ򫕒E܅�U7��1�����?ٗ2����(��+��"�����|����Qhd���*e��ؐSB#+�%o�2tX�����Xn���̵,�$��]ʶIEH���/y��˷
�x�eC��"�"=���]���-�/=B\�/ˍ�>~|!�-�e��DH~{^NzѶ�:'��pv�/Ϩ��u���¥�{>���\	�#�C�<_���&�s߲\�􃃿Q�Y�/���%����% �@����u�����6ȗ��@�~�9�����g����}F=ؒ~!��K>i?�ni�p �����HveYYk�4�ӗ��c��GK0���E��y_��,�9U_O%a�����h�b�% o� ��n��m��?\������2^O	䊟���#��C��K�ƭ��A��uS��(λֳ⸊��5{xr�;Yp{ �e�x/�6�OY0 �f"��N��x5x�w�O׉9j_�Cp�]��/�p�0��d�<Fz���-3������/�S%����s+Bi�?�'t@�2<��`���D�c�a���o�uQP}/^��� Tꎒ�{��G�O�Q����#q[�gF=�t������f���#�L��c	r��
��7ʜ�VY#���O��I"��>�˴T�U��*�ya��M] m>?P�p��6e	W2�W>"��L�����3?qs�q�����?��o��������)Ο ��#��9�����ɫ���#��С�vK��>����S��O�s�>���0:(�{TR|��y�7����+�3���w�02�R���F9PKc���#:gY�K��ۃ�����v;�v�1,�g��Ч>��s�?��SJ&�Cq�[�-
�OO����о>�Z� y��iu-K�����e��ɣ���"������"$=�ET����R�~+�e{�1wI � dpi@�˚E�`�-j�	�����z�wMF�Ǯ����A���+�@?L��B��p) Öˀ����>u�����z֙�#K��oȟ�~�ٳqe��VB��)������X\�f�Y ˿�E�.+(���՛�đ`���
A��"u��zO�S�<�(�_WudǾt ��Pbn��kƉ(�r�0�d;1�+מ>���.�6}����oOi��E�
|��7���j>�_�/D�y<��zXgd>�΍<w�|���o,/����u+7���A��X�r���5A�+�aڗ��55)��wk0?U���e���o���"X/L���'т��Р># ��!,w"���+�0�*E}4ļ�(�Y��rk� ?}#��A����n�������%qO�Ʋ�o^��������>�X��֤h�iˊ+�H���W���`�z߸B���K�l����D��22�DXh�'���j7	C}K (��`��O�0ĕ�m��Qp�E>�[`�����!J�
�T���d�JCb�])�z
���@���[sAQ�n���K�Pn ��{���8���T�"�h��`߼Z���%5��ʭ�q�
�+�����-�=y�s}�t�����E+���e�
���(�"~�|���1��+R��jK�뮊E��3d������ �h���z�g�*p�)���;�_�lg��Y _��K[ÖﳅQZo����s�=U�O�M�a���K_�� ����V9��ǖ�b� �q "�V�$P�Ҁ]��N7�E벧9�o	ErsQ�2��!�&�[����e�7����*[@M��1?�1xv�[��>��\d���5��7�QXIˆ��R��ރ��U�H�h @�W�}�o�����Gʀ�}Z�TJ���7��g�D1�_[m5�m�%����r���s�4|XL1`E��0����bU�1˸�ʋ2&,���6�� ���^��BXsS?���w,qd]Q��n���5�y��2l�ndHa�Kʔ�#��]xO_i����|�e }���R�ӧ��x��;
�!�̸/:2CcH�B���1c"f���xNQ�j�Bs(��=��w]��=p�+h��զ̌��@י62F��ɟL1@�RgI�����x��C��������[gX>�	�"5��ˇ �aͲfM�}aw�0�-u?�.����E
 �?�]�.^��pXhX�%��-��@�"���EȻo�/��"�z�;������G���@s����9/�w�5D�I�.`��}���kc�;�-��+�Cݕ	�A��G.}j�bM�V}(k���?�]RH�?\e�X����(e�s���~nqԴ%9�[��+5�]�-�NcF�لE�(�H�}}�c�1�ઞ$�g���v��.�*{o���.� K���9���1�2{�t� �.�+��Հ_V���%�Ot�B1� ��9[�?4� ���g��?%��2-���?.sE㘻+�9���#���
P�?s,ȣ����ӄM=�z�M��pMO ��KЗ� 9�~����$��
�9��^%�RQR�K��si�S�a��-�,!�Ef}��%c�
�֔����LX��#2l V���@�ǖ[fDѥ�e^�#!��'�f}XNE`�9���0c0�\+ ĺW�[s� x��9O)�>'3�m�w�QcA���;;;��|�3�~�ӟ����OV ���eɎ�����wt��X/����C���E�N���^z�ŋ/��x�w����
�mXd��@n\͈ Zu�P���n^� ��T26V+(��2��nýD���-Z�Q�������A>[��; �1� 3/��ee�R"9��g������B �Q|���(�(��#��WRh3|��5�y����~���C������k��A2�[�&���1�q��������)�^���@sm�Zx3���P��Eқhך���Ր�~hC�-���v�ų�0G+�5���3>��!s�JT ʹ�~��g���	�YʹN�ΰ�L9��'���A��e%� u?Uϰ���~R�NE2��P�3�^a%c�V�e	T]�%$g3B_a�q�(b)��0�q,Ѫ�z�?�K��`ط�͜ZKRmM��R[
,�E��K_�����|�Xr��w��b�K�[m<ȃ� Oj3��'H��}��*̓�-x��T8�wP����.���|SĸCA� Q,����7�у�P�{`��P(h;��R&p��Uω����u\sY�ꫯV�D�鸔%Ys֒�3��"Oǻl�ܦm�G�e�D}��z��/���*�Vi_{�J_���D�dw9���{k|�-�}~���m�E��ֳ�hγ�sC-;��Da�^����� x���0�:/f�/�gb.� |bqHW�
H8�ҷ�3(�V`�  �#䵄���~{X�4p�P4����zN`Jy3�tD+m)_VB_�����C@�[�ȳ9���4I�J)#hǗm�����D�㏌�PY s�m,B�깔ᩤ<`3Z2e�n�k�x`�m�z��g?��
tUg,��~ppQG�ڮ��q|E ra�� Q�8�c~�OTˢ\d9���E.�"�e��.Sp��;�O�����󻛏�tV�%�d�W�SV�؅��z0�y��(%�q�?+�>�p@�T�`�kL��hL�B�3��(e��jg��oY�
-� R�5t����|J��C�*T�����kQ��s?�P��oط��ʊ:e^ר��]�=����C-�{-h��3�d�E��	S�7��`$������5g�?�8��J���揕���P"_j�eT,�N������b�t���J@D�;�S�D>� ��D���W��ݚ�s� �o�}�}�r�˲8a��>�P�|	M�5@�3s�]hڏ2P�t@ĵ�z�ށ���UjS�-+k�l�%�jiY� _O��G�� _|<���,�����З�Q"�?���'?Y������Ui��]��ߺ�Ϩ	+�Ί��("mk�~��ƣƪ��ͷ�"���O�O�.q���1`���%�-��09�&E���c��j~�}5�pq8'�
�+������7�9��汿��LY��2'Zo�"�y�g���)�u�q�.n��g�pE��E=~��1F���^@��9�Pׂ+ꙧ[�=(j-Y� �xOv�Ȼ<�V>0�ڰ�� �
 F\�:Sۡ�|�I��J�--ea�#�,���M���&�B��Q%�f��qQ}[�z{�����nU���/�2P��<;˾�,�;����ݱI������B��,��*Ã(T?�0`A���r��UK�,���1�~8F,�|�׹��s���zׯ|�+��oY�UO\;�z�ÕG�ӏ��M��q�S�1��́��-����G��oq��L�Se������������j�L��Ob�bl�j�Ɛ���Mk��~���A{�<�?q~q��W>�>ta��o�u��x6\V&|<yz.WR�3�;����[o���xCqa5E�Fs�{\2�H��λ��ܷㅶ����1�V�p�x�������4/}���5 �ڪ�4w5O��f��l��_=săG3��6)��l�fW �ѽk[uu�����3��ղ⎀����Ȉ2Sy�YXoczO�"&E>G��k`r���{���=�Q:5/�r����TA"��x*,�A	�����ƈ��Zԋ�������v���]?m����r��c�x.LR�!���\H��9�(@�G��<�iW���V,w�6"p�7n<�@�0d.轱�BѢ��ޓY9p�P}���}�}�-���/.����fJ�b}i��e�x5N.����� )��ɍ�Xz�����K��[��6��Q`W~��O�ux6�ď�е ���F��O ��P4�0(ϳl��"���j>e+�:�9����6�#"<��x�sl\����," I�,c�7���:F�[6n��-�S�xAx��Ail��<���l,˱�r�k�),��5���gʜ��hݾ���惏��/��v5h�K-�pƧZ�[�{҂۪к�גZ�[�����"���p_M��0�8(�~iyQ["�'\;�R���?FV\	@w5 (��`"�H��8���	���������^z�\)Q��b���Il��H���m@@X�=�w,�Mϑ��R,TYn�$�Tw��@]tK6>� �
0�[�'#H����X�� ��{����}��k0��$h�X��w���>�P�����u x�s=�H����Ʋ�Q[�s�f����8����*O�N�\cG����
�*ݖ�):h�X(=l���݂j����Gv�,�R�zg��U�Z���d��9h��V}	��2�ݯ�y��c-��d�@���c����}i}U@cJm��e�FJ��A�@L��2��	h-骓d�/�Pen]�7��2�[K{�cf�<(ږD��\�-{8.Rׂ�Yj�+`v�z�����ei�y`	�
˕w�gNЮ1��'�@:L�}�0����A���'r`�2C�K�D��rB~[\EPfV}mu�@ ���XM�A��ڢ��~ �l�O�a�6"�E��O����\,`*�4@Ńn��f����j���R��z*2��A%m��E����9U=nl��կV�( P�5�|��<���%�+�B���>���" �V���>1���Z��~+�URaa������==�����&��r����rU8�\KPX � \�����$ԱP����.�҄	��p|oɖ ;��ʒ_+Jc�� ;�vW��pݧگ�:�5� ׳	�������M7��\�b�?�m�WJ3�%����+���x�pK�kGeܟ +`  ��*�q�1bD���]!{��rFW�z.T�x8�E�ɗ��� w�cz�	�t͎Rn�3!��5�4I^�:S��!s���)�dD��@����u�P��դ����V �-�Ԉ�i<�X��(�V���U��9 ����`�c	ӗsEDaG\P.��ֻ������N�i\,�+Ѷ��&W0@�` �DQ���R�!��H��C����7�<�H��T�kѷ�Z��@�Q�T�.���/~�x��j�RK�&w�p%F���KÊ��Q�V@G`Udl*�"Vw�2wO����=z�J�r�������98�s�'��VNw��R��?���j\I�P��?P�PR�rߝ1��}����8��F��r=�2�j����Vo�S�/���?\7�����,*��*����/ަ�v?�t��C�f�����؇?��u� <��@� �桰d���nJ��6S8Gʙ¤[̓�^��������ݺ��!K�h�T.�z޾��tPT�Q�W-iٵں%ɭ��Ċ�W�e&��ri���C]�n Eߞ���XQY*���|'& Y����O�<����Y���NQ��*HN��]x������W�e7(�஖�/��3�?_�-[M�q�T���(7�@���|o����M7�t��2m�K����U�x�Z��d���n� e��	��Z���z��HcDm��U�Զ���}��Mm���%���+J�����p���P����ݗ��-}A?gA��d���vv�/��-��&�u\ A��jS,�:Ʋ�[�Dp���z�ۿ�uW)!ݘ�GN��TsM}ע�^|���4FȦBz.ۺ��2��9/�ő��pK��'Y=J���5����MA��"���=`��|��,��P����mv����`�o�ެ2��G��զ�Oի����O�� \\�)D1#��\�D[&����|HN�?ϔ��X�S��;G��L��p���,�?�L���zW��2���S����� ���>��L� |0�=�G"�E�$���X�<���K�$����s�s�;�2w|~R稤F�Yx��V�d%�߭������_E�c�M5D�?�я��P����X�e�ָ�`�Y��"Le-��[m��S���?�uV�O}�S��__e��������l\Z���P��T�����[w31V�C�8?��)(��9 =�{����a��j���f<����TA��7��?��č���n8� M������L]�J���\��\x���>��~=�����"x
�_=Znݘ�%����(�^��mZp]Xd��z �N��g���Wq�9zdWc�z��j!��c�)��c�������j���|��z�7�
��Z.]Z.ɚ!�J�&�%9��d��۵�(8�LX\c"�8����>��g�R6� W�+Y�
V�rWװ#�߭��qY%H�OnS�C��5�g�l�e��+"��	茖��e��� ��Vn � T������?h�+�@�s�=�����_��e������X���R���Y���q��*C� �|R|��l�y�U�.H�5W+���E�ľ���>��z�� �ƪ����R��X�`LyT8
�K���s������٨��F���7k��*϶���[� ~�1�H �l:��
�3�E|'o|�"�|�c*�q6���� ���2I6	0�����ת�v����9TUw� �������kxֽ�gXF���ߙ(?ЩgM}�ߥ�2��ۺ��ǃ�	Fr�*�o]ݕxڛ��P�������El��ϑ�2�6�	��\�؟��#'��Ezd�2U�utN��,���� �%��7�Q2U�����C���`�4���3�ף�Q>t�M��$(9���p��LR2*2.iF�:0e�' XL��>��_u���_��w��_�M�D������.�A�����.�2{�f1���4`��+��@'������\�&����	�Aq)��,P�ũ���aTɔ�[��?Ѐif�y���!)<��s,°Ҿ�$�v �5X��{�{�w�g���f�)�. P�
,.̸m������_�z�?/�*[��rM3��w�왑=���(��H����~�������Z����������& �	�<�����e����� 
x>K��s���cT�2��س�f����x�̋�_e��'m}qmL���bH���� �����v��}� v���h��������G��U�~B��*K���:��G��E�;w�K`�yS���ɑ�E���~J����w��x�7%�P�2rמyZ����	���%)��*����ɪ�s�����C��䆘/։�	K����,P��_P.�5�B�ld�ؿ�ͷ�����5�;�ʹ�`ƀ&�a����A׏v�ٽ��9�^�ؖ���7f��k2�(���KҞ>y@����I��>� ����7�1��7�9{����5՗)�pz��f�֎��@�>�\V֔N��w�PL?���B ��2i�?��W�����9_���;���7�������� 
n++��q�A`�Λ;-0�׿�[\�rc��u]�x_�_�3ȸg_���"ɾ���r�J�c],2�YfW���H�N�뼖�i�x6_��:� n���8Y's]G�ن`92�ݓC�<����=�l?ɬ
H��B4�S��"9���b���{.�x�ߦ@���O��n*�w�j���4N��<��*<#�38A�8�Lm��I�C�\~zkdl+�4�Z�Z3 ��: 0�%���;'w���yC�M�h��n�gv�:fzc���~_���Z��<�@����i9'�lڥˍQ"���{'�W��jZ�*��0.Hd8݌�,�Ņ�m<nu�֛����X���R Ӛ����/|�m�kJ����,y���k�s7�.�{? v�rPV�Ϣ����w��n����a�	\1t���eY�e�IOO��N?�ܪ<�q����>���ZO�,&�-�-mc���{�j�u#c���k�k]�r��u�f���8�tZ0o�5�c�6���w��֥���������nj>_݊8tˆ`9!2��^�x�����\�Жh�~��O���)]���֘p�ByUY���&�Yr�^ioܦª�x��f9��k �FN���5����O�����/& �f��-��w�ol ���}89'�uӏUs�����:qU�@Z2Z����BiꩁbN����۷�����d���u�~�6Ҟ���n�/ ��gh��e�-M|���	���g2pGP�ؔ�ȓA��m�Np�� ���>���N�1�I��=6mX�ﭜ;������m�g7w�#���2� ��Ղ�����_V���.LG� ���L6=���]��G�3g�|�^�q�F8�s՝֕�!��7��3�wH
 ��:K��{��m���F�u��s�u�BD��E=3�M���ۏ$h�~��V�|/��g�\>�x���󨃸��h�. w���#C�9����Ϲc@��t�{��aAt2�ˮ�0��I�EH���ދ�K�&��#��e�HF�g����(����|)��m�����"6������fJ0�qre"t��Q�9�91��%�ϐLh�b�������_��Pv��3��J��"�\5�
P,w��ɴf��&�K�к��1ѽ�|�KM��v�mt�ȅ+� Pp����={��g�f K�"�� p|��� �-�M��|��rq,��g�^<���g �ܛz�G���b귗�4����`~]���]DU�`�o�wO�6i�sk���b���ֽ�So�s��!�1W�k\�ӌ�K����;���w�����fIp�A��/9F��� 3y�{�"Y]R��9����5\�������ud#'G2��}I�pl?uп�OY*��Iӵ�w�hf���d]ڻ�s�3���B��-gN�Dl��H5�	�'H�̦`No���|��k{f�>�n��1���儛~桕!J��
�����W��y2�����ahjv�E��s�+��`��MBzMʂ�dis\��L��瞔�O���]���z�0R^�Y�=(e�@��wXO�S?�iqG�au�1���z�+]?��e35]��8���L�&X��h5sE�ǵ_�/���<?;������t_��z\�w4�_�7�WKA�CǙ>�։�8��9_����4I84���vv ��I<��>�����;�8��k}�-�YM�ۺ깻9.�����~i�~z����gaz�|ם�D���欓Nf��I��WB��76$�ձbu������;ARIM�"ƷN�UI'`Ⱥi��Ԟ���?��/�N,W�9Y���`���V��	�)��9'27��}!���q��/��į�4�R�K2L��L���fH��TspN�F�S.ӚYf&i��v�m������2=���i�j���.��e�����3�i��d�yV|]a9�uS}n�Η�]��̆���e�t������;�	Z g}���e7�p�&F��EҷT��q}��d�������-[��� $�ʐ�Rן꟪�E��T�<<��{���dZ�,k�V�G���� Q�����"�:e�A�Ȁ7���-*�N}ng�q��;��ۗ��p�i;n�ܬ��=�2���|��ly���ҙ�-׻_��P[	i�|�n4 ^FO+S~Ty~��+]������4�wcJ���{�dl��2T��|�=��o��0� lLJF>s�����?�>�LP���[Ƙ�
�A(�a'�%��E���˜>� �wU��9k�L}~5&Z������6��wd������[�<n���v���<�	����Rv��E�uXa3"�iO��y1?�*����6x�&����{��m����A�|��������6x����-�?5�inB�]�o{J�|PM��~�����L}��~��3A�V����S���.��d˕�⓯��|�7���¦S��m�'َ�%wED2;/~����fΣ�d�̩��(d��Aо�)�����`C��r�ӕ��,ӕ�B�H��]�*#��Y�ګ��h��H��S½g�=��
V���h��H�\ٚ������O�#��m}���d؜�C``��� B�hb��`���*�Ҽ�o���fo�3]Pn�,g����3?+@Tӷ0��=��&xC�_L�-��_ie7͖[�6 Ͷ�;��.�9����)xp�ϝ�z�ނS&\0A� T]*,S���Y �䛥��ҧ��C�C�^.Y�\��<\�k�d�s[o��g�I����SF�A|~ao	:��
���3�JЬ�	 ��9t��wwj�?�PK`(e{��HN���b���l���)oe�� 9�G.�ږ`S��T~�+��d\���ɻ;��.� ���3ǲ�Bȱ�x����鏬�mn����$m���FN�0�����n����u�ힻ��P�"}�s%:b���n�U��녁0�Y�8���w'E���o���z�Ն�UP1&����Vl��ɔ0|�駟~rh�m����}Ĩd}E5EW2�����Ps0슌�!쯿eM&E΅E�<+�W�w*�d� s ^��}d|�n���g?���,�"�k���|G�{�Fb�v�3�b���A��/���y��z溽@0�7���pA�����d"���'�t`N2�K�%+��s�O�n�?u��+u�e�Q���X�\Mӈ`����|�3�w�	����A+5x�r��蛼x.V�i��z��@eT��M ��7�A�pi�������T'#���ۗZ�e��|W�q�:�k��d�+@�1��(7}���nu�������k�K��\��;mg���Fv�:�7 �d	�i����C�l�z�m�3H5��,Ϋ`�U-�U��ճ�T<y#��;�W���*�����fj�D�9�k����˗l�1�<���c�(�&!R2A�6������]��l܎�	QVվ#�%k�y�\$wE���~������	�4`fu���ߵ�2 �k �f>Y ��L����4]#�����!w/������L0",�Jy3����o�t�h��r0��d�,��ܯ�#@^2�/�0�0g*�� ��A����Z���ˈ&m�+ಏ$����Un~v"J�~m;Y��8Q�>�Ԧ8�rӓ$�Vi��z���G�E(��U6*3�$˖��6����>��\�Ѿ�E&�J�茁�[�i���a�sahy[Yg���6��ɕ��N'!Vl�8�;�"���q�L�E$Í�w��h�)p٣�W�(�"�lM�8�����)M�9Y�l_J����/�N�6m|���� W�M�	��q����so�r��I_��^A�b�,"fo��Y@�;�0�2 M�ݳ�A+%}����9�2���(���J�bS)�}�m�� �yv�B��X@-�fq ���	��i���_Ҋ�^��mˬ��,:  �}?��O��d�&p���ț'׾�"K��'�[Ĕڿ�ݞ�.���,}���덾��e/��t���7O���W7�ӍA����gF
��eԥ�NKɲ��W��� �����6q+���Թ���9�Rqzk,�{jn�L����E�Fn�d�o.������^4XA�j���"��~�����2��ߧ&ͪ��!�:����������6rr�����#[~�NTR�՟�~"���Ü\e����{�㔙��WSd&�O�&A�&J�4���{ �}��{c:����V��)}?V#D�?�:��M��1��YP1���f�S�>����,R��AY3�E��$J�A�' Rwk�u r�(a],�����֯|�+- ��8���cj !������q�:��c����7���m�0.�)����x�-`d%e���ey��f��%ŅUfQH�m�ީ���L��8h�����^yɬ*���E�m���,���,,bd�e�i�$;��b]Y>]z�Fާ�.�Snr���d9��'	1����x)׳PU��S���q��UɎ?:�;XS����8.���Ɲ����H6c`v�%�GZ;�� �]������L2}�r�	�`���\�3�
�������f��,XN3<�2&�$���8���|��K ��<E�E���QX'p���!��`(��y}��L)L��E��&]ٽ82��9���%�;U���Yy�&j����R��s�r�� �����N r���L���Ƕ�o�n���[]�V�=�6���z�<�Q_WY��H����6����$�銓���Âj�"�Y����m�e]�wZ.tYqa�΅�h�*��l-B.�7,Wش.������d�FN�8�����k�+��t�1�y���a�H��U����I��g������[��S^f��e�D����h�U1	�7��'[�ٲ��}�[�TvJ�C;�d�>m�d�\^c������o�I'���K��`5}_`AT~9�e�.�839�V�`�����P�4��3G��>���w<��w^+M��X��o~��E��'��cn�S��'�{����,l�Sn���e���T�de3PL�K�I��c�I��K�.��Q7P9.|*��uT'B���pX�Q֫�*˙.<�.�/�s��6�:3n�<�#�5�ϺG�nb��N��fJ�#�q�/i?6Zq\�y����������e��c5�;�\�.���������<�l{m?$}��nU������H�٫b�k-��������r\T������Ɯ���ݩFs2�<�5������	p7,�����EL��dT�1���v���˗.��ΘP[~�;���'�"�xZ6����+�^{��y�>�D���g&w��pm�C�e��I}t���OD>�݌�K���tG�,jF	[�#&���Q�F�60����������Џ�-~ʈ��3�Z�,f\�Ĥ?e.�mk@���� �߸֕�_�7g� �+���"	��i���H]�d���� �^�U���j1�������ڑߩo
�]��@PF4w$䜴�hm�{����-�����0-$	jҪ �����)����Y"��☿�D�F���]v�/���V���ۓ)����2kY�[������]pW������e]Z>�Y��5i&����i�U�j��{�P9��d�׿���F��S��vOօvTF{#NV�2�a��!m;�����k0�1����t_|6m����.��A �C�35e�ܟ{��f�6��=7�:�5�Ǡ�V�K���=O��2J�sN�W-%�H�4A�cV���� D]��Է�:�S��M7'�=פ�f����wַ��,f�0���2�Y�vW�R��:�d���^Rd�����������m�
�����L#�=!ʹy=����;�e9e9}v]�݌�	��S�f�H�WS�o��G��/��8�'��zM˞�����^nu��e���E��sޱޭG-*5�n#7V��g��ŋ���	�k�㣺nM-�{���X���E�V���2���wg����B�KVy|m���4��%;�
W�->��L�o��FN��xah�m�I��u�V�w')���Nl�$ ,�'�=M���x#Whn5*�")����,x�4X�K-#˶����0����
���v��8�=�ů�:o����ͷ�wmԺ��^��2�܊yvU���$��AMm��ݿ��e�S�[��-�jo�J6�D</��֟��JnG�[E�˅�u���81����E����#�)ђ��ֱ�Uˇ`����Kf=YG%�#�Ӛi�E��x�d���'����O2�2�b�M��ʬ���o]Rx.�Qw�a^mA��]�!�`�t1I�X����z\.���va���#C{]�㘃��R�:��z�G�N��S�t���{�����z�/�U_F������r�*�F�:�*a�r-Z�Կ�a���4%U'q}�c�i|#'G�qEf#�"�E�-�>�O�I��tZL2���5sA�9wS�U킈W�����I��*�9��6A���� )�S��2Y�j3=p��ɞ=sv�E�"xJw��o֫L��i��#�6J�:,M������O-O)ՠ�e}'�s�u~��YE�԰PfI�J�\o2�a��֭�*�/s�U�&�f{��-�2l��.��v#��1�M�O��7L�O� 4���ֻ�� m�ж��.�����d�������?�{Zs��<�}���2��+��x��6�.�2�8�~35&��Vp;l{�Fr^�Z��nU|��f�aqWm�U�p�~�������T�?ϛ���?A�De�r�&H�PJ2� E��V�vg���w.}<�LA&��u7,��3��PK��T��V�[��gX�X� 8GN��r�_� �
�3>��>-�u�Ns2O�Nf�2���a��X?5�dx?Ң�@�傧���������'
�/{�n�{jN7�	�L�Ǣ����6�)�Se�3�ªnS9O\U���+˝PS��b{Xf�T��g�	2`�'���J���2��\�\������Ksq(-k�}s#����q�e�P����u�,��8ݘ|�l�l'��������� %[��� �+��J]���l�*S��0 w�4a7��]w�x����+c���S!�U��W���9p0(��������m䆋;V��d����zj��8�5ȭ��:�95�~���a�����}�Y���w25'n�ko��w���,g�BI`ᄝ`S���Y��i,7,�i��Qμ8��_a��m�KV��������6V�w����ѝH�WD��2�>������m�b7}�\�d���.�o��~��	�22���4�/�=s�
���,g�7~��%Itx����zs���"�L��k6�Z2��æ��`.��Ό	� ʦ2��^g �,H�8�-�-k�.撖i��n:7{�]�m
}��9]��X���|�=�@���.;.$��2y�#��se�0���������?'@�~��5��C���3]�2G��U�BU'�+�b3u̲���S�im�{d�]��oS���"�������d�d��L���h.?m�	�A��pǨxL�s����;M{X��A7�|Ӹ���,	|��db!�E��ć2KF��5���U�E.@���Ҫ��%8��B2�IS��"��9yfpJ�7�r�C3-�~)}F3�;�ޓY��]r!���)ˬJ=@�
Һ�Iv��n L���G=S�>[�ՠ�l>g��d�,�1/7�=� ��wW�X�����am'߈~��ek;����,��f�|��~����s��
DG����&y$�k�p�F���}���0�Z"�,�l{�Ն��ҙ�a�&����kS���� @M�lA�u��|V^�%�F���Ⱦ�Q�Hna������f�9��K/m��,�Nz�U��}0u����=,�
ȭR��y�(�{=�h�wH>�B���bW�6���#�	��_~y��?����}yp�
��j��XLv-W�֙12�I�> x����޴���뛬�1Igޚ]�|i���kF��W#S{e0
n��3��"S�Q�\#+�k��s����!ml���ɵ��@+i�3�� �(ҳ��Z����n��+@����~��$7z�b�P�˴R�O������;&'��}�[�͵���&��MN�ǳ�~�o�z�W�.�m�����tQ�����#���	ꓥtqŘ�G����ϝ��-�t����3>��6}�MZ�ׅm�KBGf��^n��RL�@�{]|�֧1�'%}ks�� w�6��	��.��ʹ��8��َ�FI�e��8�g���暫�ܩy��=�}h�{X�~9�{��E,E��L��T�~v�����i��:2(�/oۚtӵd�;�R� ��z���I㭷�`����0�\9u���?���$jP�n`mB�!�,#����U� �,.�������ݽgh�@��e�)}��9ٺa��������+����!�/+*h���_�*�~KvXW� �
@�, �|�=���-w��kz]��8 8�n����H���7#��A�Hr���������Yn'�?��kfPȅ}��ʐ�"����>��U��e���z���b��[��w���#�����x>څ�u���������[�R��gƛ�$����wq�B!�d���U$�sVu֕�6?�~��#�q�l��2��+�bVO��m���w�3�~�zH�7z ��S�Q��
��}ze���ݡ�:rX���S�WA�^�w�2��󲒍����3�C� k���o�u����+�G��3'i�����'�؂��xs����Mdw8/'I@��)����Pn2�*1�d�L]Żn�����s�+����# �w����X���2�#��;�y�t����	���:�C�m��D��b�.�@�����]P�,�R���5\8�^�"�n�I�T����ԍA���oڜ����{��^h���L�[���}��g��w_+�ui9��M`�s��ҷ��:6����d������d��Z���5P,�-[5�g;%��������To.$T�EX^CP`�:��:���nk�y]W���a
 ��@Y\��D{ ����i�d��g�=d�eo����sN�-������?��/��楅�]�X�f�9�,�G=�S	>�{�3���O=�^�BS�/#g��#�(,��]Uzٻ�"�u꺋��IU���JI�eK;��S��Йw7~�7\�6�0Ll�-Zz�n���Q���{��G��6���^�������n��}��1����̝�i�=QZ�)J��2��,,�4e�E��۞k�O���� ~�O�\��c� ��s���&�Gd�)?���F7��+v��h����NF[ХiN{5�/2���I��1G;�n2�d@8��h7.�[{% L_\�?�����������1�ס]3�
��V����'g����=�HMe�	� ϸPp�\������~��{�nx	��&�Z�������e��;M6779�'��,��"E���i��/ژ�̧�{Hn�c��l&��@�K��X��O�Ü�.|�o.ެ��?��t|��o�W]{<�2;�0�da>���� � t�z�~���c�E��S |����2���.�S�Y���@����Q_�{���6U�
��RI���V'�@�fi�t[R�"2q�q�-�n�����x��1�8�■�?g 
�j[PW$��9�\YWYC�T'BY�h}�����-�1b[ �ٟ�������fϭ���
8�����X�'5�������� '�\0N���p-2G��f&
7�p���R1x�M��?�<����f�����u��\�'��l�A�*)�	ׁ����>��='�)�L���[�-���E~$��_�Uc�i�՟�ECnna��2i�S&F�V/�a��`UA^�>{2��������	��9F�H7���.d�_�F��쟸%�j�S�>��eJ$�vIFZw�����y�W�S�������o����п/��+ÂmC�� ��~p��?���k=��dv�H]u9
^�bv3�@�,������{��	p������=�b��z���/�u�*�(+p#$]��QU2���������(� �c���/_��v�mmRk}o ����
��wF����љ�2��d&8�|�ߦ=B�h��U}�������%3�ɷ��D�R0�]k�l���U����i��o�	��$j@���$�ʲ
|��9�TV�c�	�,xib�}(��C</@n�60wU ,�r��9�����X\ �0� \�����3��}��o>���3G��/��y � [� �0�=�Pc���@9sf�[@n��[��~�c��y��6�?���n(�d'��q�lO�b��twi�]�X�or�Yeʐ. >� ѱ��S�^�iǖ��c��-�/�i��R�w���`��su�;���ع�����sd�������/2Ud.b�;$�߇ep�CzsK�������>]�Yꖪ���w"nOz����T,����c\Ǩx�>(�ȼv��ѓ�t-7F��ҳ���7ݲg^�]����ܠxΞ9�j:�L����Oω�� q5�B�#������4%��Y�I0}��U���wN��ǉ��=�>��K ]�T�9��nG�)���P6R��[Һ#T����G*c������颀Ō�xH��h�;Y?������R2,`���ܪ5W��e8 1׃Y��e���w����.�sMؙ��k��! �c���%��o�,�"L����}f�6�����e��fi*���r%+��������Y3�.+�QA�>c��|i��aq�<3m�[J���n�U�_�e�>�>�i�of���R�O�6�]r'L�>��9}��Wۄ��`@��?����f���2�K2��gӎ�%�Y}���$�}'E�ah�o��B��Պ���	9ӻٺ��^��Y]WznS4wO�Ap��Do�$�`N�N��W��ᜍ���ab�Ҡd��m����1VѴH���D��Y2;@��Μ�> ��L)�e_0����(���7}s��{�� H��+g��]L)-}�|���7�zs!S�9ٱ�� #�e�rc��Q�[�fԹ��+���^�H�Qp뿬��p�<���x%�+�����؅��~��m �q/(�Z�q��0�����//��2Ź�]�W�FF�k�?����pm�-���r}�d
�~'����ǐ�ض�@mo�H�c#�U��Eb��B�̦���`�s���l�tU�O h?sۺ���Me��B7��������N�u]�&(���eп\X�nh#(����l��o��E�u�=pC o�c����=w���۰�7@��w�����[�m�i�H7%c����9V���U��1I��}��'k�d���JR��&�� ���y�E��I)#�Q^najB~^�\E�h*ڸ)\��}����K;h�̉�IL��YT�('f'�d�h�5a�4���ږ���c��U�D�yˡ�!pp����zn�܁��if���ť=����"(1bۗ�W��2�2C\�� E(��A�f�L�fy��B���z�U�>ۏrQ׀��=6�3&m�",)Ǚ���i[��ŋ�O�(F�L�~8wvv�{�]4ˤ&��X�>/� Ⱦx�bs���`�����mj_�2��z�L`��S����
@3�����D��K �.
�� �l�6ӝ���R��-ڌ����yfc �Y3p=�
.Jm���$�t��~G�0h�k�g�͛�o�)��A��,t��@\0nЩ����Z�3��G��ꩡ/o��(�=��=���f�;���{O��T`��#��u@p�֪�-22��H�ɵ���[�������$��aW쮼L	�enӨ�F��� 9X7���(Ä��M��;He{�`��y�2��'�3i�_�Wϼ���H���,n8�,7�r����M��eL�Z4w���,���0i^�Զ	�e��/e����\�)�clt��#�����S/L�<���3�Ƕk\�g�2jx�;}0k�z������eaa��Y͜�2�>e6���K}y�8��q=0�+�Dj�S�GA%��8���>��3��{n����)�m�N���,������H+�@oU2�Ǧ��׼��v��dÑ�3ر7��'8��MN,G�+uB] �<H{\f�s�cA��LȪY(�eLk1�)ւa��������C�w��0�n�����; {/��M�:�P�;:�Gwn���	��f�:W�Z�3d�E]=nY�;�[>Cf�Y���g�˪,�������zLύ�ZI��Vi�,����/�E��rg#}/�pa�����0�<5(�����2�����( ��$��ࠬ�����E��u�c����s������3��� V��9O3?�~ۮ�5aʬi�2����f�5"8B��*�}:�XS���*��_0��_�O�^(������4Z�=3.,��O��"���$�o��J�>��?��?[���K�Z߂7�����Z2��dT� m�Qgnb��d��@��T\���)2������}�5�o��oZ�7��tm]���Al���3��S����~W�A����	��bR����"�������3o����ĺC�2��&漕�w�'��Ns�2�K��V٣?��:r��BV����ɔf�(�����{Z����Ap�rv��[4������M�:ɰ�xdXP���O?����f�A�?�͹ha�ږ��ۺ(퍫ErT"1��cr�����,�Yl�R�*����Ǣ���Ud#����m}��DZ�![�����	&T�F��z˭MA�?ߣ`��6,�u�������)m���d�ڄ���淺uf�@MB:A'��t��DÒ����I�k�Pq25��@����c�EC9w��(�s��f�� *We��疇�ܩ��g�ɱ����0�g�<A� *��9ss'��!P���Q�y�,pp��<�p~� p��!΁���G>2�ц|� z�`Py�uG�^�<@4I���O�&�3gG�ob�`;L�����@J�O}�S�����l�D�7���� ��?h̥�,��Xe�)��2�E�d]=>�Rj�XmK������w]:���~)@�<��е�,�T�������P�����q����~�����	z�,�l�����M]�g�G�������c��LwA:����_p������/|y�G�6��5��C���?Խb]`t{k:��^�[����K^�zLa��`3d��ÉU7Oݫ�r�Ç��R�9�ʢ�C�׃
��2�8��r�&�tN�Yi���;�deD/
���n���0q=��}hr������/���0WL2�hn�j�6�C�8��dJ���fQ&Q�}q]SO�.X����(�)a+����k��o�;��r��.4�U|{�$�$�usb��A����쭉�[t�<�
��h�M�������'`r1Xe��M&/�4�`0i@cOZ&�cl����3��s8�g�(�D9Y�hb��|���nR2��l�F"���>�0θ$|�;�i�+eؒ;k �+�+���k�ճ�>�^�ѹ��w�r+\ g`����*�7��*�o\W�8Z1�C���ۋkӞ���#Ơ��ʖj�hmqzo�lw"�)�ޚ�ö�37�sY���gRw��z�]u<�ܶ{�j�� �p!( ׅ�7.lw&L�j��p��0�����nvּ���K/]bBd�_W������X7�RV�G�fG!+ӚaS��ϫ����+gQ���خS�=3�>O���tN�;�PB��q�3A�d��6,�5�AI�z���f#� �[�"	��T����q�e���@i_�TDD滰���o�B����i���O d�M?��5 ���\}���NI�@UH��\�%��s�Ҝ�ӕC��Ly�k.N0� 7�۬g%'���X]��=�,�dX� �h3�3i�0�]�D^�i#��bL3�=�fW���tu��	����Z[^���w�ֿ��>���}�eN�>mǪ`A���n]3 ���ַڵ|F�(�q�c�,{u�a�2P13� �݄f�#�� �M�Ež��e��� ��(o�7��ǹ��ά�k�	���I�WW'��c�67���s�t1��0����LG�./.l�[Kց�p1����c��p���s�G?��ySS��� ݘ2�"I1�0s�]�a$I��]�ή�G����Ƀ{-��z�2E���**�A)L�(4��J��4Iq.�~8f�z���ŋ�0K��63Mɶ���!q�0�Lq '��ߣ)�d��q���F�o��~�2��@��ʮ&��O�KS��2	��6�<ym�*����zہTd��-�.�������!���xs��M���,�\Uswf�A5�g�{'���X�x� ���p�A�2LF��u ��3���)���� �w��.:����k��
�P
���P���%p]g���K�B�k��`���NӬO?O�e-����`5':�أ�dRn����\��l���v<�뚹B�ۄ~��}֭B�*�����:Nw ��xu�:�\Z.�#t-����˼V�{����K�״�]@�8v�f�fM㔕�� �7��5�a<C�<>��,�2u��Ȭ5���������.�e��E:g�!���\�O��
���D�L�Q�(2�&R�-���2��FEg�T��#:۬��U~��_nu���d�c�D�H\���:���+rq
�����dZd�dw��3�@�k�.i��#i��oˀ4���e��I�(�����5�Ϲ�l%�SW�ew�wv����t�}}�N��Z�������m���L՗�S�8�)5e�kB�޲��{26~<�@cq����.��,uc3���Bi��|�2!�W�nh d@/,=��E$��N������vLĻ������!�8 �qK���?�v>k�NW.���P\TT ����j��M8ʪj5�{��/�o]S�����\��š�ל/;i~X��ڇ�|�e����Ē9M3��t"��QY��� �E��D-2�9&S�$[�B�z�o#i�pQ�)��1�H�7D��W��ko�k C?� ����J�Os��o�����W_�l�:�$!z��2��.���BY
pkE���pܒe9�2T7�U|5e#�b&T�%b��l̈́'(Q�s,����w�󝧆�l�d�IX4��P�s�噷3�ڱ�OO�+YM�N6iN5��D?`B��G8���hh�~�S������d�x-'S}N���Q�tO�&��|��K��̘��	�~v�L�;�Л���I�f%�|*�|U�P ��>����n����k�Ā!w�3 	��߭`�w�V&. 339z�����+�����\��AY&�q�]��l������y纽�P(/�S�������������׿3e[����R�郛&z��da�>5@�"���'����E�D��;M���e�ܶ�;���{^�A>gu	�����O�_��h���DVI&��U�䎹T�%�d�k��#?�S����+����~`|�n�(�?��3��/����_�2�*9>�Y���T}�?�W6��'n5[���Cz�Ͳ��yɿ#=�=U�~Q���&0�ѹ��`p1-�+4���l�f}���/���$tHSq��$���I�VS�~o��1!�;�+ �F�xq����)�}F���bv�ٚ+Nb�A��~�m2i�M��}>�u�͗�����+�F	f�Hp���o�|�X����Z��!�6� �����1`�,�%�D3����Ƙ�<���4�L> J�1��t-Ȝ��g[�kˎi�<�����|����. ��߳�����s��ӵ&'��G5�X������Nb@��었㳙�Oo�YZr�)�ʹY钠�B~�n��������Eq�#��Ww]|�\L���o=Ǿn
):6����+����ufP����xw�A'1G���{3���ۿ��ql�������ʻ{%}� ������V��Z�W��:R�Wϕ�G �s��{V`}�,��k����X�����QMk���[�oY3:+��������ia5��xg���?�ӓ���I�r�x���P�����
�f }2�RL'/���l&�9	r5Ïl��>�K_�{;�m��q25� �I�\����軹 ��ze ������fĀ��{�������9ⶢ�5A��Dɔe ua�P�k�k�P'��zKc����4{O�-͹	pSi�^J���Sk �	 �L�#�ӱ�l�m�P�L��8�:��&�7��gL�M�U����`�{��j���V�����K�5�C��G�)scZ ���񝁗<?�Dݘ�Y�U(�(��݀��S�xqc��Z���J2���)g����u�l�L[g���\����� H�Y��M�Mˌ�������u�~�9W떑Ǥ�0�5�1��d�yQv��u�����ԃ>��G���~����x������~��A�� c�m��w� =�VA�a1�2�o[�BQ1�"�`v����y!���l��rkcև]���X���*��R��� @�܁�,/
�l��a l`�arz졇ڀ�C�P�_B� :h'�;� (Y&���l��UfS���1i����i@lw [{	�@\�ȄL��v2����w������/}^�g��Q�g�[DfM0����&�9 j�7YM�՗�r�O�q���ֱ,es����@��=`&M��"!��Wm�5���~'F���|d?��϶q��z`�~�!K��p5�. �]���Q�G���Q���.t ��7yu?�O�w���� W�d=�+/�����o|�tg��0R'��=.^�"ﭷǱ��n���V����>[k����wN�d�/YT����b��� @���'��M�?���<橃n1��x�> ����Ť�>�%���A���l�!	����7�>�:~�n��MP�pu����qU�mX�#	�C����ӯ��5�˔��w�s����2�T+V��Z��]gq���T��>_��\�ߗ�[e��ܰ�ܯ��GU�S�����t(*?���I�f�n�8�<���A�<���>��O~rrה��!��Q�\ph��)WF6& ��UP(h�L��D2rm�;=���!����~��;/&���߼j���)#�4��7�j�]��~˛>��lp�9g=��
���Sl�<�a�vfd�`�4Ѷ��2\���u4���E�D+��d5����@�
Y����>� �e�'��D�K�Ц\7]x^��}��q��L�h�e�b��
���?�k)斠���M6�1��Z���}>�x��{������9��3_r�4�I-���(3k�YA���L��nI��v4q�J[���[���`d��������D�����2��\]�,o�s�+-7�+�.�IY�Ɇ�����K?ŭe�����o�2���6����<�����A�g,�i&���h?��L/�Pɗ�"?�^��a�G�%�8E.�f����r1���w��*���|=$h[�cy���o���W�i�tuƪ��L���rM��EIa6�w��{�}b8���rW�A�����5�	CR,���xdV��̠�����v����-��d���U�\�s���kc�Q���禛����]�n����J3h�'t;ޜ���� �dv���͖�u!G�My&Xm���d� @LEn�"��9�����*�9A�Ep!��vb�i]����`��e�ڏ߰�6ܽʬ|΅�.Zl��z��Eӿ�Vhꕬ	���=�S�^�s�u۱��Oh�����%D�����*�3��]�\t���O���&Md<5�rl�ṉ��G�9�]-iw$��j`��ɜ��3�eM�x�9��U.$��5d����D_�ن~�Ȱ {d8���|e���p;���8<�����:D��������q�2K�X�
�\L��P��Æ� �eV�)��o�� wb^e9N���e���UdX_�{��sJ>��d�bw0��������zO<��s�}��؀�%2���A���3���U��.���8�}��ߗ+�8�1�N*�&�
����	�I��)�\�7&@ޝ���ֲ�{9��S�c�\���։���c�[2CB�`�dhz#'�LP�[�
p����5�";�	 ���
��cljA;5n+a:6)mcz/�O��x.�.7а���s�w���-��,��d2�.��v���_,k&�Gd䍒w�
\����u�`����ʌ����q���VKR>z����|`���u�жȺ2���΁���r����g�g�.}�q.�k����X,)e0g��B��0���l���Yׇ>�h�߹a
���<��6��4���ֵu�b�ԇ\Ӆ��n��>H+B��;������tx���f�YA~��+�_��o������H�[!��\�2v�?����ߓ����b�
8+Ȝ"����-;��s���2�d6u���C�ף����*w�u��0��l�c�&Vu|��
�w7Ƚ�:�r��{�ybX�=v�}�m̈́��4L����V����Q�a��즬#�D�RM󑌈Zk߭����IS%��d# ���;Z0�93Qj-��<�e4e����)���?���Dh~P��o�L�fn�j���tO*fA��
�����Ӕ(���z� ͞�\U�.�^�`�	ꃲ1!��|�;l�)�L�#h(	PlcXG����G�r&"+��i���e��fP�����;M϶��V���ce��D�ߧi��s��,�\,���/y.��x/�Xv���䦋@��ԨmY򶘽i/HPPS�-Dk�a}[黀��/+��q�b�n��Z����ߚ�\;Ӛ5�ӧc�.��|��8��k!��֝�zu�$�.����_>�w~c��'�1�؃>��{Ƞ�����q�GI��H�q��[7�q����*S���9�,:oJa����o�E!SFw�M�\'�Et�q�*�6ML��V�a;Pm��ކ��ɤ�(& :<�t~�ou7#W�(@�<+�����u��c���7��;����9��3�4�B���
�h�;&�u�o!#�i�l�M���ʰ�`�3Sr�_DSF鏍rskF�y�'�1�|~>��T69�F�S���>��*͞2C���3�d$#���a�/�B����h���=�SU�S��Ej]Pf@"唅��÷�����5�X>���ܣ�{���7������p�����[�~��&�@�lKKC.N굳nWу=���^+M���|n��,�(n-�l��� fn�{u:����w3��-*�[s�g�=p���?ˬ���&��;�����9}��n	YO�촒0��[���|�tepl��g:AYm]VrA�nHw��ҤuH�b�tQ�N�������b���|�;�=��Û�gB���%����\@�s	�cu�j�r؞	�Va-�"S��b�\N���`�j�K�����﫲��%�^�ď��S�� �" Pih�@Q��f�dŏ�eŧB��ʈ�p���ET�cä�Q4s��ؘ�a�9?(�6�RQ ��U<�c^T�Tڑ�#m���~���1��V�^.|<N���t\MٙI!s�f�ĺ�����)k���(��?���\#i6wQf]�x��]��j�xeZ����؅�9�x3�1h��F�8��(J�)���m�0��*�U�% ݧ�>�%K�P�
v��*�JO���2Y6ie��[o�u|3�/x��uf_~��{>K����YBgֻu��ֽ�E�e�_��h�x�۰l�0[��m����Q�P�<��0v�9kI��5�-�>�(h�O'�/k����謣L!F������۸�M�q?���Z�u^��1���O���/�,"�S������p^K��La�������jY���ZW��.S�)S����[E*;���zlD��LO�m���ʗ��Mg��Ns�`����KǦ��H3X�����n�����=v����+��~���_|�����doNM7_��A���`+�G��`��������9	9�f��F��[`#L��~��4�gN�
lL%8bR% ��m��M�d4Ќ��ۀ8?ˀ;i�܈.��ϙrZ��>�
�7�C���)�6?��P϶@�_�����3���sƭW��WNP���K�[�I�a2�\ ȤȂ} �� �b�>�.	��S��Y}��|7A�O�Y���|���W��1ӛ�αg��R�"!��w.�dh��_�/~��i�K��s6��t�П8�Œ�u!k�=�1��h[t��6�mSZ��(��?օi�ƅ�����_�Z��\8g�9��jx����?>��/}��A��ɧ{�W���a���0l3w�2�d�/7��/�)3&���{�=����߾�\W���OY�yz��*22�S//�C�= �ȭ�ޔ_J���W����e�׭��N��G3Wp(l�]�,CR���{z����3�Eؚ����X@�c�Ї�$A�&����O~�(��L��)�d0V��f�1/��-Wy�j�B�tnf�-��2�f��WH��ܲ˂q@��P^L�����2L�c�1�����o4�+x�;�D��F(�;����u����2K��f0���֦HoQ� 4�0��.'{�A��P��>������+�0�8$�]��>O�i~�g��w�aqqB�ǿ���7��� ��p.�{֬u��"0;��T�#�#�U�!�"��Ӳ�nN��>�w �������3[�������K|�h[�-�6�YNʔ��|�����Ⱦ/`t�(�e�dƅ���젧����MI��k��̂`_˸�6nO�u�}3wy�פ,��>y��L��-[�����w��|l�'��¼3�A����K3�cԣC{�pb�``,���.�Φp�o_O�9%=Ra]�ι됏)gfkHOĮzߩ{/�S�M����Vb��|��x/;p::�s��{�~�$P(*1W�Lx���
����� ���;| J;LL�E1��8�u�Ne��ܶΌ �t L�$��6Ѕ�ň�SeV�TdȨ�f��Ou;0�M� +�I&�3��2�Nv0��&Q'>]b������N�*�\�)��=?�s7��۞����Ա��M�"��Er\��2�%Þ�2�<�G�=R�Q������i멟�y��qq� FQ4�>��#˯^�U�	�ʹF�-zƴ>U��҆>�9�]�i!H?VSmi�0��7��V��+��V�R�����:>�t�f
ԯc$����r��;�d�s~HV�zĶ2\�����|.���Kׂ1K�p����̸c�`Y]h_q��s��b�6���p����Ġ{��?�'r	d���#(���:KWǻcSǳ�y����)���O�����)=�H_\�2V?`p�� _e�ȭ�t���]/_J:O����+��+m}p��_$.�Fޢ��A3����0l�s�=����n�x�˿��?jE3����/��g?���3�<�m�|���'��;��S��~�����Ek�i��f�^y?��/ � 3 $M�\�I5w^s�M!����i=��%�A?�Ԛ;5���Jz��ڧs�tAGYi'\?���e���۳�,[���]7-FF����,N�s�*0n��e���F��,}pK2���K�|i�?���4.�c"x�����?=�TOG��ݣ�ײ�eES�����tv��!��	p���?�tK��Z������c�[O_}_�i�kɈ�Z<t�q{e��1��E���~�r�Ԡ�v�S��^��W-7�o7{�7�`V���U_hy��C������9?,� �cw�}��ܓ���ϟ���>k�C�#���E�7�A�t!�[QqA%���ɢ��c֑E֤�\���_���B�ײ��AzU][�G��
\����g�j�a�i'�Q�[�:Dg�y�!"�T�>`�4��C
������������>��� �ѱ������o��0ɷ� � R8�ߚ9X�"'+��{�\�n���`��rs�^(.ؒ�[�k��� "3�����Z�Jӷϛ���o�^u���k_������K�$�y_9Gp���������[L�2�{����Ե������ƌs�˶¬Hߠ�<�+��[���	�2�}����|p����&�t��b.�z=ҡ�<YL3����y~]�t�ȷ�ye�1�鏚�t\df�tAI0������b�iwa���yo����ƚz��˶�]�l+D����-�4� Ǵ�U�d
�����^�v�lwtu#x���$���u܈��`Y�g�'��aE ��0�<�}�/~�� w���ɔ0<����?o`X.��8���Ne���M��'U���"�=W�+�]�>��p��-R����C�S�Ձ�R��Ƭ�J���JFMe�b�J�A�@������s�E� � ���~����c���ŋ��1%�~�g��:��`B�ʘԀ-�!�2��IV���a"0�9�1PD�m�J΅1�kSL�N�	%����Y��2$2ϭ,�nj���朞_����b���m�;g��� ���#���U'�h��sQ&@��*@D����b���<N�5 �:��S���������{=.���A��:�B�3O$ K6^����� p�o�=>k2���-�MSz�ǂ�d����7��g��x�U[�YGc {�1�q^-�ǹ�q~y����s[�$����C��	�+�0`R���g�7P�EGK��v�C��.RdLe��E&��F���sm,���]��f�/�%����e�-�_!鮡��mЙ �k�S[��|�Ӎ`������������0�>��6w'3����w�M��0Gӯy�I25v鿓$Sze��Y��*)������>NYT��{��7�1�,�0�S�ω�	=����,�&�[����f��� ��v�[L�ߤ&z�P�ñM�|�����ٟ�c�͠T��^z�K?��O/���D�j6XJ�������I��K+�4h(sM:!Q�(���L�?��.�$;���>��l�G�����[���ټ��:x�׬(Hr2uB��l��<	\hyŲ�OrF�½uKh�C�Rw��:&rL���_ƺN�"K̢�eYk]d���7ۍA<'}%m�ʲg�`+�c	�W����FM���R����+#㟩�`��|�.�yw��q`���fۥ�N���,���:�k.N������M]`�Hˊ�����h.sV~�r-ǻ$u���L{��<�M|�]��Dr`.a��
���5�r�X�o�����/���뮧�����#�,�C�=�g�a�@}��0u�s�1 �O�Rf<]S<O�V��u�벜��U�rT}SI��,� ��St�J���_���ޫgB�{׳�N�LB����Q�L�0^2����'g@mL.
��PZ*O1S��@��~���>���᷿{��@��k�����͊Y֖���`�_c��%蓩I𠏣;>Qo*�������=\��N�+20�Ȕ ׉"M��Xf�-̈́F��W2@���o�тFͨ�x�2�������|���@�
b��~���Rw2�7-S�udU��y�XΩs�d\����2�/�e��yE��~b��L��Z��a\�NO���~zsF���!����~�)��	&�gv<u���};��������]��l2�R@�/m��֞����J�;2��|{��D������x�km3D&��|��dA�b��s�r��{f��o�y��ҧ�z� �֕�&�}:����y`<�я~��A�>��|�	t��m��󟓊�ͽ<7��Z[��T�X̝�� ��Oּ������]t�*eXU�Բ������)p['��T^eo򾩔�`�1���O)�l�ުa]�bW�*�{#B� rݺ�_����n, OXIr�+nZ`�T#���������|�:;\���ub�͠���_]x��.}��_~��L-�b����3r�M�N��ەz�� �b6���8����nU�F(*�i������租�l���N8�Ԕ0N֍�a?���U�X`� ę� �LE�$+-8�n��9_�-��{}�9�ݡ,��:�
[�K�Ɣ`,"8^���h��=Y���l.3�-�%�������t��'�����-��HO���E��Ŝ�k��ԉiM���҅q���(3��$��e6��Y?�!�/ÖQ&N�A]�響�w�z?���	6������C��x"'oZ�o��7�|��X� Q�9]����5��ܨ�π5�*��>�.L7�I.7%�.�u�#��pm��m��z���b瞔���X��7��G�gn�V �|���c�u��hS��C�gh�����Ȕ�����|�e�[�+��U��ߧȇE��0��^Z��a�_U��y�"b݇Nż�_'�8*ٌDWy�����3ln˵y�ͳ�n��EWgl	p>������G���o>9�2���ɓ�ZlPۃ�����/_��۔�TH(K��Q�&�0i�6{u��I�7ʜ:M��b1�+��d�2$�#�;���'�B�C�rO�oߛ��M:;��o�r�§1�[g�=��{�l�f��%̝�[�����,����X?��N��y�F[[��} 0`(�͠��J�E��� �d
�.�P	lz�y\���kf�'X�)L�_�؀)�Z˲lR]VwS�C�-�Ϙ}D����#�>�5�1^�d��of���
V,���k;���̲z��>As���V���!�.F�	p������칳�xul�pB�a�ⳋ��(N�cr�nP�1��t�5�tq���� ]�Ѫ�sq]�~��d���܀�pމLi�&(�0������_`�q������=�z�����Xx�oɒ���:D����W%��]�X����w�l�ྵ|p��@��\���*�If�rU*K������0��=+eLJ�j �l�`3	�D�pa�0۪�k���~��O������༮Jg(��k���"R��l�@Qм�����P���������� �R��?��֍��I(�1�&�v�w8�{H�b�/8�����$e
ƌ��6�F�dy�ԙ���r<�6F��o�5������[Z����7v�Z�ۭ�1��ؚ��{f]:�:A��"�ړ-SRA��uםX�k�k���{�:�,������Z��ZW\H!5�A�"�F(H=F`�"��\p���+l�e}x/Ǐ 0�j�A�2�.h��O�:�\D�y��2�F;.<���[�|�[��.��c+��8%]\d�a�n��{#�2��q$�]��9�9@L9X�{-������0�ñl��׿��t~��
t	��q�?���aN����yA{�:zkk��oA�����`�����10��0@v�ԏ�YG_�H����|N]��2���.���rX5� ��1%���{����d4�X��Vfoe���8�#���*����o�g����E)2�p(~7�׀�0X����XY�p0��?2(���yR��:O�Ii ��d]����^;�� ���/��.(�[��Jp��P��nA2(Y���sS��%��8���'�L%�.��;�!��)& ��"g����W^����oL�o���q�����w�^��� M���Z��]���9�~4����E�O����c{���'�������{�RMV0��:ʺ��
�[&�؏��*�"=��l�����;���G2��׭ υP���Mn���6Dwa��`�AW��p����c�J�>���d�g&�\�]Sv/�T����nPɶ�%J��05����{ 2]�2�L�	����o��F��7��} m�1�cQ�����s � ;��|�Nh��A\P���F� t������97�-��k��|4�߅����2_�׶��\螢�.w�3���w�w�����͵���QG��g���DV�&*�����q��޲{!��U�*������d��r���g<�����u�O��L3d*�\�/�˧?��v��Ŭ�ﭹ\P��:BT8($M/w�u�6�ǜ�s&��a�>9��s��5��\����Z��rax�+-Q�K/����p�6��߾���u����V�6���ꟗAy|����3q���.����1]�7�g:�ml�RkQ����j���s�{ڳ�s�=c�\�N��L��dJ���r��+�<hl�<��=3�~nڝ�{�xRI$���|��;KY>����^�wep��Y�J�kf���>��e��X�^V$S�q�m3.���U�[��=���Y�P��*�2��z� N��J��i�/�_c�}'�˺�9�q�>�.pu��1�ci�g��o�58�\L�kEf.]�#��A�9/0&o����w�1f���P��i.S[7��:J�S	�}��D�;����re�/��k�Z�|��n�yd��
@Iƅ�}������k_�ړ�糃�y�#�ȑ�.nC9.�B���w����^��́�*�g�c���:�Mdm%Wpǐ��]�f����p$�u!ߓ
�#�M��w��bp+C�S��%ST����y��ޏSzׯ�ϔJ��U3�������P.�� rQ0�}a�FK��4q��:������?��?���t�#e����'�k�vR0j(���O?}aP��� �ѕ%�=�՘�	(
j�XW��#N�փQ��W7e�X�(�x̝˱\�{9����tB��v����������}��<�ܟz�y��A�1Pfvj�-aP��y���'�־h}����JI �1��~�?\�������������������1��{ｷ�S��P�d�S�Mr���8����gO�,��rgS�_w���7
�r_�Iy��i��#2��Ғ�ں F�i�q����dh��Ahf���dk���m�]�gX��>C��W���n�8>�=�y'�ܢ���M�z��k�ڧ3e����m���������<4 ��
��C�:����������\=�u�㝧A/`��j�����l��������e�~΋n�M��[6n�}�;}`kz5�a�=.^���}��>��޸����R�zO�ԅ���>N��$-�#]��e��(+�� \��+[q���u���p�&H�/ K�Y� (��g�5��w��w7�����)O6��@���|�`LV`�H=�-I�Nى�Ք�LNT���J�����ڔ��̭4�ٍ/(' R�>qJ��q x~�;����V����?'Z'͏(��~���~�
��q�坺5p+'R��t��y�|nO��3.��'.ˇ8�cB�MjU�%�e*���th�Hd����ߎ~i�$��1���sS��ݲ�0�޴�~��WD�b{TPR���&k����R�^��������"���5i+}#&"�@-�7 �wsF3�6�~X^X褤Y߼��+�Si���y��jz��㭀DSt�����l?_on�ۓJn�)9�]$f��ԙK7
a1�Я	�d�{�6m�����}� C��Jb R�Ԕ�!���΋��9�s�{���b����
@w���,��OY=�j���^� �/���<�e���8�$�-��̓�6*��el��&�Wީ{�qS��z��^�Y>���7߯��M5F�|��:��#]�̎��^�Y�8Ȍ\�x�XݾWS����ߔ��r/XM,���d`���*�ia��8�V��.\�	K�h�2���h3-�e��T���%�.R�y:��	�	�k�ח�B��|n>?"��[��oZ�0��F2�o3ew����FV(�4MQM��}�̼0����.�����>O��7' �eΨS�-whs2��� ��|ǹ�1R���/6��o4�7v�`�n��1yL�{��2�����ZƩ�寿�~<E"�Z�u���O֞�����>6���?��튾,�&~�2��C�>�p��+��Ŝ�Y�'D}�j����Ӿ� J]�>�YW.�iWoZ���d���!D�c�'�K�E�X h
�.k��s��1Z ѡ�_ڐ���c�������62�̹-�W$Bx7P�>���u��`>��	��@Y^�,�V@I ](�k�@-�����=ԥ�q!XƔ��S�_r}���������n��Y��S�w�Ia�5*^uU1U�e��u^Y��2m2P�Q,�xQx(���o���6�� u�K�3*��Oft�R���� W�MF4g�j�E�Q4�$�R�p��p���=)��&��5�yܢ�kq/]2��2��J.�[�=���3
�~b(NʼS������E/L�2��]�6P��:l���ߝ�K���-�s�ܼ� ���nN�_�Hu�e29�[Y��F�c���>�N���~����}�s�O}�S츘��@�e��2B�d;՗c)Wl�e�5���,�	����-��#� *��N�y?Y�
���y�̜Q�a^?˃��֍��v����[�{���:.������.$󙓕�kib��� &�+���a�t�xŲ���g�L�x˓��3(˱��:����S��\�t���QO�i�,�y�S�x��ґf�Â۩Şuo;�ϰ�mI[ ��k��`�����ϴ�.&Z'�o]%�۶p�l+�S��-�o���d��:G�L�i#�,�'ο.ڙ{hXk��s���|�U�[�+������{�X߫`��1��=��z��d!���|��Ez+�ED����d��7BrbC`9X,�g�̨@@a�
����U�@״b*T�����ٙ�(�<�H��9)�`T������5��I�g�{P*x��ݛ��3b؝� I��2*� ��W͑�i�v��@$3�g8�1]1q㮀�7���-�ɯ��tY1 ��S�>�9�5HGv;Yl��I�k��{����gs�п�6�� �S6&&&
|n��[�@�]^\�+�y���C~��J�ˬ v�E#룂c����\}b���Sl'��5�~S���e@������S��� /��U*x�uX����k�4�}a�h{  �q�����c�Q.�?��~[��� \�����I�SJ�6��;F��.�W�m�)-	���p��@��nK�@�z� 	��.��E�a����Ş$��Mf>�]��<�>�0mAۣ�h_^��<#��>���3�>e;�/<��Y�I� �0�a��.��{�;v�]�`ݱ���~���/u��ǖ�0�ޢ��a�e5wY[�r\OV����8m�<��PS w�U��{�ho�������g���y��ЂS��$#�Q�f�4&�r_t!ʵ:�3��\�'�M0*ӗ{��v�mܛ�U�*J��N"<��(w��h��ꊡ��,O��e2�:��"$�Jֲ�a��Q{�W�����w�̇宊��eҝh�Y��8�~������	+�޼W}q=
(w�.��I`A��}�����:���|�3���u�IC0���ͶvS����Ӊ#.�T����WAZ��{�{��t%���[}�+��wW'�
��`�'����h�j/`�k�ZZ����5�U-s^W��0C�����<��'�~%�e<�zf����95� ���b��Z���C�5�~k�;�	|��z�.��R��P=���y�V#���pZf�iG���C�8��,S�^�UV�w�s|X'�)� ,���9Z� �}^����U�o��]���>��F���
p3(QZ^�B4�:���ӥ��2��G [-pY�JR�.�a��s+�,�9Sc���[�?p=�'s^$� �(����e�1u�E�h;N�=�{b�ef�@D������Q�SL)L��B%�X˒fG_9�%[(���\�
bL;�bw�(Ut�iԢ(U�����|~���	�$%����J�:�=L��B��LP�6�^(y����Z������D�/����]���l�b���3�2i�3A��֨�[�D�eϻQ�>��>yLnw�~G�0y諦o�����>&���d����+������*uҬ��ϕ��(}�� �ƻh��XF-�����!Х��Q� �A>gNF��@��$����ǧ����~M���5.S|�bCS.�����(ʝf�l� Ew-h��A�^#w�w� ��do�f����B�������#s7��t��U�UW��;︳�JI9�w3ǌ�$p��u^-�\4�,@�-��i��\<��Нγ���g�wZ�I}�2.����b`��ap������.�̕N?s�eߐ����̙��u������C�*�2��s�:��eeYv���S��w�Q@.r�g���Nf)ךa=�,R��u����;�w|o���y�\�9�d!*q�Uo�(!�$	�z,�+e'i���I݉�k��&S� *,����p|�K�ѷfcH0����w��1G��F.>R�i�2��I��(L�fU�:�h�����a��[G�n�g�1K��>�n9�)�- �o�v��2EXF"g���3�s���t��i�l&�����N�6�똈��~�,�E�R�K�RM�=��Z˄�Q���۹k.$}e���f]x�רL� J�R���3�m3�ϵLۗu�u�>p�՗̾��� ��{�i��}�>�+S&;451��L˒Ϫ�(�6�vO��Ĥ����e u�x0�5~7�ߺ`;�+�r�x���[�6� }�ŗ��Ѳ�8�����~��-<
y#��_$��Ϥ.Awh���w����B�ſY#L�朢��m���D�&�k�h��H��J`����%�9��f@�&�֭.��dC:u�2�X��q�o����c`SV�ǅ�pk!NBe�d�r�(�u�Y��^c�o��@M%�F�F� ���W?V���W����	����Y��Ʋ$c��prBϼ����V��Vb�6g�X�%�:��%W�5������X�B��_���l���]�`/����^5��[}3 �{[��t �l"�+���}lA���Wʒy�|��es�³	
xF�e�p�w�k����я~�M:�C�R�id}�oe4����k�l��%�g�@��Zp�S $SR!�h�k:�r�9�Bd'3#J�9�L�
p�i�29��\�i���L�~��i����\ �K0k*C��@²�3/mi��\�S��;:%U�!t�a=Wk�@)A�`Nl.n���
���짺U�G��iM'X�6��������[2z�)X5�k�1�"!c#x>�ȍ��t�]��j���s$��3��:Y��|�E1b3CH�P��kK`�BO����s�e�À�U�S��Z��E��Q�;�"k9V�0 �h�pe8�
l�P�^��L��'�L+�>�_	Z��,�	��N�
�]�FK����i9Q�(yb�1g�Mw
��rKW��l����RADO�UR�U������3X����ȠP�E��8!�R'��Up�w#��P�ȳ�i��`�3'�~g�[FM�	d�ꋈ���cae�5	��*�� ����ӌ.[��P�W]rR�`��i��=��w2�~_�&����>�R���W�veu��c���]�׿	���&�M�]�l=�P3��Xˑ.J|[����7��a[�N��e�������k	}K׋�g��׷,��z��c�4S|��.������fO����V���5"�B�ml����q���^��/��8���W���t���@6�`����d�0 l��Ԓ�zV���O'�U�����A_v���]C�Y�Ofee�@�'>�V�^i|y-B�O�q<GŇ�²�D�pon�<b�Ю�U�� �>�)�r������;|�	����v��;���ߙ{�=����ƣ�0�F�m�܇���
KDٵO��2ej_�V�b?�e 7vT�=Ǆc�O�z�iX/�����+�e�ګz߅�Od8����πd��@u�˻ԀM�ǧ�l6@	��4 �u�%$�3���A.eĢ�u��XZ'/��r+�o����tG(�����O�,MRM���&`Y34������+V���;N�l��G���Cɲ1��$)���&}��ch4���� ;*�������䏩����PN��Ԓ��G�-����
 ��Rtш��c�����[l��I���Y䱊bǾ���g`'�s��F���b9��7�Яӳ[ʱBJ���jҗ���m�%�/oe���E����ӫ�-�B�b���ۊ�����=�+,��Z���J�ƕƚ��\���[c=+y�)iU�왌G+ʔƠ���ҷ� �������nGn�E�s��]�P�X̕nW���Y�e��o��u_R����_#�Z�9����P��n�8W����4so�� ��}-���;��v����z�/�.�����q�ÿ�G�8�D=���C�Ab�����I�71�G��p�^X���q��o�r���?��R��S݋��	&K'���eS���vk�N���H5�� DD�h���O��2�o	]Y����Ҏ��B�vrk	�o~�[AA/����s���bp�a7��S[їԕ<��[��_2�"=6�88Ǳ�[�/�:h����x���q	p���^ک���5ɕ�|3i��*�Z��0Y�з�B�V!���կ�@Cuq%���#�J��S?%��Ay\Z\,��ҷorһ̩�����&Ę�U�� �|C�ڀ�c�����ם~i�u�z�zn��";�ߑ�E�sڙ�	ɻ��#��@��
�
?�@��xb?���N���^�o������D�XBш�S�2��)������ߕ�xa��gVM0������urFl�1U�Q�I"�,z߭�[��X���}�9�<- �[F��q�Wz,呦�}��-f�7���;�Qf@��G���g�I#�1�!��.��f�%^����	��:>Ҹ���t���@�%f?���U�k�U�U �&�N�Oh֑Ҫ����s<ܛ^w���!�B�c��y�2~�մs� z_zvŋ>����c^�&R7�1��owM�=�<�HA�k_v�,Ү��e>���|� _��&M63EΔ=�uwa��{_R^R�� ���nޔe+6�x��Z��VA���rRO񽮡��#���2_i�8$&*�����#�}NĂ�9���"u��Tl�	���6s��T-��@
�c���[��M�4\�/����[� eq+����SV�Ee�%#2\�O��a�*�L�feI+�뽳Op�ZpG�v��!)2HG��&Qg�8������1}]�#h���T}�?NHY�N��Ǐ�՗I3@��]�W��-����jC���'��M������.|�t�D���[>�ֺ��ux�ui�u8k��nq|p�@�|�h8������vEEh�����e��
Tf]�>��]�E˪�B���-�?��C�O7{�wǓ��I��2��[������?Q@{y��_��g )�[��uN��-��r��3p����\N�o���oܨ|	=kc��s�#���㋺B��)·=�Fl�l��.7ZϷdbOY� ��UKv���j���B%oG�}V���G���^z���]�a�`��s��i�e�Mf���'_B�`p�Z��6�Y�U^~?2x5����ݷ�-�e�ϟ���78��\[���i{�	,���T=�� ��
u@��HK_�tK��E����/��MB��R�ۊ�}R��Bu��xF�\m(�,�U>�2���[��Ҧ�v����B��c�]� �ri�@ ���|��	܏�ļY���~�YT
�f����y����y):�?�o��Bg�l�7F��$yw��"�7�<��x �?�wloҎ�dT����9���y#sbk�e`�ө��wEт����v���St2EO��*pWꬿFeD"���x��ki�\���r,���Jn�v
�k�E-���Ƞ�p *�&�,��A�2T�E!AnHzV��d�{D����'�0�zV�֟��I`t�������ˇ/!# 0V��l�U�}D�ZTrzm��Q��Y,`# Îi}�7����M9"�n1#?��=>���z�|�-|t��D�a�2�!&(vB�t�с:mO��DҐ�ہ8��������\�,���v�Ǔ�|�S��ԛ%YiE�_�K�Ԗ��ޚ7[c-��#�KН����"��~a�G�
7�e )+{o��l/�ת9����Ɯ8GWi��/SX[ 9^k�;�gV~/߮�D���*�C⭨��2������^�=3p�F�ڣ]J��4,>���^� �	1�Qk�u-ZvH��!ŲG��,)k^bZ��ր�ẉ�LFk5��;U[T�<� %���lo��|k=���G�����u
��F��|�����ߜ9{��5�#�E��2�r�3�C	P�J�y|�4�K�W�7\T~@���ei�|8VeS�؉�����y��m��l8��:���T�9���������7��z��HQ�gw�o6s���)ں��:=��� ��Vgw3����^�"��G�V:1A�vW�Ľ�{B����>�����Z_鹫Blc[AY[�h�@��l���Q��۾�V�+�d�z�"R�3�g |my�P�(\	6��^Ii�!�[M 1�C4�H%2 T̵�2
R���z7N�k�#ӼG��ʪ1�uf��Y��f՟�6����Q���]���{D��Rr�N5�g�������<}�y��+��x��mϨ���"�'Xx�~��K?�я7?��O���GS�{��L\u_y*�q��di�s���$�T�}�<��	Eytr�7}�UF�Ot�2;�h�2�E~���~���|t�ǔ#�u�ͅ�'�m$��q��K��� �S�t�����|�;3��s��4�e&��T�c�u/S y&�m5�e 2kc��ȞG|��q�����go��Zk���:W�h�\�d�.<3�]Fxn�<��(`o忄Z�m�MU��U��ڧG-��(�6�>An�8yCg@�ވu�U�l��E]�L��d\=��# j�TO����V5�����F��"/�h_�&�}�y�Zm��J(��%�٫S�~�M7J��QW�G������n����͠�}�c� 
�c޾|a����<��g�S|�wճ�@�XA?8�7F���r}d����´	s����:�����p�,K؄~���i[�p8��$�:p�tq������9?�E�_�W��PN�#֫�Z�IO�.Iz�B8UK�x���6��x��wop�|1����B�o|c���V�A�W ��yޜ/��+�T^�w���59��g�=�-�l�c�<(o�h�}/�h�ʰ��E��ɵ����٬�/OLw	(o������NK�{M����31��@F֑� �K��ܥ�}��1?W�&�ޤ>J��֤J^#�l58+����ZZ\֎��=0���^?��O�^U�z��Y)v��=}|�8�+� �,z��
�鞀�������"��� a^�?uz�/Zl���Q��-�%p����@	�@� V9��@2G�����rd1�E�9�`����� `u���16�yX0��I:�OL`{��X�q%�XWNn�M;�!�a���Q�R<�@�ek9va��v���S����r�o���!q�T���?7:�F疘v�n�0{�+�d��)ә�����O�}+�k�Qo_�w��R�������NU��e�#+w5�������,�X�V{�Wbٝ�t�y�_��wtj�*���Y%�j�Z�^`z@�k��e�������H�K�ӮN�6:�V�G��9�?{&{gI�NK��Hy�<v���RO@�_�R����f6ya���+*`l��E�=�y���gN�G�2̲=qM���q�sQ���Q�S.�0��x��^X����N����7Ym�����w��">���r�L�o �3�l$���CZ�p�4�u�������>��ت���D��Fd�BKAl	�J�~v�n��F����޸��e�1J�rsd�<4���F��}(I=l���z.��J�TX`I��d�(���U�-e#>��Ea��������zv���Kn���̑*&��n�٭�w�����`�B$������߱nQ�f໢�ޒw��Y�zy��[�����y����)����@&M���6o��g+�o>��-Y���w��� 7-���S�`���O�����q��R��7n��<t�<��3n���>���Uأ=���f������|���������P�c���R���]�+_�ʬl�⮁rCqLF��q��WsdŃK̒�M{�{�]͹�;����|��a-y?�е��I���]�F�T��ɳJ!k�C�H[�ʋ������ֵ}�+��Fe�5Z��PuZ��K&Ӟ���� _ZZe_:1,�|ee���������mS�C��D�إ��\TJ�h[����v���`+�=#����x{�0Z�X��WXe����"Q��:`�s�_�.١�����hB>g`6���n�M�{H1�rcٖ�~����;7w�q��{E� �z\d���)n��ʅB~�_�җ�o���⌛�����E�4��U�|싪1բhW���F�,���%Ļ-%�J�\W$�f���J9���JF���a��7�Gʰ����X;~yw���>�V�a�A��l�Z;i�^l���eˮg��J�	���,QO`��H>H".�߬����f�g_V��V�5W�3{oi�z��(�
�"(���w�H@	芰�b�$,��|D
��s�=s�gm�Dʂ(�oYl9�U���S��>Y��L���W���6�g5���1/�J�!���k��:b�l�H���l��hz�#�=�/�c\�Ρ8�rK��Vn	zO
Vd�:n���[|�t �n	ٵ�ọu?��͋k���HkA�.�&���~%F�dM�e<qH��.y/}w�P����Yя��������(���:�� +M�5P+A�J���1uƲ�XR�Z}�����O�v�P�W� ��)����{�[��O?��l���X������e����.`ଏ ����x�;ޱ����XVEi��Y���	/e���1[��v�gB��~�>��5��O?SJ�P��o>::�<����߲�Y�^"=���1��IwʗMezG�Y�����oϾ�Ĺ�U����gn���/n�I<�.�} ����{�|��NK�];�Um?��<vi�Keơ?Y��X��C��@F#��i����U�#ƣQZ��EQ��'��5ξ�b��~�����P�,KҮ,�uc	 ��D,{e��ޯ�=
�Z�.~g�ǁ�)�5*���2�V�2ZR�5e�CP��ϕcp��7+@8�z衇f�JL]��x��H�(V�/�/0+&�P�0j���*;������f��ow�ڵgͩ���)`�}=d� %m�6���Gn��bK��~����$58���+��7�����V�r��ڗ�-���|~���l82~[���=C��H���Qy�+x�J�[#����P+�l|���R����J|��U �k�0�d�W��e���Rh��3���V�.��B��\V�V٫<�g	�+��W&/C�Z�>le����-@��,D�m� �x��g��O�?�|K�m����0��(@徜Hr'�F%��'n�6?)��,� -�
�i]l&h�����x�)Mi�#����tp����0_����e��\����^�.H �����6�k(������ͻ���ٺ�1Ĵ��*��3�2?�W�ne	�;� ������c��#�
��R���/YY+E��Z��:R�ʌ:Kx��Ͼhy���ӌ@6����*oL+�#S�b�w{K��h#
`U��7�,�?�d��x?�VǍ�l"� Q�I�D=�&��/�Ĳ�eyĲ�{1Ϩ-e�T���@X
��4�`�ɥ�o���٥
�e}�R\��	��<�y���<*�b�1�L��o|��~c)�UQ@��_��le�eP�B�4�,hcK��K�]6Q����36;�w�}�ӵr�6@�%]O�Cs�i�,>�N8(�@��f��ѦXH9>X�99M��Gn	����,�z��:����X�?.�'��ˇ��j�g�}vn�6���(��~6�g�����8����_6wT�c�#���b��5g����|	Ȋ}��ȥe[�����)���{�|������k�u��ZnG�iՙ����5��c��3ٍL[��V�+&��Q\
��d��*gk�W��ubU�%� ���$@��ſ{϶x�����wU�]&�O��Z=��A�=��u���R�P���rg�fB�*3�P�X��5 ��P����K`M��GGG�;��lBH@`�
�������jeٕ_��4���R?VQ�YЦ�D"3P,ͱ�F��9�RsO�qN��f1�G�r���f2m��u���������Vm����[�4��|mqKPZ��U_8���l�{�e|]������@	�c�����o��}ɔUl���ߣ�|eem/�޼W�'������Gj����6�,�HU��RQ��@�y��[�5�DX�h)P����5�x�J+��K]�POʀ�IN�Ki��Z��7�U�����  ��IDAT& �0G��[|fWMwtL��(�G�l)9��Lq�oT���
@i����,����=�]6�a�ds�r*>��.Ȋ�oemD����������_�:�����1!
=��G6�E-y�9K�T^��� + ��c�p�C��q��1Bu��)8ٌ�~����[���v���V�[i�.}�'�@������X�|�/�w6�DP7�2�PV����9�U�% ?�v5Ȗ� �}�f~�"�m)�N��KK�OK>��IW�Z�Oum��(���6���&�,�]z�~�D�����$�m���2���(Z'\Qhi�1��w�}h���G����(���iD���ܐY���(k\��G��\���u^;}	 �&�	XtP	��5Y���[�-@��j����@�t�,��uƭ����{Q�8�u (	��Gi� �+p+�6jY�j٘��p��.�_�^�Z�[���/y���Y����&w7Y"���V7�e<��
��@t��Z���lN^��V��%�yD1�����͏�J���@n��Q��L�r���3�s� ���::og�2Z�}b�}�.�̂�M˂xhz��E-�7��f���ꤙ�5��{<6ji���X���⡖�a�ݑtze\J�"���	��q ��Uc�~��	D-�?��S3 �2�<Y-�$�='���� 1@������4�V����b�����Wi达����E=="uLS7��^>��2�lzF����0�c*�>*����7���(�2=�rp���yY�e��&2� ��G<�Á���O2B�o���o���H~�g�Q�����v�8�hOw���7G�Z�Z�����\m�g	�ʦ?�5�cT�h���j.��eco���F�ھ�|p��,m��'Q�ky@F��C�����yh`��$5R�� �M
�|F�q���u���L������1.l��*���`O�1=�2h9^ �G�������aA�%S���F�ظ曵��@�,�˿}_��W�:�*�4�"�x&ª��+~���o/ �*��h�>�l֠4p�P�������zx0Ykfe!���mCm�1�ݧ��}_�L�e�Ad3@y#���9�g�6�Pr�u���݇��/Q��-�W�9�j�]�����(/)�#���]�F���;˷�V�vk���ۢ%��Y�z�xT0V��Q�R��B��[1���ז��b	�䝘<�(��dyT��k'1h=O���0��Yƴ[���F��6{?�6k����
�ɢ+�&�&�Y\��Ғ������ͷܼ}_��Gn��	�1L�Q�eV~�hz�������*�T�ͩӗ@��_���xaA~t0!�p��{��F9 �s�ۍ�c�Z�)!��n�0�P_r� ܪ>*/�QP ���+�_\�o��+~�͖e�������ʝ�y����d�[�ި���_m 8*����ٕ<�N���9��w��V<�<���]ک����G'���]��(�t�x�\Y����Z�̓�K��V���&�����N�)�ȽH#u��$_M(�ߣ~`#O�O�,EU2��M�#T�p?�G�H�47�ȕ�*n�����&�����%l�d��o�e�V �>�K�.>�Xpe�u7��2 T����	��4�����3���G~��c�����9�47"G�l�p�b8��/���w�}ۚ�����=�,1�ֵ��w;k@��ղ�z��}V��9bT��6YK��?G+�%�D�-[��C���s��em�H���+I�� ��V����^�4�,�5'�8�T��H����}�Ƞ���ld���4d<���.2PX	êL=M�e���כ*ޗ�Bf5��5�V�����?��x�Y��8��d��q��,��8ӷ�
�-]��ճD^�]�])�Y��Xv�[@��u�+��1ځ��ҋQ�v��7��Ҙ��T\,���wpk ����>Rde�������|����R�@=���<���y!{>�����y-���?�y:[Y�1OO7��
�fT�m��*�=^�)�#�Z�˹F���P�6���m��[f���~n=_���7���G�N%�c�2���Z*nK[��g�--��_J�$n+��K{�G|d�2��U�9���Ů�MI7
�lG����˨ h	�8[�m��+Ea��c������K�UY�5��t{i/?Q��;��a�dy^�M�V��Lj3�|VmAmN�o�@�D P���;�t�ʡ4��5.�b���/ys��V�o-��t��/j�8�[�@��m�Ϭg}FT_����޿c�+6��	����(��w��+������z� ��,�u�VQ�oVv�O��v^��]�����d�6��(�V�{}�uI9��?F�����F�\%�>#���o]z���Ƃ� �]���'�\+M��:d-�\BK�5��*��+Ѿf?���e�,��Z��w3p'�V[�C�x^��%B�g�t�ڿ�������C�����z@W���0;�]���#��o�-(R�6i�Ch-6^�f1���U"?���Ǳ��IZ�,\(pKP��―Y]S�b�ʧV�ɲ�
������S�4�H�vcg}�u�Ѩ k�����w�[G�d wTY^C��^۶����{������[�v�Ҏ�4Z��_w��J������hf�.�s�l���h�T�C� ���
��|F�,�e$��B�|w�� )����{��8�B�X�L�kM~K'�Lk��%����w�2�v�j�-ay:����`dr �V��R��&���y@N�R[Yine��𤋮�o}�[g���w�cvc�N�"�q7έ�\�x���TT�=���3�~ ��ꧣ�b��ܲ��piY,�X�����ț-��k����<�ʣU֪�<[�X5:o�2�J>�Z
����\'I-mm�� Khm�⧞ӓs�sȍ��g��5�GQ�*<�Ļh�U�U/\�]��{�!�*��4��w�(Y_g鸵cDs��riZ��]�m�!f·W�:�����=�Ǔ���G���U{��H���Kx0K��6m�r=��K+˥ ����������h:�.J��4��:�[�Uy���E6f�"�yM~�~���O?=\]�U���J��/��K>Xr��o�HҬ.��zz�qn�'0�JX6n�΋�����Զេa��66Ų��SG���%�hm���[)E�(s�}NR9�����J)�o�'Y�E����CQKk��*�9�J3���. ���g�.��c���=K���?�o)l>Ȗ�����F�}V�x-������񚟼����Ϟ��*�]h4/ WVY?�A������*���l����?W��&0,�ĥ�\�g�7�y�+e��|��C-^��G��B\�B���C�ƪ���ǇW�r`�,�J�`�����5���po{Wz3����O��6�ջյ���״gT�z
pLߕ��?��tִq������}�B�ټ8�֡�hk;	 X�L빥�V2�$������4U�I�;���cM�Z a-x��ZM�K���g�vKs�w������ϔ-��*o�Za�z�yeA��s�Q��������Bq\d1N�2���F�0�C�{Y����ˬ�V� Y8��{���l��b߲��� \���Ė��1��6p^� ��ῦ��2�Ҍ/0!�x_�d�PW�9�A�[Y��.i�r!�ߜ����oqe���O��'bԔ��U���5��r�y��q��=	XW 7�?��D,c�wIp�(�����s��sx�2e�TsR��}��?p^��������#*c���JC 7�}��^~�vK������	�]��(c��_�GL?�?:P��VV�lp�&�*��0��w�-põ����	�����4*�j|/��^�q�`��8h�} W�����	���s-������Nv-�A�Lr��G�q0��������g�}v��b���S@�-���r]VQN������z��Tq��̼�\*����E�x_���@�k�rC�7��S� �" r��y�~|p�?���?|�)|���N��;�r��M�!��X�����Ǽ��Ju�l�(ʡj>�s�>�c�����ʝ���m#m���V�b�vI�dcn"�C���UT�\�_��-�4�2jM ����Uk��Q��qY2)����2���c[�-֧:2��W����f��h�Y9*���Y]�I1��ץ��zy}����p����d�ا`�0m"�O�@��"�q���D�[զY�H�7���!,��4�<V3`�/г��:@���u�[� �>���z3��[��U Y���4NI�`w; ���4G`��/~��c	x����ה�-���Z�r6N�:����S�E���>Ф㱎E���3���~��[E��V���u�Y��٭����l����R"F˵�?G�u�|��m�k>�8�b����\[[��^U�?��29���E�n��F)k��k���dWM�U� �(�T�q�_��>2A� �HYcY��*[��1�pw��x��Ƚl��O/ۈT�1}���9�e����d@QԮ�r�i�q7� �vo�M���RJ-� �7��mh��cգ v���O��X.g���[�.�e"�m�kt9������B��W���m�qX����ec2֡�@+�g���])����J���b�9N���p+� �Gۈsc�ƿ+� k�������˸�Us��੢�}� �>o6�
��<[y��@nL���l����y!{'+�b�
��v�X�*��:B��8�>@�`���@S��K�0���
��z�`z���l$�bd���e��]��a!�~��$	O_��� ,��= ��E`�ᔠ�� P\��Z�n��y;n|��L(F��S쇖 l���7�� �2��UO���3���	8���� ү���AF��(`�z�X�e�k�(�ŏ��[��R_X��@ �[���o�rO�p��g�@�|�����{�()Ѻ� >S^�F�WP��F��������K��!��vX��I�ƹ��4��9#�R���ɬ��2[����0atv��e�z���l��X��Nz�y��iU��z>G&�5�`t2G���/���,A�2��歷�:�F #����`Ӆ���6MI����&%�]���e$]��G�z8h޷b���Xf`YBEn!t%&k-���e9.�Ǳ^�=�ߛsG�UJ�>��U�~�ۀ�@%A�M�	�*�6���2��Q��q��qD>�O�/�D��������o��ݗ����+���fi9[�>�!#J[L�J�Qڥ����;[y����P�f�\Y1�B-��,���с�	�
�FKC�����疤�e���!v��6o�'¢�\����6�:g<Vi�= ��F}Xe)��M� mj���Alh���޸���w���N���x�)!,a� �ہ�L�w"��_	bb�����<W�����>��<#?���g�"`ۥ�n_���PV�}��*?�)��dc9��ܷ6�{"G̛�^����o�}S�N %RQ0 ���x�q�`7�����P�RP����5��~���<���U7�ݸb���)���\�5m�陵)q���ۥ,'��K(�εe\3���^�֞}�ڵ�V�Z�fgԪp�����:]f�=pU����$G4��L�Ε��-��zm����R��o���v4�m~�&�jo)
�����$l���n|�"Gɲ3���B���Ù�����+'��g��2��\�ȗK W�W��X�/<�y��W�K���^�ҶZKK&}��֎��l57d��{4"��rļ�����¾$���L��x^|)�fe`K�_)��(���&�ۉ�u]�3��=������a��[�>������ʁk��s7�/!��Dz���.�b��>84�[+�;�^���!��W���]�ynt|FZ
n��֗��z'���z�e�0\R�}jj ���sKiT1�4�����Ǿ�<��~�]�N���Mj-������:K�VVZ	N 9���J@�����9^�l�
�2���	�{�@2�Y���] �~�# �e���~�xqk)F�+M�?26���-!O��%e��WQ(zT�ԥ�y��V�f�E�_�N7�� �e�C�#.>��1��l$��U�7oR|��7�-�^v���=��(��ܱ��Q��9UO��r�dsڡ�e���!a���g�:i��O�{M���ַ��Y�k�h��~,K|�zfI�����m�?��F���D��4R�% k�=�\�\����[��v�a��p���*���~ϭr���o��bXf�0�<G-`�����K�A��g�y�;߹���f+�&#�j�c���~u�.�|�%�X/ߕ�z��"��*�++�+P��cU���E����7�S�Q��"ZK�ۇp� /���^��瑝�����������`$o�5�<]�_N�'�G�Lʣ���f�@���$ڄ�۲:�!�P�X)A�$�����!b�[`�W�0�9�$K�VRt_V枒�{��1����5i�\�h-`l��$����V��l5��C�j��woTiXtT�J�X�<�}X>F��K�oU��wU��EpWf� \L�U��ڨ��Ұ*�*Sf˾���6de��ȄV�]u'S�O�V��mo{��`dC~�n	ExaAG���E���I9��>�J�4���"��"���T�R�0��oY�p_���c^=���mW�ƈ��ytnq���?~�B��X�iWc����e�Rտꃬ���ߞvk^�Co�� K�]�X�R�[���t���x�Ǖ��\�/��K����ok�*x]�G�'p�q�:�*��,��5�x�w���v���]�Fˤ�3���> R�� �l��z���X&α�3=��r�z�|�0F#Ŀ���G�.��R�c)�,1��RK�Ƚ��#���6�]�^�u��[�L�d��-0R�D{�dVif`���� �������^x���ʊ+�� ���/ �^�D�IVj�n�׿as����l=�ߡ0�	���h^	}6ᰣ\�c	�}"/�~��@2	`aۙ<������߲~Xr�<Z�U��RƯ�ٚȫy K�ѲV�F���w<�_X\op�Ѹ0$"�D�C��
�
z��@%@��̭���{�F��
1s��H�ܡ6"��昷�u�PT�'o��1����2s�h�0�>�{��% 7������d����F�@"-P�di�{���`Z2�2����i�YY��k�#��޳�}��IlD`g�y!N�Yz�ۭI=�_�)rP���X�����q����OkqiI{+�_�p�Ĳ����bm}�����eA�G�b}8�<��m�~on�\����U�/��EZ�U}TW�%�m�eᳲɫ5�*>X3>2���?7l������/*��}���*�������C��a��9�V���'��~�=�� W����p�W�J E)��&�]�⇛�Ϥ���� ����
�w\-T7}+��
�j��y�A_�՛���h��k�f��R$���~_�����ԫ�F����S�nGh)TuN}p{@�Jx4����[�^�|Way���n����,�%�e���ܚ�� � ����6,U�t��j�Q&(�'��r�`���g�{����%	-	X���*K�n5�ܗ/l���c_�	3���-<[Pu�˛ӯ��=��E�{��y� /�9�eÛ�@9���}��1�+ �S�=0u����,$YV���Q@�K�!����1�r-i��^����1��}��ޜ�c�o�"�iLVN�/)[�&BipE�1 �
����}�9(�?u_Z�9x?jc��3g7x�b�0��RB�^����/��{�?�-�ͭ�K�/� y,M#�%޿�@.�k�z�Z�+�1R�?3`���qZi\ԍ�+�������^����/�C&l*KJ�~dUYF���UE���ٻ��o�7�,�Pc��NnՑ`��EIV[�\Yr�!̰�  c��톗_��\�K��_��-�/�l=<u�����+/o-�l��u	]�[�'�4��t����
_=��O^?P��E����֟%�U��=���3��]|Bs(�_�K��|�2���3��=w�����q��b�^�&R��++��I�o��Lvᗮ�����l�d����a��"?���S|���nڂf6�ዯ2�6>���Glk�1n���:1����#OkԀ0"��=�<�<*zI�Zig�6S�׀�k�J���8ُZ6F�j�p������=?Jդԣ�6lMD~/�|"��tze��T�5��ŗ�	;�!��mXR��E.	���5A�AU�F����,_��c@]�����`y�%/����#Z��"y��=yG��΀�����=M���ĉ=
��ؼq�_e]�^����w6�U
��7�s�j�u�@����Nϲ�^�oG� Rl�l��7��?����m�VR���m�/,��DVRs~�	y�Թ;��'n���P�'�F�����y,��as��`��0��,���2�`����c��;p���P5'T�7�Q�[Q6G�4��]r�P����� b[��L�ƾdMzUe��4#@��T�r!�{#e����,��̟M�����_�t{ )R�~��S��y��w�u��O��'[[�Rf�� =�� ]6��wCp@�sX^�߰U_›�7�H��O�\\ ��PbX�Ƀأ ]}t�e�m����u�4��\ �����FVGY�z����_���g?�|������'?���2��.�Ҩ\�2�'�� >���l����2c���zn]�a�eDx�}fqa�Z�Xb�`!fd���l�倖S����������-����o�,�kl�}���<�F�Q%u���Y���r���d��*%!Λ�zGy��K'��f�;�YT !ZȮ$��Bv={o)�l��@�i��
\V���|ˊ��#h��~69��m���5�=�L�z�=���(0+�{tt4�����j�,�?���48��DlRa����7� p�zn��n����l��9� ��'���,��\'./�P��L�>������s/��<���N��^rey�{߻�����9t���q�g�yf�����
C6O�cn��������4�7�Q���&�Q��b��zN�s뀐�� �P���7wq�6�����?:�@N:���1�>s)���. WzƏ����.�oc"��e5^"U���O/�8��(�#�uiz�Ж��k����Q<2� e}�Jg)�`>�����?��?}���.;46V�(W
�����g���kK'����w� Zv?+����@��z.N��@�W�h<ۛ`�zdy�H�(_���I�*�-A ���|	���-JK���)>���"������7�n@-��:�+���h` x�#z'��;�X�(�+�]��� �3*���_� �@���|˼T�����bx�{�b�����_V���;� P?JI��=��|���|�C��o8*E���B�y�c��.Jz��f�g���K�u��}�6S{p�'���>jGw��] W�@%=�GW`��� ���K��Q6��n5F)���œ���U���>�e`D _cL���I-�����o�/2wt�Ts|��R����j��Q_��֓�ٽ��1r��;[�U�~�7k(�]빪\��qfh����9�Cܽ,�+l����fZ���~&�^�2����S����he�~W��&�
Ķ qF-�F�>���`P���-��-�VV[Y�xq�صz'IwC���B�7#Q�̆���"*!(k�~KJ�)m�|Wwܜ�Ph	T�� $Cp�{X��CehPT�����fP����7X�9�������G�:E��Ϗ��ˍōef���C��l?�яn~��Y1R��nR�W�g����-cg>|\����g6�x�s?�`E���#�W�#^ֳ�v;��zE�S�P� � `"�`�U�n�|�������|��>.�CX�޸PP��� �G��E�h���_��Jzk\������\?R���Q�ۺ�sT��<#U��]o�!o�?+�.�@�33����%�^�&u�g��Ok-�gt�I��/^��w)�yU�V�{��/��j���i�t��l�l�]��A�����>,�rx�[&nq�U�}l���xH-˖A�5��!��[�Vʀp�˻�]�Ʊ�VD��"_CY��T#� �A����󿟟���M�7��a����A�;?zT��HVZ�"��]��|���-�R��'fX��on�ӷ[�3�GO�\��WsU�3����'�� ����O&�0x(n� !�1�İ�����-��'��?��/��8�S��ϕ�8y���["��21���ŭA�s�v�;��e�>�q���� �{����Z������=S��^�em����}�!��δdֱ�:�Zx�^lǵ�y�9�W��^�q0U�f֯% ��g$�{ ��y�<��G(0B�#p��� �!�9�~ �uS��9~��7/�yq�<^�ȏE��K���3g/	pa��ll7�Bzβ/��w����t�e��������)���1Xl#X��-S`��Q�F�Xk�Ts`�(�J- "p+�|��w��s���ܪm�� �޻�>�mW^� ��{O���a���f��-<��=��������*� mʸ�@�pqE`�5>���W0|.��+�c���9�8�����\?�����/��X��F���\{?�j^�q'�"��֖�I���+]���30,�j�q^���^�h��5�{�uR��qZz�1m�	�]�� �u��Z�����3�Y�[���E�Y����˧�`�PD.�\��E��%��B���y������ϳ^�Z/@K#~��W/��em��d�"�� ��Iy�-��~-���*{��(U�6���o�w�>�:::ڼ��-��~��g�9uåc����C<$�[�(h���²�@#�kVe}���y/n�$-,���׃y���7̊�}G��G�R�\seEϭ�<��"�p���!
��5��	X�C=�>��|�)>��O_%R:����wfs�x-���?G��q�g �� �0@�Lծ=`�s��9�Z �g���f��j�VݗXG-���5���߅F�Z�m��w ��K�"�t�R��H�V�$ p9F�C@	��W��(F	��!�q;u+F\��L�;�ƿW��-ZX����q���c��p�bn�E�J�.r�89o�BTe�jo���C�ޭ���H��< ��,��o��7o��M��?���e���Ǜ�}�{�G!�����Ԫ�(eu���	�5s��� �J�%x�s(�~3.<��.��n �׿���fG,�^O�V��>�f@}�Rh�v[@呏[��K��[m�m�r1�(]�m�a���5�!>=pۓI��mT����CI6o�����dw6��da����jnX�&�R`z4ϞQЌj~�*ĕ�����uɀ�5��K��t�M��wV��\pk)N|��ʗ��:<;R�`3E#�A�D�H�pv���N��S ��K�{��>����H�n[?��|̭�p�1��"�淏woO� �-D��pE2��~K�-N�0��u(��.�^��{-��Q}��b�o�����G}t��J9�V6"
l�yO}+��׾���W����w���٥ãbx�8��٢h�YS_Ok�b�G��T��b���jK�;)P��؃��
���Cmɗ>�'��_����sЙӛןy�v��ڊ�ۑ���-�< b�����^
7G:��ۅܨ@��9�%_���3�"��V�����|��5Uy�ۯWc��8��//��>�"��(�,������y��ܥ�t ��J�T���&�D3�,2���k���VEn��ہQ5�Tڟ���<$���\�TF(�~�&`�[ji�h��8���R$a� �z�.�<�iM����rK�nXU�@Zl_����n�U��>�tK��_����R+��"�Yl�Pt�dS���d���?�������x���U���6��o~3[mp����m���p�;�Ry�(���du��;$��M3k�{�"&@l҄w�����n���K/n��P|�2@��L��\��;�%*���c(��-Δ]�NĔ��N@�9|��w'F/s�yyY��ob�hG{-�p�ےy��[m��Q�k)�Z𖥕][���\Gy��f䎦�,l�9�C�4�Μ����ϏM�����K7#o���4(� �(N�V1���R�J�Y���|Yڣ�g��S��x-��Fk}�D��k�9�B���c?)LD�\����[PI+���.�(�We�ˏ�C�7nh�y���3g��=�+��o�_)}�CK�JC�<6/���y8�w���W�>����+�y"^˄���|{�&��G>���������hs��_�C�������_�j�o}k�/}i����1�� V�������a�ٷ��fqT�y$��iz�^�Xu#<.:�f�]\6R���#�p���5F�B�~�o���|�8���������q���+�z��t�}�=���@�3"�;��"�kk�zK[�~���YE�w�lG~��?��fG��7U�E���+0U��$�침���nݏrƯ��
OdF��lK.i����<3M�O������G��ڵS,�(�f���m1H�1LO$�$ �>>7B��s���2�T6.���Ǉ-p"rPǇ�T��"h��5�]�Ľh���C�f�)n&��.h����u6�9p���,@8FM�44�u� �; p �B�MOl ��-Z,�Sn��8ǆ�m �S�Nqy(2�D�<i��ߠ��y޿3�����6��O�GGG�喈	���Em�)���>� ���O?�����͓O>9ӫ��$�4c��XƑy8���|�?�ab���(�(Bğ�K�RcNm�1��w�C6�n��w�`���$���&L,����Tʉ�A�)�J���8�/�I��F��߫�Ly�p���Q����6������ec�ۛ��W����i�v��.#�g2p;B���k�%kZ�+�7ւ�%�)�N����Ek���s�ٻU�#4��o��a^O�ʩl"�P9�OZ�ZC�P��~�N-&�<���i��w5��t�*	Y9c:1�
8.��ғ�͟�Z�(e���X�o&�h1�X�nl,#.)�"%ˉ���ᾎA��#)�:�:��m��4�/�"H=��Y�#p �X	��W���6E z�"}t]�r@$뮢�P/  W�8,�s(�	�\x��V(�w�CW6��"/ ��O��N���<�ҁ�<��pL�~BL�΄S��]D�f?��S3������`��@�փ��2���ߙ�3� `���,��)P��F���L<*���c�՘�|C���{��ˉ/������e�>7���m��}�ß�qN�6��G̳lp۶��st�S�o�c�um:}���~�ԶY|�X�Uv�(�r�g^y����~y.�
?�R�Q4"[{@q0� �=��>(��΋U^�l�V�.>�3�w,O�ww���V�W&��������T��;c�(LZ��Rf��Y
r�z��WV�]it��gz�C|��B��0�9�#�5��8J%,���de�7�Sn�F���� ������mٰ�b���[Kﱀy�M�m�}� pp0������F3ҡ>�����;/S�a��h�=6��-�c�:pre%��y������A���Ŷ}���?���C�'��.nU.��zWǫ�-�s���n���Ě�?&}�_���9(\>޾�Y�Zl����g�l.d(�]ʂ�O ��/�da�̢���M��Oh�Է��Ⱦ��R������/;+8�V�YaQ�˭¦&�8ѿS7l����|4&�G~p�wPL��6�V1�t���#�����m���w��%�//�w%�R5V�b���k�"r�9(∬�U���qN&ݸ���i��Lv��8Z �j�֠� �3X� �D��d�<S��i�:����TZ*�Ud+����n�wV�@,n�̃��W..9�zy�H���#B�T/0*!G��9�u ��{�dMY�,B��V-�?�?�oˆ���(M=#��M��O��*nu�%P|�e��P��}c X�pg�;�:�[`����BB� x�P뀪��F���}iO}x������p?����g�z1��1��]F&�h����������~���^��ԛ��B�'�QO�CM��.�hO%��s^�j�R�e�5���[��6�nՎ�N�𡯺�0 =� �a�̀qj�0�Oi1�����+ V_��l���_��EW�=Ǣ�ʫ��}��Uvn�W.�&m�.?������W�+�Xr�P̽�#�9�E#�w5�d|��Q���w�R�-y�+�>�r���dpl��3�ݓ�K���t�3�g��R`w�Y7F�`f��g������񹪞��L[��x�#<�t���B�#�qM������lgu�yY�w7c�a�A�r���^�[��PF�"�=T��<�`�� ���}_��W��Z��&/	a=����c��r �/�:��K�����M�,؀`o{|���i�T���$O��}� ?��C4q7��K�Z��\�7�sd �>��
��=��������7W��ڢ ���-�_�¼��x��W�Uo�?�l��O]R�(w�Y��yT����)˟��)[c�{񄿷���1�*�VIģ�[��hU�W7<=�$�עB�R5����8[g��� S�œ K���sj��vE�R�d�'~����韽�U�T?Z�0�|�N?�|+!制�s�W�d��dW�)V��^�[�;S�E����Rգ��J����l��c�[7֐f�
��.��ۢ��&�]8b���e�zޙ;���2��h"����C+q�gJ�!�mX�P�]*-{�w6c���&	�Ay��� ���S����g 6��"���o��+P*�+����^��퍷]�a</پ���,����qCE���"&���� �]�?�L@F�EPs���<z�@#�j��;}�H{X%��}�6}@:�e��U� 7���K����GGG��Q�U.�A?�O�<�_̖�/~񋛯|�+��������R���,��{�۬����xK������ǽ����(�@�e]�@����Ď���|8v7 !�DQɡއ(���(HJW|'�,�Uץ���͊�4�P� ��h\���(�����E����.>�R~rc����j�-P����)���꫹L�'^�7mY^��]d��5���^��֮�Y�{2���I�F��d
�.�t��H{���(��0kȉʌ��^~��{�2��ʷ�9��]o��J��TY��2
ܶ4�jB��*R62%���	��=		B@���6�k��}Zt~Ѓ���/���G�
���fS̔�S>�'!v�<�2	�ON���$�\��8V:6� <�0�8`��*��$@��a�C�+���=�[�B������	`jb���M�?qHLT�pm�?Y�ݭ��ƣ����;�˯\:v?�}|����a�#\�7����� Yn~�}��
�Mj���޻d���r��v��������	�
n8��́��~Q�2��U�u_�Z�g!��M^�o�<���ϟ��m FƢ�	���C�qMce�~�P�?T�~�����U�S>��W$�S{�̾���UwQU~�����_(��8�T3�T 9���������`�^QO��v��F�^��<4ȭd]K6Vej���]c��o/r��a����H����
��]*�����4]�֣&���Z+�]j�z��|cE0�1t�c�N=+PKa����/g"�%`$�,��V�)�|�ܺ��ݲ�W��+�nQ(q��,/�� ����)�S��==	��<��^ϟ��'����'�4_>N����ON�='�@��*��7PK��" �~�N@1��#�F������n�Gն*�^ Am*���ѼyK�	�|M[�8����R��K>���ō|[`k�g���z��e��2n�ӟ�ʾ��/��E�UuT�jW�����͇>����3��y����{������}��m7v�}E{�
�:Z�|>/D �n%��n�mk����� GqB�eB��<���ծZ��X�V�g�s�������[n��|z�	����~Jm?)b��6�'�5��Oymw�����*�i\�2��S��2�Gn�R��efu~��	��͊��۝zcvw`\��M��Lm�9@y�����|�d���`z�����9?*�zi�V�[4�Tm�jkO��+���
�ge�pI���ّ>_pE>P"����*����:c�ac:Uc� �����.iU}���~��V�W�����י��H#�Գ�ca6[��*���v�>����&���4V�i��+K�Xe�0�����'AvvJ��{��'6����_���>;��O`���K�*i����d	U�5	t ,>��P&�#�U}pwP~�5K�]���T�eɔ��>z�����B�kXh��G��|X���w�xT�ܕ�7T�&p(p��d_���gp�6�v�M�`��X���?�F���ѧ6�N���x�W!�#)J�q?#-��>��[o�u{: �Ҁ�o)c���Q ��M�)`G�/�x����}�ݧw���9?���R���V}����v��ON���?�2��S��4���c���H���;����E�&�ҌR꼌�v�/Xm!~� ���	���N� �Y�q�oKʲrH�=R�i�J�Fj���(�����$��h����%�LL[��4Q�*���!�^�vxL'>�1ھ(�K���Q�J��z��q+�H�F�>�>d�P���qn}�ޗ@e�A�2�o��,� )B� r�����������LB�	j{t���Ϡ�g?��gdݝ�~iO���uN��l��]A���t�Y������u?\ڈM_l�Ȋ��S=�O!`H56Z[жeB�����;��zy �����7 �h�ĲF���L>�rM�a?�я�r�c���e��O�����r�-�+L\r� .�p��8���n��XW�_N�	�=���_#���V�R&�k��ŕC�K���I�����
�x��V���q6���S�>3�k�q&�����g�y�/~|*۬\
\��8��"�:�7<�g�WƢ��5
~�Q�Mnj���v����LZ�7�$ ̌2���-#�0lɶ*�J>�)c����7��SD\�]ۅ�-�=���0��cyF���K��^F����+�~Rǒ|Gx���a���]R���t#�w� p� �r��iȭQ P���r7~�Xl�,@������N�>�7���$xg��I��,p��t���?��l՝������c)0����'#)�o�_X�� �[� �"�	@��4ܯaMĹ 
���[����;�w�d�q��_�J�h	�?��O�'����[�g�����pr/_j/��(p ���ӈ�|�TI�]9�(~En)��^��q��UQ@S�l$dl�S��+(�G�A�uEYU��&�� ��ec�ĳOL�������@�^ǙӃ>8����zJ�0���T��kW�@�{�Js�p�`<��OJ�0�]�_s�څ��o���xQE[��yk(�k��}[[[8!�q�ei��EU����xų��R2��~g���Be�w?�D��V��1c���~|�]Im����#\��$��WZ���[ G���!&�C��Ճ0T{�3u}��%�2p�����m�ԦI�|�mo{���9!���/����=�ܧ��=*����0��`�W<,H�����/@�7� 4iG6� p�J��wU�=ژ]���E�e+��6Gq�"���6��+�����x��Z�V�՞Xoe�S�b��y���|��|F�(�b���7nP76;Ÿ��=���n�u76B�%A���,S�#Ȃ����Mt�y�䦋�>���K����u�mTj����a��E�\���W�{���)��WF��{���''`��)��Oyb��t]�8g}hC���şU�M��0D���g��D�B�s�5���7���e��C�(@m���	�%mx���`�2�q�Ȼ*��գ�]�*F�Uk#���#��=���w#ȯ(vv6��}3z��!4�JA��G�٢J!��>����*�e��x����)� �������'5����|�$l o��O�����O��NB�7W�& ��Z>5���>1	�ٚ+ #�/2 �ef�BRϱ��}�~���Nx�/�&��n��ӽ�n��/)���(�#py�����j��D@���[� ��W�U�ZYlL@W�0�tS,�z_���t_�u���%�|��m�F�^v����%mw��l���wg�4~�����������[����c�Ϩ�o`D�xS�jw]?�OL�ͮS���u:^�yb��L���4o|bj�sj[)���r���-�M��Ӧ�Y����*8>;��\-Z��ke[�n��ׂ)�7#�j�̊���)����O�2��g6+ə��i4�g~	���E���;����GX�Gi4��钶�Cܴ�)g+��s�r�{|�sê�Ѡ~��[�<�k�?K���X�0\?���f��6�z�O��[��S��G��VN�&�;�	|f�||��'���g����Ur�:��J0�	L�]��A�����1&0a� >,WK�AGy<��Û������{������t9|��t�'�$ $�*I���R�2*��������х���lz�2���������M`5q�������I�`�����MN��z Xe��V�V<�2*����;>��=�=#>�R��6}�Ֆ�������x�-�1��ɩ->��C]�&b�d��b��^����Tߩ.n�wW*Ѽztf⃩�8�+B�����E_mj
�(;98�hW��u'I��f)�ʼO���>,��|�ꃑ�V y�Vܬ�{���k^Uz��{4�J��WG����L�K� ��w3�u%Z�[��,�U�c��I�*c$M����h ��	��/;`q@��N�E|QYDzd�өWw�}���0~�j �NǛl���׾v~*ߧ��xT'n	�(|�����p�r+˞4�Vp,��zV ��r+-B�*���/p���
8��ɑ���1Sټ�|�������K@Y߀;?}L�)p��o���◿�-��	��<�g�nH8�E!��Ei��^���]V\���;�������~�oS VuP�e閛��@m���8Ɋ��E�Mo��� 6�`ssѲ��U�����6�]�h�ait+���+�s�$��n�|���K�Xn�
�7�ѓӳ�]-��i�O>��ӏM�5��BB�?*��+�h����q�����eYQt�� .�_?I����~��>��e+(�.�Ce�#�Jk6�T�R�f����(��fŊd�f��Eke�=&�:a��E�d��h2FZ[�H�?vUb[�H�9��#�©e�*�Z��m���%�B���XJ�'��< ���w��؇?��N�B���|�g���������n>&Рv�0�z	�t.�,��@pT(��pG85]S��WHG���ʠo|TU@2�W����}Yʕ�,���
⧩��]y�.�b%pD1H���G�YB�v����:�@�p\l�RyU6�ᳪ2�?e��Z��o<60�d������=�e}�u��2�tvy�f�W7ۣ�U wE��GuS�p�ㄥr��Z_)A���­�*cw�������S�����?O�����v�=���O~�������S�>*�ꍲ���"?Qq歩�u����j��+>��G;��?Eq�t����7"_Z�dr/{��#���V���H]G�XѾ��U:���
+e���������b�1�c��X�5��l���0�������K��L��5��U�N/�I�<�]�ͤ��A|��^�W�������YH����7@�/�	
�"~��:�-a�\��b������=���}�;ߙ���%z6���Xuk-���Q%����g 	�P���@`�#B�P����}*�#.XA�� �$4]�F@���O�rq��H�}�Ve���n]S����!�# Ky�� �v���_��� -���fQ��[u�u�K$�Y����G�s+_V�jlB]W_ࣺ�P�f2@..�MX�ٺ.�����������G�����~���L�&ӟ��?�?P
D���EK���%?d����!=� W|$^�������T�:������#-���[�*�Q �oڥ���wɿ�Czu[�簋J�
��61
$+�_��|��o�@��Ycu��.)��P�=��ץ���_B�~N���x�"He�%��.�.|�X�g��E���'�w�������:�6����q��oՕ�H9��}�?\>�O�w��$������H�z�����L	{�	`,������*����$���_RB���X��J���e�LfV!�ǚ�Ue�; q���$�)Gв�>�(]h�����X�X��X~��r�Ip�������r|��e ��>"R_+m�Ҽ�-o�"���"m���W�*w���x�n����$�T�ˢ$����@��Q�lE�ώr���Q:"��,���g��o����?ӒEkereE����֤]M;m2kQq�g���VyWe%<#Ly���e𲍖�&�%TҞ0̀��w�x�H�#�]`����=�f$-%K�N�<&���5FGGGO|�{�{|��|ԯ���,�
�
L�B(�����Y�_���-`�������<
�(SHȞ˻"@����Ve����#����7U:U�5^}l�*�\; $l�Ǧ�<u_��<��&��M[z� *��=U�(�(��-�kԋV�r�>J�xr��'�1wM��~��O~�;�Q��sJ�Q���6c�1^p	�3�O������r�q�3E����w���o���.W���w��O�ӡ�"�L�\�tȲ��l��2��!)Z2 �+��ʖF�O-����rd@�Z�����M���n��3X� �k�!�v
�<q�m�}j�ל��&����.������o|�[w�9���Ϯ S�@���i~��TN��7ƈ^���V {�0x��E`�S���f9��Cj��'��Wb>� f����ǵ�p���Q���M����I{���6X:N������p`n�$E���n�i>�Ń6�-!w��ӵO]��� �g�6��;��G�ݿ,�ګ�^����*��P#�9��S��(k܇w��dde��h)�mɂ���n-�ɝ�u{_2��V��F~-���eYC'p�wo��>�e��Y~�rf��ך�����Z�-�If�Z'��I*����į$P9+A���>}?~-�[����?}�o}맧�?�HrWP��%C W�\-�Ǔ%u	Y� �O�9�U #�q0F�BW!l��9h�1�8`u�Q�W�w�G��O����*Ś|�o�sKuL#��&��ڒT���Rp��� ��5�Q"�!���]��]Yn�t<����W�>����H�>������k�d��SO=��7����{�s��ͯ������$�+z�O��L��>�<����侻Q��d[+ݨH����ywpFY��^�`�$��[�^��0aU��Pֳ F��݋�(�8�[u����Jd�W����	��>�}�=��3�_�R�gGp�,�;_��Ҕs�O����u@��sϓ�>��cw�}������Q� �p��1V��+n�%�~�,�z;�'��lC�����A[K�9�>�e�I#Oǹ!{~	Ea��#.k��hF����j���o� �W:nJ��/b3�Â/T�{�WJ���k:��g�y�u��9��&W�s��|�H�����W|c�ƫ���(�Şev�s(���K҈���Ʊ�����Z���Ja��j�� �I�,g�8�f�'2_��-�E�VX#�x�U��s��	櫕��l=���侖~ʕ��F3Dv\�����Y�7�|����kڢ�ttt�䗿��Ǧ����f��#(˭��BM�K��%P��\�����	��q]�J� �\wnᄲ��󃧟�b6��X�*�:>��o+��*�S���=�]��'�A���� ���~���#f��O.2>~���_��A��v�N;�۩^��+b���j;)���u����~;�m��>����rD6���鈼\J2�╯Q����%;ZmS�������/W�d.�+�W6'�j��7UK	�s��[	���'�L�]��ݯBO���$�b��zfi[���=k>B�pE�w���	U��Ã��}9�W��%4�4�_O�R���M�>��� h����܅ ��/!m�d ��_��������f|�~�-E��j�3�C���sE��d���<�y���~H�h��={�[{���q�� ��7n�%|� ��&(�4.��-����Oh�d37������	槼�&��R�C;^~e�/���U;f����G�O*���A�[��*3��s���ʖ�����U^�s�8ه����ex�ٞLΞ�'��� �P�@mi#d�O/��[�ү��bG�J�ܞf�ܭ�Q&�t�֩� ���"��^� ���`JD�&B/̟��au�A���:��z�6�)j�`C��O�\N/(!�*K�j{6�Xj��",vQ�:eքJ��x2���ّk-ǽ4F�� W>⽞�7��0^����8qk��+r���	Q
�|V'E�Sozӛ�;e�����/|��:�Sg��Q
����-�>�"���j�œb��
�83>��EټĚWɑ�߻�]ݫ�RK�]��������~�Y��BsQ8T�N�DQ{��b���R��֠n��?�w�)2���CfZz�w�Z�L���t1��d�,����U�����ON��\�4���TǏM�����U{�X�޺���H�!`�<�ul����f��pD .�K]�~���ҶK�#����\)�#e��Q�E�*��y?�� E�b���Q�"�r����n�	ܞU}�R¡1A$Z���R0�p�1��ZI�l�'�ܺ�xUV�����<Z���+m`����'#8&{fi��h5�a��YK�,�#�|�J��'ۑZ�Z`Մ��W�W�5�� �X��/�;@�B��$L���>;������\�$��7����w�u�9Yp9�UV] ����w���?���*�7����=���[E>o)w�߻Ү�}S5�窹%�,�5����ԟ��� ����nЙ�7\ڐ�4��r�w�;	�����Oc�co|����m<֘1C�� q��\��a�ˀ�E��H�Z�Ѩ�d���EZ��Ż�wv�k�E!����<�Z��O��57�`�j��K�RZ��Ȓ�2bm@%6';��6�S��x�"�jv��_�N�����>׭{t��U�	dp,~���2�����K��-���Y^��
�û��姚X�L���ӵHq5�kq���T�G�� =���Z����\�G�n��E������]#4�Y��%Vn�;C�1p����U`/ZnE�W}d�e�(���֑�L(�������H#��R��E�,��M�� �Q �2 ����ZY��M���Ȳ	kW��R���Zf��(N!#}��bqb���#��ݔ!�w$h�]NO�^�BW$�׽�u���˛�`�Xhi����X�b����tE1�,�Xd����e�3�������h�Gn�g&x\i��콸J�2Cy�����^xyy��g��6�N�����u�
M@�'�q|5'��s��`"���V�\�UMQ+�y1W�r-hY�����'ߝz��ʭ���ai۷��5p{�k1�}��(���v��U�����Ea͠m�}1cLs	e��x��o+T_��ݽ=�)YEgN]Xp] +|�����w����uN����o{��=	�s������]��76.�b��}6�!�Y��pn�֡�����^ɥ�
�x��S͢�q�+�,G��߻o0��,�䭿�p'�qB���ic��R�D;NQ$����sn@�u���l�n��Sɹ*�Q�|��<jէ��#Ϯ-Kk�8�y$�QŢ�����z]� wW�V@�X�w|_Բ:F�' [32Y��h�A0b�k�u?�P%!�G������H��W/�D���t.O\/;��C=��?��?���Nc="\����a�:c��eiO�ͣ1���+->u`�dD��.t�V�L�v ۲����rE��'����L�ʼ4~��e'�y�i�1	��w����������L�&ƚVK����ƙ�N*�GnRR�}
E�r�h�̂���*y֢�`gɳ����H�#�?�r=R���:�k��w��
p[������V��	(��iU������+�pe%���ꛖ��G�V?��g�V�[��X�<�&��,��mt��e~G�N�p�ps��ꥐFXR�z�-��?::��-JN��=��PJ�*�ڃ6�v���{�ѷ,�
�����ƣ.�튧S�|�C�Q�`���}�E��+ ���Q��y|���>��PLp�0^�@��?l�X�l>.�T�3��W���� M�v���~M�5m���׿�h�~�_ly���~X}��YC�cQG�r�F)}'Z]�g�L��Ҳ-�=�N5�:�k����rX�b�d��]ho 7��]@nf���vr4=�O�(���٧F;�^�z����I$�=r�Lo������ad����^�!txV�חH��q�rX���ew����ToB{i���6j/�}��3W��܇��.��v��;�Eq�
�����(��d����3��S�R�>��� �8�)�Dh/�>��N��h��߀0}��>T_�[ ��ȸ���}#!���MS��J^Sc�o|�)��7q�`5ʕE����l�Q5wG��㽥��Q�Ԓ1K�9I�Y[Gd�.sC�x�$h)��*w)�� nf��'��U:�*M�eE���������� �(��gG�z뙪�#�<ӆפA��9���K/�4��$�ٹ�p���4	��n܆>���B��J�}%�o���c�-��%1��7��\��
��XE~�ke�u:�p8������7���no��֙�����]os� ���Mdƈ+(�/)3�. �% ُ�u��79�Z!�@}!�|��g�C��J�
��!iɩ̲ےW��Q9Y��ӻ���O�i�^��9��,g�%����4[xg�s��-���}��!_u�dˢ�2B#�\�F4�����s`d��kY~ZFA{�,��/K�,K���t�- ���7g�Ej~v�/�y�5pu��,�+��jK�Ǭn�"A(1]����nn�c���Hn�+��م�w  �3���ա�}`��z�6��������t�X� b�7���?(
[���p��|g�������[o��Qz
�G�g%���,Z�I��p'�+����{�����y��C�D�*�~�"��lu,���ZV�h��:��]��}��^;�TK�k�F=��>0�j�۲�e�Gޏ�i�˖��]��;�Qp۳L��lR���J��[<֓�}R��"�fgy�=?�A��(�ث������
��^wSS��	L���ͩUjO,��*�%���.x\Y�o�������\��S����f?]��H-���894�l}̏�4��utt4[���{6w�y�oP��{�+u"���K��_�s�=�=�N�r���; �͝� �[��1ϯR8��}?6�<Ǹḇ2���?�L+"v.���Y#F��10�DV�F#Ȩ��$,�# ���X��^������}έN;YpG���ߣ�>��"��/[z',a6�N��zV�����&�}�y�pm�[�q���u�[�|�����9,�V�/a �C|S �v}����|��>��[޲���{gP�%u�%�_���d��u̩@������/�>�Y�1�,͑	x	�od��W�	�
�>��#��~x�r1�� �����&5��U����?����}�����#  p�\�7�Q
_��
^t���?�����O�:=G,����E�s9�M�(0�|�x�]��{ԒW������Ѽw�����- =ʏ% ����� �H�vMup�Գ�TT	ܥ�j{��}�ƒۛ ֖��}$(|y+�S�<�y=�}l(���$Hu_`���l�{��aX��� �ZB�;ޱy��߽�뮻� Z�������i)�G?���~����`�C���=�-лJ��D����6>���]�z׬8�t�l����g��~�8���-���N|%Ғ,Z����FrCd#�~���4�?%@.sA����DY�,ɲ��$��٢(��<��[|v���g֬MJzkca�5���Ӈ�����������Dѯ�]	�Ty�l�rk�/����z��C�fܺ����>p�i?���ȳ&�Xy[`z�ڇ�z,��3s�'����rj�_��C��ru1���Yc�͛����S�� H���=�L��������l���D�}��z'"�-�K'���t�P������@�����B}܈%g�����j;YD}c fN�?�,�pu]�X��=A WK�:r̯���qT2�wXxk>��+�]���,�D����]Ej	�oT����(毾������ߟ�ԧǏ�.'�l�-�a����7ˆ0Yp�OEpQ��Ic���3>{������x��Ǖ��}����-�ܲ�(B���IƏ�{�ʿ�p4�VSye�2ů�KV}�Z��������r��s訌i�����B����?�42����������;e���?��Y�1/���U�z��.=�!Z��qr� ��P<��y.{���Hƒ롱{�Cc��ヶ��ǁ�B��'������������U K+�]mZc�iI]V[���Q.�@i#ԯ*��~W�
ܺ{cI>��ԛ��dc(*X�hj^�����u@�����j�{��'�X��'�0�xt+�ܥD����a�V���N�lI|Tzn��K���ן�z�2�q�4>.4����������_t�F)
/]��H\<�>�"﷊�<h���H�2�����U�g��|�z�2��k�鑧��cT��۶[���ڠ��6Xg�'��X3�^hM+H�������s�3{&�������ίO�#j��h����0��ӯ�~��'**��+Y�<|	G��9��`���X�����c"ڕei �����?O}���}e�8;y��h}�s�.����{��'Y�� � 7���1�=�hJ�GF�	���shJןƴ��~xtMP�0*vl�v ��X;~�����nXn�3
�(q_],�z�㜩�o(��( |�H�N�S|hh�sC��X1ٴͱ[��SIq�/"��b�G�:�V<ب%�|��b���T��_��64W���P�%w
�����&�M������=�^E��E �>�ĩrz4��/��O��6���x:ϳ���Z�b�s��S���Y����߲S�DSm����|b�<���S����q��w�cY�8���V'��f26�	|	�:��b��P�7Ϸ/�gn��lO���zN&�%�Ǻ�����|�	���r�P{�A
�>�ƕ���#��~惖�}3&ώ@�����~�Ґ>�D��r���>N4���㘿r���X͐B�p��`���{�op�ts�@���q�7���~/!�sV����������d�T�S�Z��*��n��%4�V�Z�(���Z�搿gvR�Y^�V[�z@����Li�-��e����fֶV^"��2�"��J?��B�D,.4ʀ[B|�F�%V^�V�e���5�:�	����5���x�: �T�Hܪ�E�vjY�Ƙ���[�c[ʬ]j7�Q���6�9 ��r_[����Ga���x���4�{���x-f+a���;��y�Ń;�s �+����wW��{�s���eC����Pk��/��ͱzV�.3b�7����U�m�l�^�2�fo_�a�jYZ{��P�Go�l�w�ne����iicgV�L�[�����K c��F U��6��ضm��Pi�-�a�����ʒ�%������n��7��c�ɏaMEhr���E�%x9�W�3�%RB/&w��ۗ��{�w�^����������˿��X���2�\�o���^��rT0��"��R����<��T�,}������6��q����@>���e�,w��#8RZ�]����r�!�E�2�8��G���so��ַO�:���G�%b����9�� ~x����.J�+*���&��)Oe�i42_Q�lzY������5-|�K�Wo���S�G�V
J�K�Ɗh��B̸ň���:����,���V}��8�޳�_l�%m��N�Re�����2�a
��>K�Vl�p-@(*�'��X`��>VV%��a�d�#Ĕ������E��g�a�<�,��W�����P[��K#Ap0��㨒���at�y��)u�z<��w<{��2���2�B^�	��V�	�'��Lc��*Vo�W^ye�Qa?
��W�^V^,����DX168�Lʠ��7��������G�~���sí�<��Z��a�TN�s�#&�H2�3�U>��d+O�8�4e�ˌYY���S@��� ��_vZ��r�1+�O�ȓ����S�Z@�UO�C깝o2[JSڋ�J�T�UYcg�vv6�3ZY\���d��gjP�w^KY�ʩ��,N��7�d�����_6d�E�%=�cajn��7��=�;��;�|��{���]h�W�,a��2����� rƔ}!w$���/��g�����n:����#����P�-��,�����3�>ܯ7�4V�;�	�q��MY�<z��W�q���<`�V�(��������7ëvwr����B���=�L(K����1TY�<�d/���O.�B����q��=����=r�OD���2��kY�9���:J�p��n�Ϟ��s�p�(lcXt��f�ZZ����ߴ w�,(�A���7
���,�)�c��9Z_�ߖz���g�&�1��Q�t@q�������)C����^C]|���2*+���"��Y�� ��P Lqo��b�����.\�����/��Ty�����d.?��7���0����SDQ��.���E�]�W�^�?^vk�>�1�R{�]�����}��_�����Q�%���/��X��4m��G� 
�D�ƺK��/7?�w��X����7�9�Dr8��~��3�����7��� ��UU�rP���|]��A!>.�6�̥(S+��\@����s�/=u�C7���3�b��ZִF���Υ��r��NOY����9��&H���ʯڶ7������*+
�8�+p�Ub��N�0]׷o`����(����q�����&c�""$6��DX��"��q���/mN�����k HVDŭł��f���1�l�WB`n������կ~uL#T�=���V�<˄y�CG?_�:Ơu�JY���{�����E~XǾ����
��������?<����@ߚ��jQT<��ǌ���-����=�XN�'Q 4'�J1�@��'O���*����/�_}��sZ�P[��嚀;�ĞfѾn����n�W<�p	�\m���O��s�AU�P�ʷ�쪬%���.S��2�d��/��K<򼣦��e��� n��>�-�[���4�V���:DA���z5�� ��ߖ*���|<��O�9�8P�� ��O�@,U,{c�8�YN 6<��qS@�%-g+>�� A�0U;��̭߇,6{�V�/@?Pb�� ����[�Va�b	7�B[�UWņ%j����?!�ܥ�쀾n�{���b���R���2�Y�|��\:ju`��8Xm�x�>w��t�~���_Y�q��kl�ˇw��x�}WRf��/}i��G�>�+&����_�98��5�F�/Yw��ϻ��n�F|�k���G~Mݟ2��ȣJylɡJ^m�\��IW�ͩ�zA��<b]b>q>z�W�F�܌�����S�h�KS@r)���;<�8Q���g�k��Ι�ST��fB�m�r	���	�;⫱C:?:`��vX��XL_'6��� է>�����^xa���^OV��h"`1,m�m�8��?[��5_z�X�V�l�bӓ�NEX�ʏ(Js�̙�B�ūp����Tp����Iyd!�b�&$�� ��G��.^^�����G����ɘ�'���k,��z �
�SU��7޸$q�g�7� "�Y�[�V���5�*�	w\DD�����p?�m)*6�R�Z
c+�x}[P֪s�v���\ڦ����"x��8�g�ၣ�=�?��^P���wʂ�6 �����NQ�k����){�9�y�:���)��]lw�Xj�?3�
�T��'=��""!! !�A�|�7�`��?��O���	������#WEqy��Giqw1. ���%9��9��"PL�G�2Y{���^�\�q1hYp���u�^�G����S�s�I1T��ek�6/�#'8�� ��ٻ�T
 Zp�e�w�>.B^7?���U��r����AI�HZq��u���?'q�DӮ�[R�p��e�~c�����v� W��-1v���1V�̈Qs֦(�O�o�N)�Y�����H��]���j�j�J	pP�NnՁ-��Kk4����NYi���걎O�6�ps(�gM��V\/3��Oh�8X�K�]�"�r�������ꫯ����?L~��j��1-�A롶�s���������KP��#��V�" K�*����z���9w{Q�D��{|�ޘ6֗H ę���h�����!Ǳ?e���G�+�_;
���{�y(���%����K/i#�c��S�<��G��]n	���VI\�eYo�W��C�
<ʍ�Cdl��(wQi��G�Ĺ��b>Y2ٱ+ �>^��9�W�2�g{뷔�w�׏��P��0�^Gj�݅�rIGLYZ��[b���ԩ�"�W̴*BKo��	�$�5����C���b�u���)k���=7�'����� ���)��&�i<��Ab����$2���M3���D�'-(�����C������v��YH���U�xg��/9�"s�4�,{� ��
�}�����o����ߪo��<Z 7� ?�~��(,����Z�%���:����O�S���v�m)+��F�muVVj6��DE��T8�%�݂�@�r�������(˲y���KK�e��2�w&�צ�9�c%��Tm����q)U��|�F��
{L����q�N nl���W�n���K�湥 -�g�f7EѲ�-��Y���Vaʍ��C���G�CB�FX6�x tƚ�8�)}K`��Ah�@�7O�>��������>���?�8������,H,�Fh�Q��e_�}9N�8��nY ?�о����H �K��q�WV���c���̲X�������(��[?��)�pm����*�S�d5Լ���5+�?ļR�Д��J�C��qY�S^��E"@(k,�}�ݏ���+O<���z����9AV�/p�a�`�fo ��F�x�sHD{+����?�j�E��Q�2�kL?e�1[U����a+K7e,Y"�DS�|3�3�*�L���OF�֣��͌�gI�3n�&:����0�����3`}2�Xk��ce���tkO�l�� xU���X����W�IM�/B"߭~�L�D�XL�vv k)�� H���[���oϾ���p}��ǋ��Np�����eh6��J�
Lys,-1C��Jy���E~�4~*r@��V � 7�ԘGE^>��-��s��]��X^Yn��t��������}����9P}#�R��k찹�~�z+�ID���k*CV\�G����?�Ϝ��7?���}����N�ŘǴڂ�Q�%�Õ4�|��[������u�:8b������ϔr�)���^9?��mi���,�S���V@�����sh���.�
��t��c����@�&����s��">^��ճ����@��v���S�)��1��sʩ���W6�"�径���B*��2,H��"nYs�M�%4d��cO?�����z��h ?�����ge�hX������AcM��vP}�/$�%�xtM��b��ʚ���^xa<�@y
,����9���"�^��1��#n2so������[��<���4^������תvT��!�;g<�I}����"�CsL�MV\|EU��W��.nMw�Q�P{	����?T���������<; ��4�œ�_ʀŕH#�K|��Z�th3���ꀖ�lE^���S[�����Y3�S|n��+[4��f�Wu�s�R�[F�^��u�����k�]��~o��˨U�� 7N�,��U~)�ݦ�{������o]��+�)�x�y�ٗ�{Ax��G�f���o�PD$heQ��թXX� �9��A��BH�X������Cޏ�w�}j���Ϟղ���??��(����c���v�ǐS1Ě�W[a� ��;�3�,�T��� j�����?�S$+���3~Dm<�4���|�EK�#���4NZ��;���z}�c��Jq�ڍ�jo�A���_"��=<*�w�+~�z���˿c�6�� �� ^�\�ʤ:��R^DR&5&����p��_��W?t�m�[r�9��������F���������xl͇ҥt ^ͭ���w�/�L5���d�T�2��i2�����B��-�&S�׃=*���1��E�O�o�2��=�����Ҵ�l,n�P�S�Ş0-��6����Kʎ̠g����@{���5򯔚he�m���1�0y�@����=�����]� �Z)����z擟����������?����C'tE����yYo�|���� 8��.��u��c��-���-�F�+�� a,˭⵪�d]����ە�&������@�>8�h  ���.�A�����pN�O&d=�@���������d4%�	!&˭�Ms�e�4G`�Q�̨�D��-K%�ȡ�?^\�,��4_�63�?�s~ ���@�k��vv���笔4���/:8@f3_D1~1�Y�.D�@�@����*��s ���ͳ<��?.-�(����i���z6�����sճ7�2���N��uA��λ��h�Vߩ��ޯ��4�%��C61"�u����&�6J� f/A @����~o,�� ���ђ7zx�R���+�Ґ����뭷?u�ԇF�����o~k �g���eF��#8��e�U�%��H���?�<Z"ԉ�vģU�+���B�siF��W�,EE��tz���/�n���w_UOyX<*���2 v^�Ȉ.�=np<��Az�	-�QKA%N���NPۆ�7n
jo|�	aŒ�����d��-��sP�Q��uFV܁���?��s��+_����0�
�@�N�S��V�DX����,�1GO��i�;n�c�K�z�q�S�W�,�-��4'����7�� �(w+j�Χb~sdpV�m��\p����a�� s��Ziͻ�^Kn����?>�	�X��M3�\i�=�����w��;y��迉k(��m�o:����eU,��Wֱ�����
��>}����"&���$�ֶ9Qi[�\��߾���vh3�]���Ը?�H��NB��D�pH8\������TT��=p�p��@<�/,��}�j<G����^�����Z ׏��/<��-14��iN�O���(+�Ɠ���Ͱ��5�_�MyC�G�(nRĆ�8;�����ǿ���ݴ���[s_e�YB�hWnD�%��Ǚ�s�C���c۾wM���s,�1����zڥciW�Ă����l߅���"S)��3�/3�mK�����d��=`�Ѝ�.W������d��|qEp�����j�8Ӆ�K0J �[�eO����JO�� +�a}�3Gi�GK� ����{oZ�+z���p�� �I��dM�������rk��-N�����&�#`�6UK�_�"@%���}l��:�¸N���c�<�KM�ĺ%�8�{ĴSs��"�!�p�,=�L�a�+cG�5�de��_��J�ٱ.�
It�P:=��W���
���wu��3g������ɡܛ�8_�۷�~��P_m,�I�y�w�\ �j,z���)�p�.�#�]��hq<�!;1/3B,��a"Z������T���)Yk������z��ߖ����2Z��&,�z��l�`�- ���/72��e� z̳Z������c����v*�m�
������#P8�9�$�	�k��!�Mm�}���s�-�MG��B& �����\���DU ��,� ��_�\ E���-᫶R?�2=yG��9�� �~:��0�/D~^6 ;��[a{������Ik^ �}c\l_�_�<�@*���V����/~qwD�9�{}�F6V4F5f�y���?�����o(��|��Ϲ��c�ѡ>��0Zn�3zgN*���K���fTPn���u���9�vC�<��rH����U�����p��ڮ����]Ҕ�ڦ=z �\^�)(kP�x�SǞ4[�	���X6��UG5ŉ]1���V&�$��������㵞���fV���U;W��@�b�fa%"܎,Xq���0f�@�Y����&�hg����||j7\�:���+g r^��{���UVQ�	`-1�B���K��k	j��ѿ�O���V`�L�\�K�\�c8S�|����;˩s�I�.�)�ٮ�
����Q�6 7"S��ҁS����z8�__s=���Yml{��Ʊ"��q�4�,���|�{�N��զ�������?��?Ț{C�����y��?���0������fU�CP�������D�G��o��F�_q�!B��h���T��^��s�"�XLc�Zsl)XݵLπcK/�7�_�镳�����Q���/g;=�a��z:�j�^1w�W�̣�ڶ�92UVg�[�~=T�9Lx*]O�=�6���4HHH�&~,->,)�=�Z"�Phs�M	� �9;���{�o��on
�;�e����L�$@��N��;_���f9�-A*�����c���Ƭ�+_�Yo��ڔ�{ns��t����	k�G<�m6~]�t7	_n���]f�,a��R�3��˞���峛�y���q��]QdMȓ�����q���|n�8m�G���7��4n���������x��w�������������[�i ���"��}i� kc�������~1�4s���n"�#�	��0}��a5ֲ�e��=eD�33�T4�1��6j��M]���UeT�V}*~�����)�^��qi�G-*As-�kPV�������9�S̡����An��m#��r��IpH�jS��ӧG��Ě��D�����B��a���<�]��;��ֳ�>�� ��:s�����~�?��G_~���
��%UV%}lea�hP����@+K�1�+m� \�N9��LY��;�]��6��2�����w�R��{żQ�y9U}�]�έ�w!�{���X�-;)O{ \S�_'*=�*��3߬(�=5G��1$�I�R>����7�z���{b(k��'����ǝͻ���:����.�^x�֊��Uc^ _m��#Щ���Ŋvf~៌��iJ�ux��y��W[F7���̌(-�V2zh	�nɈ��Y5������Q\��SU�0��[v�sz��jU���a�K�Tp���R>��ΩG�"<ea�L/�Ke�= 5�fQ��W��GC\���eM�@���+��� �,�-� C�� �':��@�z6 �'~��a���K~�����!e=�@�$TW�"�O ����o�����M]\W^jO���\m���'da�2�̍&g��^�}WuYC ����;'_�P%�@,���d���T;�'��HVH q"W���,�s���)�m�C(�� ,�U�p���y�'��<��#��6��m��ŋ���0��5�	�&p�����{F����_ܜ.ƻy�~�7�_(�Nσ��9�FsK�G�Ȍ:S�)��)COf�X�*��+ۖUድ��eq�;UX'ޫʭ�q���/�xl�i��̖<ۺ׫�m[~Kc�u9jP�u^�&
�֠��͹_������ky]���K�%�e]=p#��/��O���{	؞ӝ$^'� �I���������K/��� �����>�:���� ���W��<�+�='p+� �,�X�6n���]�|����8�l � ��_z��,�ĥoBI���M�: �Y�-�ȝ�(�Y����&O��͚�k�5)MR�4�4�4�r�oYr����Y���R�4_8���1
�Q9�R��U�ƚ>r�8s�����ؿ��>1��c�0�ux�7�|i����������p��g�=7�m_J�,�DfQ] ��'���־1�Ց�n��Li��e�?���x�=�V��s��1rB��[J��&�o��h��f�Ve�Es�-��5|��G�m���WTu�a.
U s��d�zM⻤
���X�"�ka�CkM�X�9
NOY;�f��^�K�-iJ@����A��}�fY��y������C�����[��e���'>�?��`>������ݟ��׾�5�}��7e%~t(�A��K B��cr9���n�\��nUUZ6pLV[	m���7pZ��׻�=A��شXa��JSJ�Q�`W0+�/*�\�V����-����V���--���y���8hб>��HD,t�#���"�+J#�
��Gi�[�+n�n���e|��a(���?��a\��i(�ʠ�.)�����5��֢���Q�Fu���<&4��<V1s����៬g�o�mWY"�,��ukIx_��lLU�e���~�}���Ꙭ>G�nj���H7���R�e��>����٦>^�׫o�]Q����ے6��H/�)A�s�Ų����;�����&~:exX1}����|j��B��4!a$a8�Q� ����O�;�B���Uu��7�!��GA,��,d�*Ku#$������C�W|Uw�]�u�>��6��/m .m�|�|�շ�'�-����ע��]�8z6wf�#Kۣ��|���=|ƣ4�!���*� �PO�7Yw�piÙ��<h\a��oV	P$)��cT~�zN`S�*����R�TG]W��a.�;�R�5�P\q���^��:�}�*�3�:�+�P�Uұ!Vi�3�W\�|U۩M��t�Urc�47��ݦNkY]{����~����-�1��
�޲[���.yK#�З�DsA���n.y])?�6�Z۞�<..!�>�?�[|�/.�bu�?5����>w"6�躄���>B��:������%O6�>�cg�� 'h�o<A��O������+��'��V�����r���;|gm�2��5�/=��j�M�]�R�{� �W.6lj,	�j�0�J�-��N�wr�2���7JJ�(����1d}^(=`Re3����rø�c��.����P�K��o�|���EAdΰB�j�}�{�;��1�Ô��m���1���yf����a��b1ϥ���*��`���V~s(��]�M�?���8�Z��g[門�p�ì��k	����o�����٩gv9�[Ka��XL_)=��k�A��,�JXL����a�U��@V"4p"�1  �U��gTY\%�X��R�n����ǰJX��(hyG��.��W�@�����
-�*��0b��U����){�p1v��XfVz��E~�R����\�(����jnok%Z���o�%�)�U�k�?Yp5e��ԉ^������x`t%��?���/"`�TzwN!��z|���g		�/�� �2�T���xE��|��ǹu� ��}���VTpq��	@�o5�����JY�iWW Q<5��:�o;m��@S�?U���c~ߕ��6+{��LVx�Sc?փ�Z����%��T�K�tO�mKY�E-��[�b��S@5�+Pӛ��^F퐁�Ke�������)P'_�޽u�Ҷ�1�m&OLH�z?�o+�0����\��]��u��P�� \	X,�,�eR�y?B@&ea]�o�� ���J���
����[�6˴,k��QM��p�Ӭt]y"�%�o;q�背�  ��q��pm�7i�%�?��O��� �q��Xb�߭��o��P�ٸ�2{[O3G��䛕�k(��T ��]���o��ҁ[�8N�.�Z����G�B�	���gP4���i�9��ܐ��5��h�n4l�"�,���0\:r��5ޠoV�pC -4�; ��7�,�2n�x�F��^�ܪ�p-� [�b��ȝcIfx�yE�v6�b8�8W���g�e���3{�ˢ������x�[�V_T��*�����.A�q`D�ԫ�0���Q&Xz)��*�����ɬ,����M	󹃹%���W��ԩ��Y;�����  ��Z�@�[����l��<��O�:q�:r�{>T=�@�~����R p����H{ v�3K���[v��QEW�n�Ѣt�u�P׵܉O�wܹw�����'�aaC�˽�kl�q���-����v�o��l�����>2���%��� zL���gz������ӆ3����Ɔ�q5�t8�����/�>����?.b@K4A��yw�C��e�~d�q�~؍�E������ Y�$�8h�/- [�<b��ZCZB2vp���^
�\@pi/��9��x�U@o��n��l���s�8ߧ�75G��*fw�G�<L)��̬��٣��.U[gT����H7���g/Z5H2|E���XN�9KL�ջ;Sqa�^*�ZT1�(��)���5��ow@ e�$���������������%l�6�9�����o��fl�rk�Ҹ-����� <28��ٌ| ����/u�� �qG���/��|e(��-��}$�x�5Xi�4��S	aN����5�
q^�k@̄ǜ9A��뺔b}��I��ᬾ�?x��ʠq'�QcAsJ@VV\�\��g�}v�l��x���u�,c�yC��o'A���MX��UҢpF��ظy�ĵy���(�����4��%D6������kU ���
�jS��3|�����h�K>�R0��V��n[ ��s���zВ�K@��U����͖>������ކ�~G�P�jӊ�h�P%�N����0����%9x�V(Z>�o=��id����YW"�����-�'�A	--"\�w*B�Q�]#�yExA\� ��J�c:n2L#����ry������ ���>ú��V�Q�Xwi3��T�j1AX��$��s�lV[yƺL�׹ �u}�|�@x�#kQ�|Gb����"0�q��"W�$躀ڏ~����9sfT� ql0s�w?����� = W�},z���q���Z�����^��B����J��0
�+�"�~K�V(d��9�L.j7�sȧ9�-���2����V0z�iU�% )ʓ9�eF���qN.�y-+mYҧ�n�[)3s�YJ7]�� \5��@���1[�F�#�r�h��d���C�d��� $/�ÚX�|{�t�>�Q(z_ �-�?���,M*�J���ح�9���"��]��^i��s@œ��j�E�z�]	I�=���ꍠ���ѿ�}rU�Md�h��0^��5||q��eI�8��饗�^|���b�j�Seݩhj������Д���(+7S�Z�m@�.�l���t��N WcU�E�Mc[ M��4פl�
��š�_6v���t(�1*�E�/���`�%��`�������{�޻xmc(s���RVa�X)�D]Pz)��j^�5AJC�?��o�6V<�5*cM�2�����.)3l8Um��&�����vM�G֏�A7��h� �i�rA��ɿ[��;�+�-N�l��<Z�v����{Τ��y���	�ITe�����̚�� l���?B I�H�����\�n0 ^~g>��9���nXH��fB@����X��M)�Os L۰���w��/�:p�MA�
�<��#c{a���O~���/�٭���YΡ�<��n�
`V�5�*�P%� ��sko��n-���d�
�I��/NԓR��"\��ո!�����rE��WCPҘW<?DBq�A�H����;�v>p��+��]P="i�ӫ�Ǖ�e��H�03Q:��(�����ukQ�K����s�Ȕ��w�E���P�R_�g� �|lWc��J0,a�s�>�`�I�����;%���#��A7������7E��#��T�eu�@L����߳K��ޥ�@�<�K��%lW�܍}�-�������vF���O?r`K�ۚ8���l;v��5��e	A�ϸ�{��3�/�5��FJ$��T� ��=��te}�cĹ0%T�����;������Ε��g��R�c�Bښk�={�6S�I��_�r܈��s�c4�7�ǏƔi\ �	4���D�Q�|��+�G/!m��ǰ�l\�_��ݍ�]�����˯�2575'Ug��J�V�	/.����8���	*Y]�ʠ4e���e 7�S=s1�g���1��;E0[����\��]Q��[ w���a 7{٥֚$K��h��b	e ��W&<"�[����`�,d���O�������`:*Z,�$8��� r�]���b^�k>}.� �\X=n��!>�H�o:A8c��j<`� �s�I�)H䩺X.�G_�'6���G� d� ���w��ݽ.�˧X�PV�������CKǴ_�*��)�{	�mե�z�Ω[��rAFe����Q'����
%'�����nR���܄ �(��Nt���	���Y��B���tE�_,�����̡hĀ���~��x'&���}~� a�䏫MzZ��:a5���TIr`�#�[eM��Vz�� ���R0憑LA�¥}�����*н�Ųz7�A�;�9W5������� m�'YV�5hʽ�}b�+�H�=�d���&'u/e�{�U�[O[g�|&P+-�5޽�`�� $����y�P�����_C�tݺ��	+B�H���el^�!�������r��9�A�/���L*7X���|�t*�+`��3όa��?��Y'��q|d�5�cZϣw��k�@���l���SYYQ��xb�Ǻż*�VZZ
x��=ĝ��o��M�Y)�rK�sZz��Q:�@�@��*���OZ�9�Qt%�\����=�`u���:��RO�W\	������'�0{����E�7|�<s����{ECF��ȧ������%��*�<V<��[J�Z��ޕ)|�q�[��λb~�)(VhI����Z�K�i���(�v�4`�E��_@��Մ�ޫ�w���62���*���[� �l�L	�W�#,K"�9��?��cx���x�0E�7 w��ɪ#�`��9B� �L�ŵ_[����.���(� @��UZ��	j������2�,��x-�c5�[�?����*���ȟ�3���mQ�v/ַ%��G��Λ� :Q���?��v�5k���1�<#��0����S��xD1%��c]���C|�-�C���7�d��S|�QrݢL~�n������W�O<H�V�x���-��e�(�+S㢕�=�֒^ϊ��읓�r�ռ%+�t��{�����r\QY�E~��3�9 e-�nE���)c	x�ʬ���j��V�nM�Y)ja��q�c�(Z"�"t�(��E���E��ݯ#�2D��}���'�yh"���%K�.���*����[]���8�Xo�s<�s�������S����t]�V��ZR��b�b�"�
�����F[4%�*��2���z��(d��Z�3S 6�S�%������� �T6e���^�n�(�ct�.mƷ�7`�B�(�UE��X�q%^��P�+�V�Ϣ��QN9�(ԏ�/�%Ȃ����m�� R}�ýM4*�5�S�'������{ꗥ�dt_��^c.]�z��5�7|�ٮhjd���ѫ/�U�=���-&��*�\�թ|����k���V& RV�q'�APw�\�&�Y�r�υ�X�����?��
k�� T��-��<�#}��p�uW�1���7��,�	4��_|���?Z�� e	^EKx��W��r��Eա=�H����X���^����{�ee�R`�(���Z���H >��(�����q^]�~ I���ǡ
������q���B�]�Ň�"x��Y��WH.p(������O"�u�'Yl5� �j�k�\߸G[d�af����z^�>�7� ���LYz�Z�*9�T���s��T~��v���k�G�A�ָ����|62�WxS�s���k�-��!�N0v���J������$p|����'O�VM����?��ҟ@n��"x�`���N\;6W��e�K��xW��s�1��F��[/�y(��_��B�Շ$U$,��>��)o
̗��JṴ�Z��T��1\1��ת��*ϣ�3�����-��� M:�x�,�HyH<�ݺ��f�$ �l�b��WX|���˯�}�W���v��F�	1�	����7����F���x}n��@��r��E��y�D9��S��̝k ��= y	�x׍��sh�ᮥ���Sy���-(jcЭ�D���&i�����^�|YoMM���ɭF��.���,��ߜ�Ѳ=�P�!,�����G��Y�7W����7 ֣�F�6�hC��8^Ng�GQ1q�a�4 �P&T�6��r��@.Q �Y�Q��(Xjq��8xm=ﻵ����k��w[[��hjno;�[`���d�E�Y��8"�� �$�=Q�X��FM����u�t��qͳ��RD���uk0����mGJ�#���w�_��k-�Q��wy���7�U}2���2��>*p2���ka���ʀ�����z�Il��u��S�.hg w.�ZZFfI��lEѺ�V�,������l���k2�
�,N��+۸�Cp
�z%�t؁��Nb������"@�^z�7�r�L��Ji9��C���0��]�%N�*��*��b\4#���"�s���@��,�Ō�t��mK�]2�x&Ư�5-�S<��oT��M� pVn$\D(� \E�eW��S9���q<�A����y"�/y�DR�`>���;"wgrW 6�i��F���N�#"���-ϼS$o�m�0|��L�1�2�R%�*�m�20Ck˝Xv�?���%�m>-%u�2PK����E�K��j\/��1��t��\����mFQ�'c�ZK4�Z���m@�Z���8��\�0���c}��)k�P�L��Dw�q�3����[� �z��r7�ѿ,��N໿]0��z�?�2 U�qY���VdB�)~�>J���.�+��귊v��p�0%L[�żw	,�� p�w��s��T9�K�>6�!��ƙƵ�)&"w )���k%B�<���+��:���s�#p?.ۋ�r̦1�"���uMs���cל������;�3n��In�c�w�[o��kY��7��G��
a�J�����R&cעp�vٻ�$�%د2����]���F��SX&4�&�-e�s�"��ߛ,c�5�cvo��{V(2G������hs�����>0��T�J@p�"@ � �q<��7q)?vH#��W���� ��w�˂�aÌo���4 �U/|ٴC�1	e��4�� ����P��-M\��Nk|�wo?W �x���{=��ˋ֘#U������ۿ��x��gx΅&����s������>�w�'���u��Qr��
����-��>7�K�NX�����뺦���a��\A1(�2S�K
�,��L�o�7��Q���� RFZi=߸z��W�X�<Sp��\y������dMja�]�٪KF&#}T\*CR|�J��0B�	b���WF�ܞ�+���%������y>��@���j�Ǽ�<���22��@��k�О�A;�&���^$A&�$�Ge��ө�ea�{��މ�Nl,�� W6����������#u�~�ڭ��QY��eN/�mr����$t%p��Ʋ������蜑z_�oc+s d�s�g�-�y�1�*�����J��h#�T}z��x�;�g�����Mh��R�� �����1���~Ǹ�"�8[" ������p��+�Pz���>��H#��P\�j��1gq[���bGk�iæ�G�H�d�ɼ����ɖ̉���1�Mo�ۘ���S�- ��c[dϬA/T�����ԩ��
t��s�C�e��{ܟ�9�����4���T	�
����L�Ί�qW����� ��j�j�T@aMF��,T�j�o��JPI�!��@�X	c6��:�]�R�I/�����A%�U'���X��E��n���`�G%�emx����_��~�I��wc����%��y�7m�l)��c��z15�e��P5����Y��΃��3��x�7��b%�mF�Q�ͯ�~��N@�����~�5�
mL�R�x�������9}M$���a��>l"��{h�����Jޭi��>S�)s�뜍Q����~g����Q��x/�.S`�'�%��U��2c;���^��u�l�g-�K�� L���PYڨ�������dX#�)->+׿��1���Ty�j��R��o��Uޭ2ǣG���������emz�G�4��H�q���� ��%����/a+�I����]._9t��(���{=����OV$�Y�-�gc[_��� k�nnd�l��'
�LxoS�Խm�G����m�\r�R�?.
�3)�Z���N�9']6?�Kϻo:�U�LK&@�;�<޴��� �=���L�D�U1��4�T���R<�]#O��7U�F���ܪ.�.�v��T��<�*ϯ���]����Y����֝��U}z��깵��E�������l��kK��pSV]�vڄ���(3�VfQi������Z 4R������ẋ��*7�*�(��~K�Iк��,���蚄��8u����1�Ê�XlِB�L��$��Xq���b����-��U/j,� j	\
hV�4��<|��Ż�X�0K�m;u}��@d6�x�R�J/�Z�j�����nCkX	����G&K�x�a5�d�%Wʙ>����Í�q�&5"3�[��Ϗ�e<3���l>�K��
pKqd>�n�k���ͯG`����d���\�7Sc�wlr��6�qO���ɭ@j���lɼ��ხ�AS�����Q.G��?��	�쥹��4�V��%�c>�ON�K'j�yG��ƻ+�a"դ��89C��;�Tx����&��zk�a�M?wb̡���T)�P��k1	JYee�x�o�,��gΜ���8I8*=�l4q�͆0|a%�J	���Mf���Y=�pD.\�{��ƺ������}X+�=��Gb���3�y���kQ`���4��[^+�ඕ�~7e�X�~-E?�	`��4���)R�R޴j0{"�D �F9<q�G����Xd���z�#`�b�F��﮹���e���Z�:Y-���9w�����~�9e�"��o6��p�)ј�Ϸ����4�ŭ�s�Q���4ێ��~p�)��ii���@[�#�h���>J��l��{���O��fy�:ƺƓ�b?d�����o��ڔ����]��Q֏(�G~be���c�R'Ɋ�Ih��b��Ǐ�KPk9�C&$�v���Ka�����o��,�hl��\_
��e���s�q��q�-���-��}��M�"��H���f�`������j�D)�^|���7�>���7�e��}��^sIV[m�6�>�S
���e}e������
�"�����\���}��ݞ���.���r���ylbw3����_)�kS6��*/ʣ��Ìz�\�����oK�94�Z��Y���3�L�Ui����l#U �wR�20������� %�Wd��ļX�>m������g�� ��}�4S}�����g������LBO�L[6��#�1m���B	�꺄)a�\��B�y �����KV��~U�M��5���Nk�ܬ=�i*�6�6'ߵ�heщmǪQ|q��^�&XJqUp`���g����4 \�=?؁�w�#T������M~`>3_|��󮧭��Q�"��~��'W����X޾���_���� ��=�[Q�4(���:ʏ�}��U�r��+�R��O�yĲ=_>�2������r�*Uk�,�����AKVa.�u׾HSi���~�s-a���4ϣ�j��h[�{�Z*��6��D�����z���1����t�3]�@�`��a�D�eN��Ƥ������6�Q��z��$Ζ�����Ȣ�eG�P�bJ��Hm�Q��?\��K�Ĭu�L[�ل�F�ȅs9ZRZs:�u��j�؇���������K=|li�S2$���n�tg����Zk��g�x�2E�@|Fc_V]����y'+���X�|X��~o����%̇(�V?���q^M͛)9�m��{��dl�l֟��������������߽\�e;_�7�aџ:�窽���������U9=X!˧�l��Y�(S2��>bӬ��A�-k���§�iOe�6��-�˿�3=L~!�Q��^�Tݪ���+2��ld81�O�n}YÏq��N.���?q�'�ؔ=���P��L|��嘥��g�6��u�ߗ������ i��Jy~,�$yH/*Sy��}0�����>�Y�c�M�/'2���y�yd��0�
,�-@������Gk�T�P��Sn��)���|��̸���>Q�< e�́�S7�av�,�o���@~)����@6w��]>g �e4��{����9��`wk�����-�"OG����y����xxO�HSm�b��11�^���!`ͮ�g<��^a����U���=���8V6RP��fL��e`zɠ�T�,����j����X�Td�����k`&���|+���_��-�R��Ѝ��?��-���2f���I�_˭ _��E~2K�n�\�*�75�3 ���m6�R��k����Z}��TZ`8{�G�L)�՘�Ʒ��외!�y�(*|S�@U��]�w�����u�-��g���܇?���kl�x��Ll"(y�(�bd�#�6������e52���5�|���)��S�ڒ'յ����N�>�YF��C2j��T��J��:j��&-e8���B+ �YU�e7
�5z��N�V���o}s��I�M��C&t*�jY��̜�^�ȭ���Qb�bapk��������i�w�yF%��n!vK�O��V�� Z�gm*O��ޓ�_{~OQ��-��Ի����d�p/�{��P�өgZ����,
@5���2u�����8U_,�D� ���?��l���r���p^�'*��ܚ�N~:��]��u��V[�P�&q�N)--9�F���9�������E=#5}p[�	�XH��&箨���Z ~jPd�=�$��� ��ge�;��F�K~�&j�0)�Bz_�bc���<��_�@[�?�?�k1�8FZ
� ��9�Y�)q��[1�8�tX��)���<����;�����wq�@�����ʧ�n$�q��`;+;��(�[
��#j�z�qo�d�Ekd+ߪ�S f�.Ss+k߹��A'nT����7�⊖��%-|�F�h�LZww@����s/�/�\~rR$��:f�a���Ȩ�K��Q���6��S���C�	s��=Ln���G��>@8��&14^�wMZ���kԾ���?up�����?�U�N������˦3�#��Lӏ
L=mo��0��ޔV[	��4J:��g���Ǽ[�3�]�A8d�U��{s��>QUڑL�T�gV�`�E`w�� �(*�Sc����3����,�8���ιT�w��K�-��P 4�����eL���_�+��S!ݴ�Ve2��<�2�� ��{\F�{�o�p}���ylֶ���Ut�V��������Q�l�[Yg2���d�$kPԄ3�_V�)F��N�TC�Ä$����#Z`�)�Џg�ǝ��1W���x�"�t���~�b�(���|���́�L�@}����!��)p�)= 6R�q��{˛K��[`�e��3�=+�UF��c��x�PV����띯 ⹌�M�>�S�-��}	^�%y�B��z��/*�;GA��n����l/�m��.��v��XN=
�y�E�I.�e��]�|ß��&A�����p��3�R@���P~K�_��������1��Z��f��.
N\p-ӂ3��"4=Q�����:gږ��m��yW@ �E��V���5f&lU���sҖ�K;��d��7b>zNIL����o2�}`}ĸF�H����K;�tx�C�y�+e�%�b�5�����x�[n3��M�T��d�:�9H�V"H�{�.ߖB�������:�=���m;&[���� ������m�aWJ*�8E���Ef��u��%���>��EK�J�/����u'�u p��b�pゾ���ʈ���� _�+�2��n��D䆎h~������/���d�Ut}+�����Yb(G�1��g}U�Y6Ǽ�Lql���-_�ʩ�э�� n�$�`� ���]���e�wr7�5�T�.�	!���s�}Ǩ�w��R�eI��c����r[er��!_�R�0@?p@�_����b>����n�Ɋ:)o��0e�)�T��MY�Z�U��,���}[���RG�Ff�&���W]˘x�z�[`��U�{D�����V=��
��e�-�h
���
|;U o�~q�M)	���?��q�Vc��'g`6>�j�xT�z)+#3Uc=��9x�����Gx6���r�{��";�N�E���uN��wأ0�Yʐ|��XwE��T���i�-�52�(Ģ>2��ڋ�%����C�{q�1�ሇ�|c?�s�"�����hݯ�koy-9U���]��>��t-�eN^=4n3�;/c�NS��֪D�V�` �x�$���;�Eb ��C���gƣ_ńD���OBs�sbH*Y|rU����16��ha�<��bh:?^ /��71�����,�枾X"�{��fdzYz��S�&���-�,rE"�H�;���E������f`���f��0�yTJU/��Z�����,��s�{,g����h��9���/�A`����OVV��U��2��Sc2�p����z��`�ik�+����`"٢�d���Z`�hd�g�!�R>��AN�ت� |ۉ����5���'�._��1����?:JY��}�iCQe����q�d2a�b�����V]�����UD��V>��S[5I訐��%��1���.�5m ���� ������ԍ ���y�b80�9-K�M\�ŗ�����\�\�X�mO��3�
���-�bL<��/���X|�p!��h/�����|�3� U1�(0[
]�.�g��n=������1���fm�:e�)�-@�s��ES�N~�^B�����}c>^�^ �j�T	H�SyW�;�_P� ��y��q���xtp�R`E��z�����w�U�q���n�N�� ��� ���icnv�8�q���I��[�߲���;����ul#;$���� w� )�
V]�މ��p�b���YT�J	�UJ{��M�J�KS�U
ٮh��BKsy�.�����[�(��W]s�ܭ���#P�I�0�wM�c_5��l �Xb�-��YD�V0|�����B:4~��E���UG�g� W�*�w�*�s��%�p�T1�L�e֖J��"����|*�[�a�x |����
4B��#.��?��צ�3�MK�j�V^^<[�����l�J�h阏��f-���?��1��6�U^�̪��f%��5���)7�z ~Od�KVļ�_�ܞ>}z���eF��GOG�(d
�
���X���_d�>ʓ�%Z� �tc��o�=nN�,�t���j��O����'P�z�T�;�z��%��j�k� v�����ѕ�,K�\ T	�Ш�yeL�WLB�I�]&>�S}��j�j�M��a����KNb�A�����
�图܉߁-�K��\�v�%+1�ri�ZR�G6>�0^����}���e��P��k	vQI��"x��|�  �S��y�:�Mhx8cc����'��:.��VF0������2���X&�Q�+!����6q0��O�L��T)	^߬�[`;>�*3+����s��Ĳw	��|p���������)�l^���a,Q����s�������K�o?��(���DK/�F�>#P�J���җ�b�o\�/��$
�b�U����}A�S>l��[uV���#<����� f�z�W����%�eڮ�D/�E�FД�iAE��_�ҢZ�g��ء<_V���:�3@xY��tl��ՇgYZ���z�~�͒��9t�ጄ����í��4�`<b n�ey�ݴz1���zk\N��-?*����/ ���t� ��d�}Ќn&.'�G��4��!ʫ�Ϊr���7��t�����ǰ�)r��:'�X�,Ԏ/ozeib��X��Z�(˧��M	�����lTe{�ٵ*�yS��O�r3���ž�eg
_�vj��\���;��;
�Ǚ%�MK�з��������W�1B�����%�j�� H�I���#0|8��n���h� 4�+|�ظ�;H�HFHF��z7�]��I���U92� b��ԆQ��b贬�����:���=<��{=��������Vt�+�-�@g��� �h��Z�d����2pK�>8���֗pa��X~<���u@T�V�F��
8����	Cq�B\z :��-r��C�����3 ���w��5� �����ob�*ߩ�g�}�8�sov-�5~�hG�".&1*E+|�SK��hl�sA����2 @?fs�
�_x��񑽟�]�d�b~�+��q��}��8�����l���wVG�IU�J�Ƽ�X��U���|��1��1ME-ٴLG�Ue���5*"Y�������JIS:�O��|h�s5��kE�qd��\"����>���|��pE���C���w�H>�o�z�W\�$oy?]{��w����?l,�<��/�}2��3O{�ԃ�b�<7��f��JT/�8JZ͂�j�9��3Z϶�_&�2a�	��VKƈb�^_�Ħ�9�t�-u��_[�l=��8�38�8槢Ep�o��yG�T�>s.m�CP��fo��eR�v�;�#W���+�KVB��x����vn)]q�F�25vQ ��s����d�%c8�̸I�E�	,"q��Ge���o�����!wEaD� ��8?2k������G�7T}X7Q�-��"��C�"6�_�0�xqū[���\���9Q�1M/8���-!�����w��e'���qf|��QƂ�|h���S�x�x)>�JC��E" �(�~L��Y������(�.�1�x������L�0�f6�]���]��zG��g���9����W2gJA[
n���*TQ5.+E�F�Ƃ�-U��{sG3��z&K�i�QHeyf`#�ր�h,�ú���&,b����<��IӔ3�ɓ'G?[MJMt_:a���l4^_ҷ�	���,)� _��y�@�p��EP�)4�����Gu|��6>S�Q�)�-d��}���43��NƔ �?��w�a�R6T��T1H������;z��%X �?��J�7�/S�[}F�I���B�!��o��=�������}�/>�qS�{�<|�d�y)-�qR
�E%��#� д��-��7��d�v�K8g`3��=�^#@)�"���"�Q�Ot0��V��k�_e|�E�B4Rpz�R���֒�纁b.���U��o����Y|���ܳvs��}�	gΜ����??��7 ���R�ޱ��py��n��,��@��姡���Ä��n��U��	lFCN��ݐcJ�j'V^��2tםw��~���<VQ����Cd��Y*�囨��ҫ�e��~6��P���r�Bk�lKq\��֪.
C��O���̇.�)+E���2?�,}Kz�W�[��a�%�C���7M.�(B��K$3p�2j�X��H��7�]�.xa0��}���G&g~�z@��7	t=��#�屗^zi�K�-^�`��l�s����YN)W�-�V ����X}��Cu�W�7�|st��*o���\u�Oe &��� �d6�!|ܲ
 �2�!�pYa3�L�:ч�?���FF@��7��0c<��Pc h6�C%�s&��AD���ݿ�!JV*H_j���#��	��+>��ׇ�">禄K��y�����S]["sz,[����c"�o�#�W�kK�2}E-�C��T��A�ĳ�W7x��N�l~g�E��;���@	y�K�!z.v��G�����WAI��-�1�+6.	�?����9���0��:����?�֘��w����-S�20+��{����T�WѪ ���:4"��5�)��J۲6d�-|�:�� �5�A�tbF=���4�t���pE��U�VNBn�Y?��X<x�O���D�ڀ��;�=������w�u��q���s,��3�ݰ���ƪx� �K˅����	�4ƈ�:q�����u]����ɮ�ʗM"��@���&ƬD��t@� ���
�u}�@�J � �j���QyZ��W�7}9�5��m�a�P}���"��-���[�\�f.�\\oK�+c�;O����ʟ~�����~?n�f�f�!��?jW���+W7�,��,(-p8��/�˽ed��e�ʏ����X�h��T����Ȯ�NS�_���;F3q�#�)^���AQ��#|o��fR���a1�%s���䴑��z|�����0�����A�'�ԁ4u�d3@2��J��!���/������\NH�2�\K��٥�K�@�S��m��t�Qb#�@n��޺W1���^�#Z��w�L��ŉ��R��/f$%˭@� ��lB�u���P�l�~��3+72	�bi�=_���b9������G)�����;F��� ة�j���C� w-�_�Ug�\w����8����W�Wc���o U�R#��~`n�=v!B/�Ty(/�6�����2@?�CT7��h̹��j��5Y�nծ t�MϿ�⋛���t���u&'m�v��<�-��ϯ�y�4G�9�u厱W)m>��{��7���pA�� �盄�,�Z���x�=*K,Dk
�� :�aέ��hy��3
#M	|�or[��@"S�*#��}����q��:���ĸ��ͭ�J�������!��Q������(?n��Jþ����g�.{\C�FY�}�6�~P��������' �j� �5�ә�)��si��8��m�&�w	ź���.���:Ue��V���[�Є3z��F?)���<5��cq?$�`�G�X�l@/Ve?T�2�a�"���8�v�5�C��p )n�{�����PL������DZ����q �W�lc��k������
@�%���3�((��.�KS~;��Z����Ǡ�
��
K��@�Nn}P?�)Vb���b�`���1���Gʒ����D��e�B�Vm+�M?RG�Q�V2����3�����	����y��V/ڼ�EոB������_��_��"����
�o���L`g
>����-���[�P����1^��zJ��g����S���Y' ��R��:����F�Ĳ1��+)�m��X��_8�u���퇀7����0�S�;P�(
��h@*n���p�Pz���b˪������G�R)"� 6Sn��� ۻ��6n�@T �Ҽ���#��zOYn��,糔���7������ZM8��c����L�� L�.�#�2�&(�K���wa�E0p��E�`,;�O����|��[�h/�U=�f���ǁ���/�/gyͱ޸O��rA�&/�G��c��[��{�[�'Vm��MO�mx�3�+��� �M,[Y�&� 6oh�ʺ��K�}��]	�.�.Ҙ�"�U�7�D���^<f�L��6��8�6����r����('�M���5��I[T�f���xoEsAn������[up~�5 �KY�V`�J��>Ϩ]	�ŉ^�`�2]q`�;���I<�(8�!�i~����<PZ��C�� ������@�V5��ȜY�w  �Q�Md4.zj7�6�V!7هA�E��A]N:ߩ��=�\=��f�S#��ì��z؍�s%�|�f�n�a���	@�tl��ʂ&���*p�C���Ű��q������ b�b�u�6����D�Do��V�f1/��)`6n���x i)�6%�@��LR� ��y?V֞��\���0��5�^D��/'ރ��mܥ#�oW��-(�(��G �[w\�ѿ��i�p�
�b���ր�D9��.���1���� ��ٷ��6.|��2��X����O:6����6k���NY���OW-�5��hҢl\d4e����~$���;�Q�cG���(�ίP|���7�r��!��t��H|��;m�nf\c�����ܨ����$�Ib}1�(o�r�m����ܺ^}���e��߸l��7�x�L��o��lv�W�ݖn�흄���K�Ψ5��L@���R˳��H�&�i�
`�G뻯9�����eo@���B�������z��Sh��)R���.��\�9��خ���F����
�e]�Y,�w���[aݏ�-}���Ue|�?�	�����S߾���7^a�v0���<�P�]��aI�L�X����Y@���l�U>����J���)ДN����4�{p�rD���e$��J1��Oג	���)�ɕo��~k��T{��q�+W|S�qT)�{8��(A�q/�<�]̯�d���#��,=��F�r0_�_w�b�e^�<ہ��I�%�AX�U/���k���k2�>H�w�?��ZTm�Ի��9ً���5���v96���J�;�֚_#�]��ߢ�P*+�ԳY�ͩ��w��Y�Ù@�i�
 �#ޗ�]cp�rș3g�o�
(?��z+P��$` �5�	p��x�����5_&1Y��1�~д	���f'�Arz���&���9UB�eug� ޙ��8�~b�Cgܙ��ǲߴ��ӴG �OTt�0�'�,t�ǔ2���-��Dē�`�ԉ2�rF�y���[L��`E�D�aT��_��~�WHK�x[yY��z��d6�3�K�e �wF����~v�
�&��M8�����w� ��^��|�ߢ�S	�Li�*;ȕ�]K�V�������'�yTV&|_�YrG��9�����L�+e�J	�%w&��}�����[7�U�q�G \ƺ�U���.�����;�g䉞G�1��e���#��̜��]�|���V��Dm$Gِ&��<u�q�m���sF�x�����6| �1�{��Z }�>����D�e��4�Z �}};�� P�5�OiYo�aC�}I�c11i�H|"��n�T:]�KZ����GUi��#��Eރw��xO=/_T�v�X�Q�Q�lfS:4vv��\�;�ԇ �h������=�>z7?��r�!��cx2�3��jL0J��[[�:YY|�U���7}�� m�M~�}�p��ؒ�\����6
��.�f�>SH,�#�-R?_-p߹�b���@/�2xo/�g���d�2�&c�w�Ǿ�~�,"���Ɗ�&O�����Ʊ����^��2����3�?�9q�:�r�Xo����i܈������.UY�E·���k��߱w��u�I��9���z������!l�ᢇ�C��N���o�<�ַ����VV�p/T{�/�?��'?R�jnʭPu�F[�y����7�L!k���*�1�����?J����(d�ԫ������y3x�~���F�N��V�Ciq��E4IK�Fs��$�q�u�CF����K*X���׵j7N��ɟ_TG1�+�@�<�(�_/` �8��	#����bٜMO���7MD��o���ßM����NS�|](�?g��d��W@.���;h�t��#�%^>i:N�p�'��z��,+,��|l�\n���v��wup都+W�l��s��*�!�F`,S���(�c��1�K��`�u���9H��oS�o��
�̺�uqE$���J�ϱ��ys��"ʀ|T�}��>V��&ne��G�O�+����|�_3���y����{Q� �CyO��	ɇa�����\H���D>p������:W6��bݦ-�@�o��A���h��NД���#�����8�_h?��v��KŇ���r{yL&[�{K�ۂ�U��@{�/��]��ʜ�ܺp����{c��`���cwI�I�Dcy��I�:�����޺uSu�ĔŌ����rˁ���C��:�~z �D�Ͼ��8Z�-\�ǲ:�B����h)~�ݽ_��/F�C�'=�Xq�[o �
�|��ҝyec,ZP 4X����C@�������i�?�Ma����������=��U�簌|�����я~4�����b�X��3��|�ͽ���cmd	����#N�_.D��>؄��b��-�����a�|�6ʭ�y x�� 
���i7 ��rt�B�=��{��8����m�-�V}e���uK�~gV��w,g���5�2��D;2� ���e���jl1^���R����^�uD����w�����n�m���G��`���KOs�s��uH��g>���
ܷ�:���e"&�W��ѵ}�Bwa�� {?��9C��x�6�ÿi7V�$�<T���ќϒl�<��Z������}}#�R���i��h���f�(D-1
Y�C���(�:���Y��w09cfw9!�4Id�GJ�p��&��?�����|��3�&��e�GK�ʛp`_�����&���=&-�`g��h�kOWm���/��g�䗇�]������XR�-�#�"���}�k�EN@�O�wr��,v,E��s7	.C��(Xnal w����c:2�L!˴�Li��U\S�U�����rc�g��5�}����e�2���I^>W=�[�>����g�lJԻ)>���h�q�J�[�=ړ:᛬:��7�-��Oc�C<^�FA�ru��b�q���`��������|dY�U���E���HT�<�'J���}~��q)˧�{THPn�~lj�Ko_��5xlE��Ǎ��8��:9W�e z��7U���� ��񬈱�f2�-W ख़�s��W��b���R��,���;6�`NDWyz�������ӧK�����~V��,� �=|d�cC���}͆lQ�F���o�v����rÃ+�>Ȋ+��,�1�@V���^�)�����|���[6��v��ӷH��4˂�7R����{�F?����{ꕁ�5o�[z�&f �x�0Q8��M$K�71�Dy,X���ɩr����:�O�ɡܧ��]��_��!���[o}{���8\���o�qn��>�Jd	'u�g��_c��xwl����oy�7j,�,G}(c�c1q����Hψ�i���?���M�^� �S�xWb�s�i�Xx_��'m�@ y���jl#�)�(�ow��@-ZB����w1K`H!`..���1�"��xo\D@����G�T$}
��z�g��Ee���P�D�ɕC���|�+�ܧ�Lq��s��[=�G$��=�=*��O2���hT�v���)�Ғ���2֕Rw�q%W�߳�ϑW,ã� GPΰ�n���U:��r�@����!�!��2�-�h�=��կ�@��/��e�pj~ɨ���f3��@0ql����ǐk.+O�_Ny��|�\���d��
�6`�F����֯�Zs�e,\B] �%��>�i��oэ�T2�:��[˼�ٌ���-4���r%�;��dG=Z'̋	�;[��,�"�Ui4�4ɱ���A֣X��vH��C=�
��:u������'���/��=�uRG��- �"Nc��I�$x[# ���U�M:�v�;ؽ3r�(�(������*_��^�{�g�w�*�% `�>׾A��d�eJ�/i"X��n9�v����F>����L?8�qA�ׇk�Z��*Byå�-\��EXr3�_d����!�C���F������)Z٠�5gY���Bm�a,l���x��6��׹��C���7�~=��̨��<\�~=������O�����oW�P��>���!�ũ�X���2c�ݙ�e	��@��T�+W76���;C�o����#��f�@���Ɂg���Y�)��
̪�lx�>̏��s��c�&(*G�.��������ע�(�c���L�]�� nŴ��bp~/c���GAs�=��J�K�XoY�1��})F����x�}|}3H�a���UTe�����@���&�SgΜY�V�/��/���ou|t`(�����F��b�hĲ�u�ü� P|��FA ���mN=2�K�(��Q=�35�`�Db�1b��w_���6���矸���o��$c�����k�����c��с���#��s���K/�p}����+ .���Qļ�m\�u0�u�3�m��'�SJ��=��_:!�~j�+Vq�@i	�����@��o)v���GP�m<s%>έ�۟u��#KzxA�U~��}FQ�b��P���mV"�%�*� ��Y9��>�?[�-�7��h���={��q�(k���C�'���.�m�x�;���7�w:7�ǥ�3��ɺ���8�"�&�w������ۼ��S[��	6��z�r7=��W{���g�Gv?��~�A[Yp�*��H�N�4��qҏ�MG�@v5�*���o�^��0,�V�E�ǗDc9���3	O�*�H�����N�>�� H�����wl�,�O���A�=?��Y�����.g}����E��
K
�!/`���?v��#e����׌\8�{����'�$�>��/q�`9Z �8�o��P���h�x�5����k<��1�sE� ��i+]S;�=2K5e�GL;b� � �}����}L#���5mN��L꛷��M^,�z}q���Di�UX����O�O=D�^�1�0C�� �0Ɯ����r|�<�D&D"�����ż�����(+�ZY��P��hZb�Q�Tu�_�=�wo񛬜('�=T��S!��;8���h�u��R�
@��/��G�-�����a\>9�n۵�}v�h�_�ysV�
���}@߄4T�x�oW�}�^��$ƽ����4�%�8�I�^}@XPdN�]��.�P�Zإ���l��m�v6/� �&�]
l[��1��Y:C�6��:Ek�6���#�q�O��{�1�}��f'����ߙ�jgL"1 M<��LHi�ĴU���7����/}g�����W�/{o�k�U����܁����U�v6��H[l�UQ�\�O)�s}n,���(���T��`b�#��q����ccs��۪�Y���ٯǘs�]��T}���Z{�ٌ9��}�v��{�I��{�yh �'�6�ڷ����&�̾�9`�Q�&5��V�t%P�� ��L� (�\7OHJ�e�{�+J˯�ԗU0j,�B�!0�Ԑ;�p]�xN�ݹNO��Y ��1_hc��;���)PY�̛�k�'HUp3L��T�]Z2W�I>C��Ω�Z򷴜�Z�2�J�+c�ӳ�dKl�ܼ�{'?L�� ��Y�4V���.�P�?�i	�v2g�����&|=�a�'(� �uϖ��Q�Y[߷�j�|�vU/�c�"�:����G����u�kI>����9i���n�`�ml���p�7o����U�$�{�=��'^xᅓ�sn�����]5�T��o��䍮o-��1��.���-��u3wj>�o��oBK��& �b���\JUQ��tSM���LudN�<������+��c�-��L`PdMPk�fI H!)�Q����&?[�`� %VQ�Ή��J�6�� ^�90�om�wx�m�j��g>���yvy~�T
��OM7S��!�P ��m�,�)�y*&ާu=�w��T�u"����o���Ѫ�Xf�I�I�%�����Қ	X�o�0e�t�7C0l�q�5c��E�-�����~JQ�ߍ!����$���M���i��s�9?8z��Ȥ�
�r��u��fz^ҭ�[��Z�ox�S������9��~�|9�m��%�kH�չ>%��\������Ӗ,�O�����m�\��Z��[x(^<<��sk�� 32�8y��W�m��
��7rl����$p+�v�m=��c'>�ό�C�&��V1�T:{s�*L*��o�/(�|�G�4�P�TL����~�^�A��S�>u�� ��ئ������ί �����K�}�T��ܽ[��;�xd��-�I)$eH�"� 
�����dQ����}�K_"��-��t�vt!=���@~rx�-,Y��GWG�:�._f�l��jۖ<��}��--�5�*A����,H&%��]�z����Eh�%�H�R���+�r���gbK�Յ2t�v�O�(��(��� YZ�XWAs�֒;�M���b֝۲lN֑��8rM��003�3�.�ئ�m�y�K!��?3�,�K�`Z����^Y�WA�uGAwų�rι�6<����Z���?�WO@��س��i�q���8T�xmcm{~7gᒼ�g]b(�)�B���<��G�_� �T����	�$�W�ޚ�DҲ|�칳�cy��ˏW�q- �QJ��(k��X������3Iw�u� '���ڽ��#��y�	֠Vp+���|N)]����:���-�un܄��BF[}S�i&��:[�F6��"�R/F��m�S֧���=,]`~7��=�^&;0��-k��oZz����d�"��ͤ�}d��0quag������_s>��8O@�E�%�~�� �n�n��Q�&.w 7[�}��x}7Ѓ�
j��E�np�aR
7�;�;cV�5��Z�v]�ȅ�����b��1̂�-�����Qr��ѣ�pk2D26K��*�ِcW�m��b��܄��y��@$ږ�x��O�Mty��Tp���
�,���m-�'Պ��!��E_poc���}s<qZ�Й��m�\^Y���ܙq��A� gܯ�윣O��[���yk������N*^yL&Ր�u�%���z#*�ͶdXE�8e��5�	?�Xj�]�kR9t|�?��:W۷��ԣ� ��P�Z&Ӻ�������9Ϋ�M���\����D�u������cǎ}`eL�́���e���F2x���LZun���<N�
듾7���E�w0&Y&Tl�R֣ޚX��B�g����~�F!
P�c{��p���;�չK�⋡�YJ�I(sM���KF��H!�%ʅ 0�1>�����9����G�����Ьp~b`'_}�խ'�xb���>�)�?Z�e�<�5h��)p���\�Lk�nx]�-�a˂����J�'�����V@�3�0�T��r�����V�N|&�q=�a�p���.�a?�O0�'�|r�8�c�,�n{d2^�]ZW� 1�σ�֛��J��s�y	���N�1}ٗI)��5v��^M��$�����X�٨"-0w
�����ʑ�'�ᴈ�W�M�U��g��>���+�)��ρ���Y�2��HD ����|O�v�sߝC���!�ZA�5Ń����uϓ�:��iA���beJ�{���W���XG����T�2�4Ϸ�m^W�e췫���j���q��w����1I��������G�\�(�'���o����(��B\/��/��\%[�;5'Zƚ�������0Вg�(Da�by������K�V/�,�u)(�c�{$8R(�$d� �ڰ�,Y"�w�VH���f	,N  �;� �1�p+��:}���N���+[�Ң�x�#�$�qǯj�K���#�0�xt�K=�d�����M��P��q9���7�)��رc#���H��_��� �c��uV��M�#Ų�c0rj��^��nX��uN�(�����*	���*BH��f�nyw�p����90�*���d�{f��"�&(
4��oֲ�rJ,1�����b����賯M��]�o�~��y��Ь�P�*k���V˱��:�]G����A����U���y��L�s#7��X�<Z�u�s_炉�*u+���U�FZ�7���I�1��+�X5�1J˵ ����d4+�d��9K���!!o�����<#����7��g�
t���!�5�IU���Y�:<��-KiS�ަsnn}T��I�[L�a�|������
J{V���Zz�U�@F˒{)4�%�Q�j�Pe?�V��1�;A��4)Ee�+�X�p߳(�Y0;5e�	�&�>d ��O~r��UG�{����� C�9aܐ�:-e2���R��8�6��*=P�����>ˎ%����jE�)�`M�x�v����;����(W���k�=��`�w -a	�4fR� ��;_�
�f�-ca��V��<���V}�ނFc۲���`���1�&�)�����kז)]��q���:�2`��rc�\�d��m?y>,��5k�u��8GΜ]xÑ�Ǭ�P�z�Gzs��QZ��3�`�Am�#/� پ�M�#�Q��� ���p2�����G�f7��]k���|(%�W1��-S� mݫ��7�-�[뻩���Q�����^����lu��7�����H�IZ����GRƤ��f4;����w��3��a^�xꩧ�{gg�M�$V�a^j(HRaw.�7���_*^�0+�q�Tt��v*Da/V�sz�>����E] ~nYe�B-R�3�!�^�כB�=�\�i1������j� �Z�vi�w�Q=Z�>����KHP�D5t\؀3�ƣ�>:.�(���}�C�t���/?�ӟ��}�����2i嶮 @�~��Hu1�J@(3�Z ��%rK���9&
s��3vS�TZ�2&�k�^�l<�1�2W�'Ϝ
RZ���xy.7��o��
�T�|�j5�"�u )�LX�V����#iȒf�uH�uZ']K�L���I��W3-�&�������w@�@��n�-�sG#� %��8��Zb�
ڡ��8r>�
��XH+[���,Z�8O񫜳�K���o�v��G)f�U/H�MC�^V!�1�ܬ��y ~&�UԽfU�^r�rL[2��k��>��Mxޏ;�s3+�0�"��6������}��= �y���aK��g��xӍ�[n�e�f��,A�Jt�����Kn1ϋ�]�;|�~r<Vr��C���w���6;L��T�Pf���k�/�"��j��i�pse@z"��07G-�D~�������i]#�D�y[׫2d0����B��	 <>���:Ď��Ӱ7m�&�	ȭ�$c 3�ZF�u�2�9�����<�}��k��ň��B�w�w0�Sfp+�����?���Ƴ�˓�Ϩ
���s.-��0��Z�R��y۲na��R��km��QiхZ������k�;l�n�dY�!-�?�����Y�Ƌ
�j�i&F*Դ�d��! C�?<V�� ��f��)$�ʈ]��#wcR��y�3�B�*^�Ck�a����JX��:����wc��2���d��"ō����ln���Ĭ�"���p�<� ��Bu��|�+c�>�����ZJ��c�a*��_�lcɪ��ŬkCj"^]Ǯ��D�U�߸>�ᮻ��"ru	�r��_K8��>S�V�mY�ɧ�9%��K�\y��e!&��  ��IDAT�Uu�g�C�!����K�z���g��<8��24�E�B��3�<s���	�B�EY�V5���T�U��G��7`@a�3>�U?]j��bI�LO!�m�����P5k�Z���c��ΫF�j��������+mr����t��Q+$��Ç���t�P��#ݱ0-��%���[���ȏ�.b��_��'�~�o`��X]`��1f�~��l-��
^���,��J��'�Дb��o��㮇t!g�U���k�z��K��jk�q&5�Ak�� ��/C*������ԽoV��R
*��k�-#����ݖv��2&6����s�
	�u�{?-����O�I%�#`�2������|�/U�gz��-��"c������ ��k��9��$��>Xmy=zt/�R�2�s���
W
̱��6,�uA}� /�/B�$���e_�Hi�D���}_���wB. y�iL�nd�	5P�zR�����M ���ʄ���&�z��9����Dk����^�y)����������#�׼$׻q�Y��Z�Uv�9���JCʺ��ٳ{��T�Q5:N3�sO!k���Z�5ғ�=�2�_p{̬6.X�������u`I��u�s�����΄�K�k��X�������3o�-B,��~7A혽}��!��m�\�wn�����W�	C������6 
 e��lE���i��y+3	 �e����������)g2X�F���~Z�2,�VpH�%8�*�04F4]�&d�'�+�o�5�6k�D��9+��I둕C����w͊OF�p�ǵNmf�ˇx^+hQ�+�U�x�\Cb���j?�w����qf�lx� �(XX۴�<���k������m��/|�c�-VM�V+zkn��Sy���T@Ҫ�s[�y��k,2V��uv����вNR��w�m��x�u�ѧ���b��bE�*�t1�^Y� �������}iy��8�ZK�:4L�$��R�vu��
�{o����7^c����i��~-�����dP�c��p$�5��s.U���� ��/�n�m<����6�ඨg}�ƥK~��-�8��=4?���h�L��.�!�~�+�Hkٙ�gve��c��-���C��`Ը�p�y����2���o��
�l@� EZg+�U��5�5cYӽ-�R��n`t���
_Ǝ�T݃5����3!��\���\�?�ziq�Z��_��s�1�yo]�V~ ����1�� ,y��9�� ���V���V� 7B�Bg��؂5��5�;�xP��7�����׷�`� I�y�����L�3��9a"�Wi�����-|���qˎ������8e���(VfO U#�}�[:C��y���	�JR�y��bɥ�U�R������5���b�X2_sW.-�Z��T���x2^��K	.�.V6��s,2~��ƽ�T[�8yL�AV�p\���w�3��粱�J�}��G�x�m7�P�Փ�ו�5�9�(y���XX�B�7/vɚ� }��3RN��q�m2�[x�w\b��u���{�I�������Ki
h�ڼ��[Ee���c3�%��9�[ӽ*�M�V0K9�t`^,@���e�Pi`ڧ��e+߱6.��X:�
'�Q��VT�K%C+b-r_㒪��*(HW��C�(x��)x�5xs]�	�<�9������9�8W���@�*�[�c��l��f�s]�,��&q�߱Fr<	E&����D�8��N�	�AY�M���7ɋ�t3[z�W�A�ߎK�)��u �<��Ҍ���/�ɵQ�0q��?�^�繣�B+A+�R�O�1�Cs����i�ldl���8�y��9'�}�	EΕ<�
�I�!��$��kZoz,�v�y F̬J�J*J��,�a�1ǣ���#&,�˱Y+C�xg��;N�ђ�V>������d�Ty���/n�b�^�
�3�.�����w������4��^~��{�>��(���^�0V�.�z�P�X�����Ӌ��o��1��-��.�o=o)�k�u�E w
�������X-`{Y�{��u������NQ�E��^��Զך���B��6�'��-Ǿ߃�>��ix����?� �}Clӗ&�XW�{��3� gWn��!��nYa���:�	pH[�1������֘���)�;�Y�57���x�~-A�}�`_!�o�č�?�؟��~��լZ}}(Xݘ���n
 �-�;`��VK��6��)�M��0�jg���3�� X�`�5�(~Lju�3��ga����l�:�7�w�2�7�0lA�%-�zpT��wyj����ʓs�f"_�wZ�SX���~�s��AS�GK��kM����זW�C�,�����k����r˜�|���v�I����/ca�V�|�)��}]ǩG-�4�d	92�[��L^Vk��X��mg휺�bo+����}�{cX��(5Pi"D�P������p��y��2������Yp[�s�|l����BKϟz��5�����Y�BP�K۲bNYQ� o=�4�ڸ���V�k�	����Ȥ"]e��2�\+E�r�Z��b�V��Ig`l�� ~��L�c��C����OϹ=��>������!c��;���*�ݪk?k���d�n�D 9�C9�W�����ڦy�aH+� ��2Q��HI)�X�Ӆf����>rޝ.�l��b�E�y�k���J0�Z��-C����%����p=��� �=7�jY���)0R!�^�1��~��F�m��J��jh�ʆ�1�Z&̹�D���9Vi��3�3P�Y�\�|�s|���Q^��U>^��L��{��v�& n�J� r�O�7f�XE>gȎ󔹄E��,w�B�or���`Z.�|Wפ�m�~Yw{ f��<�e8RZ�{*�u^8��>7��J$*j��RrYz
�>s�yi��|v������7k�:	 ���E�D����u�e&'���E�6���������M�K��������,�K�[�)�z�1�!	Z ���o�L�)��	�I�"5{[Ғ$C1]�m"��e����}�ݗ=���A��̳Ϭ�|��u�!�:3��F-��D=��1�YOTp�1�<��[]�X��H�)G��C�H�P�N˺%�5�&+07z8x��V���L�������K״Ǜ)�� ��VҀP���u�%tC�&tc�=z���b�;w��u��Xi����} /�{"�A!�bq�U5��p�U7�Z&����7�˶;�xw=� �m��%�r���_��jM[I*Uqp^$��	��	-���{&�f<y�����ڴ�疺���$��g�U�������M�����2c����K>	e�?�3��٧��m�q��*��R�|���&`7����H�����
%_��;��hg��\vYz
���<5�կ��6�!���W_s�hH������6|�^�T,�:�NtVQO`��0V����	��P�m�[w�"��[L���KL��jֲ��h/�h/f��w��2�d&
Mݕ���h\\Kf�%̺��;~�rIF�p�C����}�i U�x~���ܢxd�C׳�����[Aƻ�<��|U�aƂ�@�aU|YF�몘h�4�Q�7%�<�Rr
�t���d�֜��� �x_��X�L��N�$-��.I ��q�4�s�n9l\k�$��;�
�xv�sox����k8�(������.N�c��0-{[�����Pl�aw}j��L��Y�,p� X�ƶ�*%�U]�Y�z�l������]ݬ&�%Ы�b����OE۾��x	���Z���\���ʫ��R&Y��s�8 , �����o�%���J�|��S��1�i�m%j��
V��=R��=u���������\�os}xM�M����٧p�.s���;����j���ԮE�b����c�F����}��H���PD��z&r����9ך3��}�A�cb=~�NQoa�i��
R󚕁�']�5�hM-+�$@�cji�s7%(�P���c�u�"p�50��.sB�����so����U��Y��Jᯰ�d\�1���Đ�>
�LRx�1�:��׬;�%%PIWV,HA�u�r_���z��2'Hk�:���i8D*Ʈ�W�U�p�yeW�-�n����Xб�V�� V�z+0 W�
�]�_��������RX�R �q��v�ʃ��y��M�����crL�c��_&�	&�bO?r���%�� Sp��̾u����saK�>'��.��!�O��3y0��P�=S��>�)�� ˸s_����v�-�n��TX��\����]�~O֥�q�9��3y\]�>K�� Ĝc�4�3v�q0�ک�z�KM|@hx����zW�k��ꥢ-/w�f���G������V�̫�i�_����k����B���Y)�RＪ�|�@.4u�RxK��N���.S���$]���Ǯ���O>�䩡���2�!!PO8�\,ϻIk�(��8�ZôtdX�c��Pi������&��ݒGZ��|��т]ݓ�-㎹�`���+�v�7i�i���p�O������ײc��1i	և�[\�PN[�o�����#��Mh'���\��l�ϫ�1��s ��F���$�Si�7 ��(x���j�w���/�W	 �2�y�T�>�v�D�Y
�l?$ U! ;g����img��A �U/T��o�}X�'��V�p�z�L��k��2�V��y�oZ��ȹ�  ���F��cX�{����]���R�Y�����߾�>.�?=D��1�̛����S(�_��X�:yz+��D���s�NJ�;☹��?.5"&���ţ�����/�K�ݢ})��z��m�:;A�T[��5	*��iSy\�t��IR��6�.d��ݬ�r���`��Ӆ�F�"%sq,҂'�O;��L�I+��������8���ێTX2�2ۖ Z��V{������0�HdH@�u[��f��H�+pM˯��Zm�U�C^yy�+&�3��>-�(�a�`y;�Jj9Ra0Y�k
���/��{�ǒb9�����L���X�d�
�� V7����s�
�7�p�d�hΗT4j�m�}�Vǖg�5�|���א�ʇ���h���׿^+>V�H0̘8?�K$�� hz͏��Pr��&<�������*��ڸ�_�!��k8�`���MY���,����Rϸ���~zu���ι�������CZ���>����}���;���[���S�ٝ|��l��2��;���2TI>�8a/�6)Ͽ��Mڳ�����Y�7��}��B��Z`5'X~WM��{@�Z�2�ȉ�q��z�r1-n��f��B0��ٿ>��v�Y�qO�wi�l��n�7��ҝ������&�V��*`MP�0�׬@j\pM��w&ҭ��z��\?���e�2��
�1+9�	�x�O�������`?� ���UG�o��Ղh���;]�!�6�H�I��}cI+�p]���`�@���A��h�SH��<�Z�Yr.㟳��;�m��j<�	���X��溷�9�r��&]��p�
2�
��ԧe3���9c]b-�(6$�?�2n�T�4ǜo�w�nyeZ��S�-��~s=�ڮƇ�v���MӻF���ن���s�<	�2!�k��*���Ⱥb=���K�����������m�l�}��UTR�� ����`�Ji���T����¾)�X`|���f�mYV��;GX��o]{�VQM�x����<O띀E+�B�JnZ3��šu�W�����������z
�+��ݜ2QB���+)f&�����$�K�����P�o�fZ,WېV��
𲔒��
��0-Si5Nڲl������P=��?����e� ;�i��ݵK���X�(��裏�
߻قq��W�r+_��q(u�A^7-��a�e��L)T\WƠ:�����t�]�!C�IX��Y�v�����c{�͞a'�F�o��q�_%��%��s���c�TZr��WZ�������!�uAH		d�l_��T4��Y��rnx�[�X�?���ϩ�8g=7��b�Zp�z����u.��-�(�����Re�
5�����P8i��1e��˝����R���w.TD1�G��J`zo<F��)l�S�Z���mJs�m��=���D	}O n��<�-�R��f��$�e�5[�j�3۔�[L<�E�+�i�Ʉ����l]]A��z��*��M�w٧�t� �e��w���("d�0��Z��.d�SV�����x�xq-�L�~�^�:�8k)��.Ӫ��x.�#�Q]�ɐ!�� $��	f��k��ߍ�\˘S�l�Z6Lvs=h9�l�������Ȝ�^�9n�j��k�8	z�U�f�����q���k9�e�	pӥ%�5�~��p�:��UAr8ՂW��״q�M@���6�*4g����ʣ�F��|$���Nr�\-�u�~ɄC�Z�|j?m"���y\��<%OZ�kY��3�0�_W�ؙ��G�U��d�+���/��/��1��+�h�S����}���v�Z�>�:��z�����z�R`����*WKs�_j�������M�\8s�K�� �:w�MS���@��L�U݃2R�ڌsb��oi�S �����+�m	x2i&����1��$ֻ�<Ǆ(�/�CM�ʄA�`K��}G@t���}X����Ņώ�ױ�"���h�$��ː�|���Zؼ�`�fA�}ax �s����ن"��@) 8��%^;n��yk!u��mY��;n���6-�zQ��ʧE.� �z�&��{M��x���_Ip�eZ�U�t;o�*�5F��2�>���`V �1����K�.�J�	Χ��kJ�4�����þ�A|�T <(�#�����qpS���L��%SǶ���:?[�J���'�/��Ы�\K>s�e�pI�+����r��L�L� �!�\��'r�<l	x[�Az8ij�T޿�����N.%�^p����y��	���S��s�p�D�ixZ�Z�JA2�]�v,��7x�{���L`R����;m���FIZ_���ljz�ܥ�!�`ML+��W�QfrF2�0�ΖsS�Y$�f�C�`)�Z�h����ʲ}	��9��s��kve�{���g�P��n�L��2!P���hz(8?��v>������u�@qſ{�wc�O {8h�K��97�������2k!��^9�5-��5�f�UV睤U�s����^�M��w�[�B���f�aq���F@�fuN�2��0wvT�y�G��C�2 �D6�fN�E���:n>��T�>%�zB�r�����-@���>��ώIο�N�}������h�s���.�A�����P����!�Rm8�����^k�����9w�g[zq�Kڸ�1�|��гl�=u�����$	��Ե������������wuBg�_ZZzt��tad��O{Q .R`�(�W��R��%Jm:w1�x��):� θѼ�@"]Ė	�X�.iy��qֲhy)煔�6��?<���kWo��ƺc��fhGRmwZ�2�#��}� i�u�[c)s��\����K���~|�
G�W���jF}�-(=�쳬��2�@+�	X�M��Ϙ��R*dV�HК^�ʟ�  t{a�}Ο|�c-(b\ZV�����䳻C����Ee����
X�Pn��ӷ�n���ǮoK���6��R��� ���=E$y�8��|k�-O Uc�kxD�g*�*W������̯uŗ#W�%s��I�R�|]��W˃��0Д��b(���Z�T��x�E �b{�yN*�c[��"��y�b����&Y�y~�M&R=>Am�C�t�e��n���<)�y�4�w��R2㴄��(.�qX?פ��P��6p�b�s�7�3ߩ�R55L!A}��<���L`�m�S(S�K��!�G�k;2"�t7�jY�����5s�8Ob���8�U�t����d��nD���o��
����L��#3Ƒ^u���)�k��>�ܬ���ղ�w'w�K�YC)�q+�O~r�z��g�ތY��+Ж˷�sBαo�nK ���y���* ą�B� �${
�2yʸp�g呞�������r�՞��� �����:�� ���c_�X�˝�ys|���i�%�v�3��wc�5r��J��f�e�}���|ۏ�Z�����0=�^{��p{���������R���s�m���}�o��),�z��ҵ���|��b��{E���~�g?��q�т�u6�j'X��\B��n�)W�J9`v���Li��:Xn}e|\&����,&>�Z������;x�Z>�V`-���2I'-�)�_iQLnZ��b���x���)�a1�qA�x���k[n+kH�nk�Yy�)���tT&�
`� n�
%�Q[*�����{`���\��Z��zE���S�j���iK>o�p>�e�Z���jq�9O0�����5� w^����%�>�QΗ���Z�I^Z� ����7	��$Ur)�r޳e5kY�k{j>�[�ݱ������0�4�4�@�$��Ynw�w.����u���'cxp�gB�sUϡ�ܓ7=��8�b�ƙ�i��櫆(��R���3\�u4i�������z�)p���:�^���%��kK��Զ������^>sN�zʹ��pe����s�=���o���H4����d�uc+�2��9����P�\k|�{A_&�Uڥ���	�0-yj�Y٠�Nj�N��:�C;@h��"ugݚs|��;j�Z�F� I���s۟�>p�|�
��nZ���w@���̨g�g�!@����9�D3��p�.�m�<�r����Y�����*ԌQv|s���9_3�s��wk��Zs�Z�!]�&�qo_��⇻ OX���
3�qnl�+��0�����d<h�N��e��=�{U��cg[Uvs;j��2���m�$S a?�޳r�*PM�7C:�9Q��Z$ׂ�hXԹ+�e�:�/��m��5�]#i���n�s�5)ǧ�nP;�>�y_��)���ޢK��J%��^���`�b(v*Cm��ʸ��j@���8��� cI�nƪ%ɠ��Ƥ�h���+e8�� ���ua��"���q�b&x�"R8��oZ�7��)���Q���7^�(4����q]�B�GW�ΎeCo�rg'���������9�mU��2^Z{��lZ"��8�� ���&*�r��U�1�̖� d���Z�k[
h��B7L��%�6�~I��Ie�q���KP�h�!������!���	Z���q��9}V�K%��HW~�s ��&������T�z<��e��R�M����~��-0Y�8�Z��II-@1g �ώeZ�3� �=��X�u������������VW ����U��KB򿆍k�ӧ����x�u��u�H��@U9��/��^i�-���}����s��¿\�,ɛ��h"�g�� � �b<`R
���+i�}���˘��8g_ۿ-nZ	[{��}&1*ص�����W޽�Y�9�^C����e��k�(��_�gײs��*&�3�ZW�H��"a�w(�k*R�����8��xZ�`�~�P������L�R���u�oXq)�ŵ���U��[y�T�a�ߪ%��೺U0�d���`5������q�	ps�F�IZFs>�9[-�f~��VfZ6Si�^�<kY���yO77�c<�!)�}�)Y��К��`�&���~SJ��j)8K�5r󷖥.�@~�X�1y�֚p<�a��G���
1�}u.���w�����J1z2\��[�5Ix��9�i�Z�ߜ"�ĸ�ϸ/ w	hܴ�S�{�L���P���A���b���E����Z(d ���Bju^p�����J�I�s��kH��R���ᙏ#���4�ʸW�gj<l�h�-eKf�g\���|i�J�$�62�]�9��rd<�:�t'�k|�3��[�V�oi.�,�-��\Xf�h����ݶ+���C2/�V[���6<A�h)~���V++8�Z }n��9��V2��q�97<6�@A�� X��:���x���M %�HkmZ��N|&��u|��۸SZ��UK'c�垊�3�\�x��$ٯiYNU�s�`3Λ����V���gVǎ;_�m�Z+��� ǩ�o\�;�s��s+̜��Q�=sv�Z �%�@�fN^����u�:��S���o"�	M���$]��T�܎����_��>��0��5�}�g�O�>M�ߺDan�n8Ln8�!4���VJJ˨s���F��9[�h�~K�)�ջ�^�G�6Ve[B~��>[�׆�w	r����oK�ɉ�ר�MM�	�+VK
BJ!��F�NH2d��0��܇D���~��I4#c�m@��-#0}��(���Z�HdB��ָ���֝���C�Ƨۗ���T���p
μO��9�L3-0�{��U��_P-�M�h��YSV�ȷ�l��1O��A�
�����VbC"�.7���� ��#��< 0@�Z�z��o���sxcZi�ʃ���S�j�B_�u<C� k$s/�P�Eڇc U9�R��:9/�W
�?w�@��9�_�qI�7���k�s�+ȩ�#� ��b�QD���ha��s���X��z�X܍�Lp��O�e?c�[��K���ѭ�k�gL�L�*��L������^�h������pk�}�la^��B	��2��(���O���0�e{�w�}H��7�����c���ʼ͒�;ǜ�}x�B�c��H�nr�1E^#_�zxj
t.�ଠ���zǶ���{V��s,9���&���{b��¿Z]�Js�g��]���E=���B�76Q�G``P�LI��{I)�����/��� ��s�7^�Lgxֳh��ɬ1;��9{f-@��C5�zn��H d�Q�'8ƒkù����y���H+��|p�B���k+́���S���4�.�$��8-�Z�j&u�0�f�`0���'����XK���]�����!X٘���Zc�������jZ]�h���r���T
X�*!��峡 �CcO�O3ڳ���u�V5��� �+���� ����y���>r���@w����(K���~vu�]w����p���$�U^��K��g�(r�V��RkP��Z�殽�;(贴2o��;�3ԩ�^��krs`���;���>$nP��|VaJ�iTX{^���𢲗�|��l՘�(�e��OJ����sݴ�_Bs��9+n��c'˄���iY�c8앖XS[�٪��k�~�/��K7C��3.�#(�P�K$��U�:��򰨶�s/{�������Z�=� ���P�՘�)�[�@0���/���Y���o����� S�*Պ�닶�-��]co�"�se"��9/���6i�P��X��6YAkƮq�{��gWO>��a.f !al������5`�:c����|m�
g�@��`�UP��J;�@Զ��A�ϣ@s�z/7@�'��s�*n��c�V�f�_�(�,�-�3�xW <%,T�xv�D˲s�����!X��{�Ԩ��롶���S�Ĩ$���qC�	*�Y.��Z��\�S�ҥ�=�jo�>y��EƱ��<ʺ���Rp/O�����-��x�Ӱ��I��[�\H^+5�ȍ��5�C�"�Ω��+��jͧ�W�����]�Nz�y�rs�]=/i�����k�4eB��\�I��u��6�k��>���[HA�~�(($�堆stæłc�� � ��{{u�Ӌ/�82�tor@�i=���L�#-�9��*%ê$�I���s��M#����1����H��!>s����[c��c[�oA0aM��Ϝ僌�M+X&�WB˙��9��5n�߽7m$�����7�-/BO,���K.���o����+��-��;�311cqUN�n
��y51JWp�Q�W~ޭ��VdnL��9���=P��H���9jI8�b*8�<� k�_|�/V�{n]�P�k��q��v�m�O�ӣe�1LŮ�v�0��CַN�>�������yl�e}ٞ��m���,=cN��c|����Y��1˘q�[*�Uf��0g/됸���g[��Mňu��1�9�=�ֲ���ݸh��<�灪��RPo�|�J���h]k��Z�/��Nўbp�Zj�-�S��)P;d�I4Ō�Z𲦠��|���Ա8�Ъ&�q��=-V��*?>,��|�_�,����կ�~��_׺��,����L�9��6��~�uQ��%��BO���w��d�L2�8ߚX��&��sZ�^5|޳6��\`ir	�}�k��oZ[m_Ɗ����~�O!g&Tq�}I� kZ�i�K/��z��g֖����o]���O��q�����|����oX}�/>�k7%w�2v�L�Y���>O��/cH9Ne����u��ُZA�.�LL�]Ȃ���e�CΙM�q	p��s�T��ɑXd	3�%������6cHh	��J(������cjrT/�3����`-n��%Ш�OY�=�7�����%Y�*�Wu�]��������s��?�����s�C�ˌE|�駟�ox�-�m�n\����Y&�j0�w׺�#�&�/%�5�s�b0O���ދ�\�[��\d
�d ��	%@���e�2��U���{Ͽ)�, 2v���� �"��Ѳ"q����XL��{w���,���=<�}C_mѧ �j]��ә�6�9o��J��y� 4�,KA���t�� �x�t���R�2�:�	��Rk101��M.�BZc��3���s������� ��VZ����9֮}���C�=_��i�O��3�<�Դ�shǠԬ`�>Nak�.`a�q-7�d�/��,�6��W��aٳ,E����#�`�j�w\����^�c�Y#���ki�Ty�T�����%���Ӽ� ��w�u��ƛn\[����9���T�����g��MJDӢ��4�UjR1H3�Q]�K�fk�]z��̚�h�y�3���Ÿes��T��p�ٷ[v�G�YurXs���Jސ�<<��/~�q2�����iH�G+�5�*�7֒���r��I��}��OU��rhւ۲��w�M�Ҏ�60eZ��Z{��dR�ֶ/��ߔ�Z���,pcg�,�)p�ou!ru�����������¹,����� ��~����`7�[!M?�{�j��U����M��ZBI@�	@�^s�
p3�-]�Y"*��2Y���� V�Hs7-@$��L�c�[Za�{o�#�"�#�=pp�2~��5.���j�)}���X@��b��ϯ+��q]��8�c��ɯ�p�5�\KU^����J�k�����J��֘3g����J��2k��hͩ�.�։͒e9WL��myL�������L��C_�bQ�� 7�Q!��=��ŗ�NWx�f�շ�� ��_�z� wN�^�Ew��s���%��9h5,�1I�]�F��P��)�3k����n�>_v5q�9�6}�ҍ��r|�&�R!��VI�|=�V��zk��2+�n��0�T1����v�~�^S紌�y^]�s7�x]n��0N�l歆N5�Z �^Kh�S�N��N�o���'��.��ED�!����ݚe����� ��n���c�=v�]w�uٸ�����կ~u�SO=52��o��]� 	��
r(����F	;V1-��:H�E��Np8&q�P
\�}&��Y�2�QF*h�-�����$d�c���2۟~3�3+x��n��Ly)g.���d�iE�����]�$���UF�>���X<�q�����C��t�W�[�Zc׾N�d�܁���ʺ���x܁ծ��Ω,�&H��"0���2ԥh�
�Z����.C'��|��>�Y[�r��sMy�����eLo@}N�Hy�y��VP��b��@=��b�m5�,9�\�o��|�,_�g�?\�2,��(״q�����0O�=}��G��,@�w����'�x�8��>a}(/LbM�� 7��3�2>\MO�;
z�֨ةEu��dX=gjnn:���ޱَ9<8�y�߫=Re*-�S�aK:�G-rt2�Chh�����T[���9���	H���V�Q�i�%D���X�ܔ@7�@DP��F� `���?��_�⛟���?�L���w��w[X�F�tr�o�=��w�o+h`*"HK�Yr��E�7�X��d%O�o���*+�<ZQ$c�x7OpN�G�_A��u��f�"l�Ib�A	ߙ��4�i۟.�7��*T3l#�V׸Ve@Y�Mְm)��&5���)CO�k ���Vχ/���}� ���:�c�����9��w^k�x��|��B��Tynܶ�Z*#�#�E�����ղV�����LR��
�}��K��׆�`�\<���#t�ߞP�"���#���&�v����94@7��}�Ҕ�o���ng����ܚP*�k��3�O>3G����Rw���Ɗ;�O<���?�ռyqV�I%�>[�6�P��ҞZ�Q�\�&KWӢ9��1-�ۣT`ZXiꞭ���g��d{[����)�O^wQܼ�(l5��Y-�U�]c�Z�u^��^�]�h�4h��2e9�Bm�����
k�
֌[�O��5|�,��`b1yN@I�c]�YM���ġZ�t#�2ɡ
�d��ύ�V�(0���z��𕀺7�s�'�����278�x/���XQ�������O��K]���cVC0"��%
���}���\���2f�ly��#�}���Tq��U��ߟ���>`�f<~h6���>�������0GL6�|�_�H�k��7"��gi�� ��a��&�_�%�%�[�����w��r�N	A\ t�CJ�z)������7Z�MjF|���nj������������-�G�Я��L�'ɵT��5\�c��83�m����=������?����~v/�ĳ2w��d�o��w�{�s�^6dțkW�c Tc��HΩ����|��eB�gS��A��V%}���~��SAҔ�
자��v�}
���U�_ڙ�����we�%�3�T�����#�ܒP�9��'�VÖ�!�����ǧ��|h���O?���SOݫ�����K�v�mH	z�w�� �r:&��1I����' �:����t�fuA^�hUo
�g����<��QZo}�ַP]�d�젴�	�!@�}W�����X5�G�xf�4���Sk��#�ܰ��zr��pW��@Z��^�����9w����'\C�k<���,_���f�c�E���7��&�H��B��i	)�1��jџZ?u|yV,�(�k�����k5�ϝ{�\�x���g|�(�Z_=y�ƈz��Te�^�'S�KR��oᛄz�[�&�o%�9�`��3.;�t��9y���'�~��	r~��-<�SHze�"k�}Ր��?���o��:s����q�i��L>S���)���r��r=����x)in�-�}����M���z�S���j S횲�%���Եe$k��!����K��ٟ�ę��Xd� �?��e���h��=Г����~���?tLgr�s���2@;�c�}�,��]_�)��_��-���\�Ro^Ky���{����9fƇ�̴:U�P��{_۝^ 7n01�.H2K����������ruß]��Ӑ����ZB+�Z�B�1�u�؎��T�Q�S�ۗ�>�E!��ʒ�� ���sZ��ś��\�f�/C�,���W�>�2��c����iM����K��>�1�|9����������Q�'|�P�L³?k8����y�w2��>��koKQz���oN�����;��N�ތ��k���z�riH�dIK�3�p��u��O��Pɛ���'[��ur��[?��O�gG!�er^U*׼�Ϲe(�L����xTE�G���s��a�,�u=������Qە�XJ{1*�9]���|_r��wS��^,���n�{�Gu��=��A�Ow�`�	��ӿY���?_kǸF�=:.0c"�jh�04���>�:@��aў�җ���b:X�� rq��%��M�ƻV͌U��+��4�֘�ja�㟙�i}K���k��6���E�W�P�k��Lfִ�����!w�	��s�\AmF�!$��@:���ܔ$�"/�.��ވ��>C��t��,
���7�0{�#��=V��Tt��p�����h;$��3��9F?zϱ&�׭7���s�4��r�<���OP��4R���Uqr��BIzJY�OUL$׀�	Xo	A��w5�1�1�?s<���b��	K��u9�S=�%�k�ۢ*�Sf�|C�'|�0C�r��q��{�T����n|�bBI�Ço��|�gN|�S��PțӧO��vh������F�7k�
4&4g�s8�hs]��L��<��k(�[4�[��@hOA��T�]s�v�͛ܥ��M���ܖV�Z�y�ڈz�����i�s�R���n=ok����2��e�À`��[w(�|���9�����L.f�50��?�яN|��_�P0�|p�'���xb ��`�t�N�ݿ����Md��ܳ=�EK)���k�Q�P�E�CY�A���|����Z���L�^3��ps�8k4�酙��)�*-��]c�������%	�2�w�)z�B&Q�[U^����ĸ�%e���,e�j�� sMǄV��<���+Я�@�#A�|"������Q�Z��@� X�s0zlZ�]�~_�5	3��w�<w��v��U�ۢ��j=k�s�U�2gtI� e,.�c^C*� ���̜���O~��ҷ�=zr �'�;���7�?����!�08��m�y� ���ʚ��f&ov�^�f7/�4�ZM)w��F*�a���Sϟ�S����$�Ӣ9�5E�!g�G�{�E2�|O-9G��^jjYc�B���M���*��w��dªd=[����:(�ͭTy�5;wץV%�;U�㶆E{�G9q��w����������'�5Ga�U�g������ٳ���M�/��S21�-���K����	p�_�#�U+�m	͚�$PLK�L4�L��_�"���x�Fk��V�/�d.2wpq
X����,��5��0���k��%�|��m1��:���V`^Z^R�P8gk�c�ͭ4yi�ҕ��H�zk��my3�%B3w�cj��TXZ'kۥ)�v��TZ{[Ik�����2�EE���-Jp�b���If��r�2&ۗ}�j/^��/S��@�``�Rj���=kk�ʨ��x���|����'�����
�3oM:e}0��B4���%w�o[��{��1~��q"g �$�����he���	n�����T��k�7�ISރ��U=E�7��z�n���� n�Khj���EK��y��͹���-5N��1	�`<^��,D��`F$����X��
�xw!i�0��$ �9�ck8�䷾�������c:���7���#��H��,�2	�9`
�*��lF��\�Xzs6�},�� �k2�@�ZFXy7�CWrVc`�X��{ZW�����|@,�J�>`깓�J��tk�}�nt�b�7K�8R�AН�Ur���
f�\Ӓ�@݄>}@� �<#�a�&�I�2��w�o�`�5�Ҕ ����^�o�y~�@
'���q�-��=˟9�*���bH��Q�f���*6��z��wc���|�\�V��*1*k>W��c�-�I���O�b�Mz;��j�x����z��h����(E��zmj�7禹�柲����_��S�*��!97X�k�����ߣQe�����N��%oN�:E�������[?�яV����1�%Ç��s�ǲ���,�h�?߱V�w.�*�k��Tګ՛����,�����}[�>G���I��k|�I����]�R�۩I��-K����NY�Xl��9_� cApϤf��[YXn��6���u=P,X�cQr_~��A��7���A�<0�D1��ن�����r�u�ri<�E�G��ι��,HL&�B5���|�%�
x��طb0��2~��fb[Z\[��
$\~�>�� h�%/�-8�̖zJ��u���	BL��,z��0c�㘛$��^k7B��m�7@9s��3�%�wZz��:n���u|�f�xM�a�s�q����A������]�]�)�4�De(�y�v�.����>� Ƌc�>cKH��wZm�}����9{z9��
PU���z}���y���$�N�+�%��:ގm�����Xe�ϱ*Z�:��1��t�׶���a%�ArKx�g����)!?EՂ�)٦j�ޤ�|�X+* k�W��Y�_K*�O����k�/�K��ְ��{�������a��wy�����[üxoę+7\�.�j�>���ܪ����}�z���	oD1���Np�	&�Ĳ����r�*zs��w�1w�\gi�Z+cS7�tA��~�X(;�vL�z�X�ޫG����w~�U���]��ذ8`�,�#W�u=�1�j53{?��P�F8<�c� �>�?�������W�zР��02>} �Y��
bJ�K��� Ra���.�(d������e#-ʎ��?���hsA��x�ג��X�T-�
/ݷ&6Z���r>�ҽ��֘���n��H������j1̾I�[��P^Cx>�C{����gWG������:�f8�R1�5V����~X&IX1	����%�J���g��YR�9�me��;��&4fy2c��$}���Tf��}v��y�92�y�������{��vVo$�6��z�*�\L}��s��R�	�����iɏ
<�}z�J��k�NnSM��!��qW�m?��������=�t{������?��'n����\�J��0�� �큟ǐ�:dmjі7�?�WP>`�ɧ=Np�L�U��My��`���3Ki����}��m�V�N�e���Y=7��V3u�
p��s�j1���<?�Ξ"-t��x����7\�N*��������`����[WW]{��ͷ�ܕ���.����2q�d5]������n�ftr`B'������Lg��P��ӧO�K���e��r�&`�����x3cy�2L0!�.Z�]���T"(кg�pJa�����%��1�\�y����d��y�~����j_���LK} ȵ��Y��G�|f�w^�O�[Vb�ἇ2Da���J	 *@�=�5��88���v�26��l��d�(�L�����j�׵����
�)���r�N@��8�K��*ȝ�:��ڟU
?����x��v�������?/xW��ǩ�0.(ǎǋ��!hP�ʄ6�6A��Ps���q��;?���Q��&Tө�������Z��#BV �ss��K� W��q�9Ny3���pߓ��o�v����3y���[��o�[[n�<���be��� %����56p^-�/AD��*�5/d��ථ�Kn��ޫh[2|�LX.�ނYJ6d	�鵧�s
(�4�t]z��D�@��˽�i��}K[nh�&���!��ʃ�c�n�q\����p1�2�����9�w�!;�ɭ����}���f�#�����/�iМ��p|X�oL�8�
�򤍴��IPWP g��<�fj�*�Ƨ��|ǳki�e�|���<߽�q���-+c�+��-��`��?���} �d>p/�٫�`�C�j�b�B=i�SXIA�IZ��f�+��e���I*+K��֚���
��x�P��s�;���  �@�B�8�@p h�o�mW��=�?�+3�m<����9��e\��ܥ+��	���N�9��^�Z'6�B����5<�P^* v�? ,�*c>�Ռ���׷�~�.儱`l�m�b��?ЖQ9މ�L@�<�ZY���WQdܬ���_K��Tǣʛ�k��n�ʈ���Th�/d��|-�������:�ZG�y�E}����7�|��?|j�a����[n�W�s����a� �(g �(f� �]��S~�Z�kP������2��;z�\�X#uL�]�M�`o����!oX]%S�G-k��C�ڰ����j_�o˭�-\K1�
*�g���e�Y�	m�C���d�#��`��u&0i�tAr5W]���g/q6� D}}`D�@�����=<{|�;0�m\��`���q�MF�u�gI˩`&m0�}/�5��,� C_e��M�WH���N�G�ly�>W���lC�Ģ��,u�glb�d՝��ݵ�\;����k�I���qh�v�7�`���!�9�n}��}]��j��u�Ϛ��Z[
]C-7`�G�Pc��^W!2,�{�FGtaJ�f�AV+�-zT�ꔗ�@���s�:?Z���gK)-R΋�J��Ⱥ ЗZ��6�o�g@)�^��wٗ���H%��M(�V�H eB�W2�	߁��9�ݲ�r�D����:v�ye��u�'O攌�1L�Rc�{ ��^�a����3��z}-��1�VM�
����]y
|�5��M��������y����޺g���FC��s��A�x۶�`�S!��mw雬�-�u���!��9����8��b�`]�k2�b/����f�h'3?���^A�^An
���Ն:I��[-i-�Zے���-���?Ȁ}��R���b��i� ��;2'6��ŵr[V��4+7X�k!�L;�9n`�������cG-{��6,f>Xj��ɜ����tF��p�b�F�k�7�_�O ��]�/c��k��K��>7A�~�dx	.�h��) ����m	̵�ee�:�w��K���\ό���}�W��b:�5�.��V�j��;��qHkr�C�lOZ�k��yN}��6&�JK��� �Y�u� �E��-�ƌE���w����O���u�kx�~遡L@�0���2)--x��$p?�P 4��[-�9O!y��BzG���V�S�#q�� I��Po��	V���op,�2.V��O�ȵT��e���>�z����s�N��U�����ψ|A.��%s�Tdk� ���~�O�q<�9��Ayq�A��&Nw8������p�A�y��xh��)��Y@>>́�*ϯ���AN���y�1�Fk2ʓ���T�]g�X�um]��t�_�1�/���E)4i-�on�\�4���K^V��\�s�~�ȭ����Sz�|��Z�S��[e	��,R���b];0 �/�T HXH0�.U� YLZNl�]��@W�fl�c�=F���n�j����z��Ю�
�^��l�}|��m��e��cb��Cc��1�Y5"-
��Z	��К����	�e�V�rOy˅�u%�#��W�֍]�.-�@�� ����F��y�����t�2n2�-d!x�������K*+� ��Aο֚��Zۜ�Xױ�g�������Na�,y\u�f�fRYe�	�39.�w>��Z�g��:�5)��y�-u��\`�Thr�Q��\N�GB��a�yQZ���˻� ��WTFY��7��!x�_��_����P��fMܜ�~6,�N��a<�w�1���o<Z7[s����H�K]3u�'Ue0��c���ϧ'���,���=�<9C�L0��8���U�m� ڵ�K�	�*��}����~k ���X�Hn����
��S9ge�G�iz�lw���'��9Ν=���$vQ��;/<�º�u˘q%ҜX�ȶx]*���d6e1����z��i?=��vH��-kq}�D�V�ƭ{狅�Bg	�x7F���a��`�h��2%�%\���T�.HH׊�dKO�?=mх�5���ݡ=���JB�{�i�l|�|�]ǲ,o���?2R������ �VE��2��� ��:y!�tC��[�:�ʉ ��3��u׮>z�G��^ �3i��!B2M�\�@i���.�.l�cR�ke����<'�׽�E�u۵��j)���ZT��~��/��g��@�g��$��ͤ�j-ϱȶֱ�ʬ��zו��D*	���l�k�<&?d,u�3��:�_4�[4;�|��>}z]���!"����nK�q]�3� �,/� d�hQ�p{��Q�]Jg>����`�@��[nѤ@���ܵ��Ȼ�9��\�Sי��<����Q`F���f�
"���f-��U�Fc���y�5��r�=�Tx��@�[A�1�Ȧx�F��|��5��yq�[��ך%��2�U���
����Q!|��F#�
��y��������g��Q�P�	�:i��2r���u�=�`���ρ�V#��KJ�,��Վ*�R����5�Sϕ׬.�͌j��$���B��c2��V�V�e���M׈��zH��X��]"�1�N� \��X����xd Y��~MQZ
����sD���&ml�}��
34,�vU��Ը�,�i�������>�qN�dq{����8	�lg�ZB�'뜇2�&�O���,���F�)���Vj���1=�g��Պmgr��˰�k�uS ����)!���}Y�c-G�5��M]rnV��׏	p���m��րv�	JR�̱4vӍ0rM�3�n�?��W�������{FkZZ����̘c��X*q'~p��LH��<�[B��������R鲞��q-�j�vg�f��Ԓ�P４WS�`	�c�9���l#����ߥ���C�dܭ�P1�9�8
����m�Q���I�Vf�w��KO@�v��3� �Q�>қ���oٸ�ϜW��|���5�9�X�k�����g�{��(S�^{���Z�nK ��eoQM�)�{�s �ՎM���zϖ��[���OW7�
�C�X]I3�u�g��W	C�l���B�Zx��j]r�Ba٫L�R(�*@JK���|HWh&9hM�1Y���ZG�d���1�9�=��g)��A|�YưU�dR�1���V�ZL��y�u��j�9�}�������ǻƭU P��S
r�UPA	j�7�WOq1,��V˞�AY�>C�Rp&��d�ܽ-ǔ��(���%�>O+�&����K6ב�ƭ�0	jӕ�u�-�X�����7^_'2+���bYaCσɛ����-��%���U�ٷ9ƹ���c���2=zt\��S& �K�����������L֒�y�9 ����jkH[��w�P�K8@�c�R�~��3��L�
L�����$���,n�����GP���`���C�!��U������p3�������P����m��k)������V��u����~npsa�xS'OK����Aj]��^{{�S!.�C��f˶�~�뮻Ƹ\���]��&˹,:~7�?c�\���dR��$ �k�-���1�������ĥ��/2�3��3�0���یiܢIc�b�Zuzc�����I2�j�2泺� V(3�QD��g�a���X��znřV�^��ᘶ2�-y��P��bL��I���u-牟s�������&rnf_��ls&zL�����P�<v��:����4�q^2��,$ص�amb������x�������;���k��1f�P����`��w�:ǰ�G���Z��c =��;�q��ĴhcJ�%�tN����Թ�=`L�ȳ[���,��O�Vp|�y�Y����;?�f��F��A��P���pz���������X��ζel����Qc��'$zk��P%Xny�.]��A�)�[���6��N���7�봬+-��˰�:-�R�t�6�Z�P��B���vf� HK����?<
 n:, ���\��,����X$]KZ`3�P�h�2�^��U�4e�Y��*()�en�X�p�x��J�.�W^=ߋ���f�r�����ʸ����)E9wm���&&�붯c��Nƌ�'�Ф�YTJ҂�3I&]�2�2� 0#��\�=@����d�E�eb���2��e��]׊1�Z����DU��� �y�u�k�B��1�D�ũ�S^��y����[��4d\nby��ʷ[�'7���Z�]�<�]�K�3��j_�"�f<��E3�]��x�WL��de-�*�y��ђ՛��e_�~-J޷�����:�Y�;�X_ZT�`#o�'�Ғ}���W��|�zS�+2ɹ�ᣮC���'R+Vp�a��,(��%�Ey��Ko�ʲ�3���H>��c<����N;��~a��N0�dT��KA�����u�Z�3��Z�Ni���j�����[V��{��g��Q#��R�#��s��}�PV`��iQ`!Y�_���7}ru��,��eT�Y`Bn����6jM�;�F�#��a�W�+#�l�,�����)%�M��Fol����x�N�HA߸k�qy�+ɔ�"��9����
n�Uxs�`��gl&('�W��[�sR�����׵W�?C*x����v��R(��r�^s#]κ�������N���a��(��݁H�M���H�Y�:�\Z]���s��*���=��9f���%�k-�y�G�=/��O��p�Ü�"���I������V�<��}�k+�e��y�N�/��B3�M@K�]+P����po~���s�V-�Z��Ư���Is�.�@T>Ø p�����S�R7��������s���#׍]��b��X� w���YN׎k9��O��B^Ky����'�e}��yM�R��/6�9s��:��}��o\#��Lz���hn�~� rʜ)��2j�K���juPN�`�۞��gmjuD�>{aD�:R5��ի>o��뱐 ҍbp=/��[�*�����-�޲+��z��u�9���,e��Zl�x�����Q2��ӊ�ڲFk� Gf�������d��'����Znm�c0ES�' ������ؕ�� +JZ�u�2^�\�K�,y�� ]�����{��go�-+��������s8�7��N �貫�S-%��Q�s���X�-!�%�|f�έ��셭��o�B*y�8��š�ٴ�ؾĭX��S��u�3�O𡅩�W/RK��5��ɘK��@f�l)ᄗ��xW�f�z?��׭�~�/�^�3�o����~������q΂��gPOfL���Y�r�@Zx��0'���8w�V{7s�y�|��%�>�oj�L��z�;����?���Q�4}E���]�5�"�
ju��Lg�}o��pE�ZBU�L���y� ��7�X?�!	<�����O���k����~�y~�ϕ�_i��-\U۵oe��0=�㹭�ꄮ�����-�9՞�<sm��[]���j���W]��:������3�����q�!4Y��A/�& �kv;L��R�lnM
Up�Jr��$�H->�0-�Vh�������[n��۟
�xn��#|���-�+�T���޿Ʈn2_[�8F���al�����O h�_ϳo��	��\�*0�n�T8����� ��U��U��5�Gj�f�\��]U�ZA�_~v��@`���P�*�I�H�����8����W*`=n�I	l�e����ݲ$�r�E�n����-^��Y�"�N(�/�l�L,�:� ���g�{Z�j�U���씂b������Aa1�gq�S�ol����Kb����]=��y�}�ř��-��4N���q{2S����%�wi�CP*!CD�3X���sz���}n��Ã	=�����zEfA��P	9�Sq��f�TKA�9/�K��u����x<g�;t��ZY��q]�/��0
s���1֕���y�9Z����oz������9p���^:�["�7�:y�Y���uW`�����֣\T-���-���5�OaP�n�Ԟ�X�_��5��a��4�*~�k�[rm ���0+�Ѹ]^Z����T���grN+�Q�0��dP�x@Y&��Tu�R_���2@��}n��'�J�1\2�[�j��;� �X|
Y�	���	U`<�.n��OfS�W���A*b�^ݹ����Z�|�K�s��h=�I����n��|v^z!�q��X{��cB�\�����:��S�d���ײ��[��ռ�x|��q��K>����l��g�(�� �u��̠P�C��%+��%+���a�A��|�ٹ�aC\��%�Lu�C�g(�c�¢��������qD��*�2��!��j}L�5�}���[��\�S��9y�1ɯA.��v�Zt�͆�2Fw�qǘ�5��N����1.�Ɖ�b��RΧ�P(W�wi��-�c]�!k�f���g,�| ׬�Xnb⺲/�"{��|}	�x^�{\���˛η�c+�	�l]����,�^��?\\
v�L]X{�)|��s=����[���~�4�� �,%�}:��ֵ�z�BK�i�[]����G�d�3L@�uPK� �"�԰Y�Y�[��s���[<]�	P�!��������L~���s����E��&���x��,�#Lw����a�� w��y���Y�"�ı4V�*B骆j�g��O�j�Z�q�����&������K�6�X�����zR�a�YW�2l�����?B��H�?�QA��)�e-t��r���V���9]�V}������U��pMf�_����Z��iaP�0gYkn��W5�6�!�X�e�c�z!��0	��k�6�ֲ�&���(��c�q>���]��;�(�|��?�.f���h� ڻO^�~��mUN��û�D��r�7=5(B�W�3��o��oV_��WWG�=-|o~��F>i�h��v����k��dLDS�͍8���V�p�;=q���L�G����Kkn�)�4��fK�h��z^�ST�ӛ#S�iͯ��)p��9�;�s~wC�\��-Y`S�I��u�S`��y����F�o�3��&\��������%�ж<�`KA�"ĚkR 5.<��f��>c�e+�.H����׍�MZ�h��Z2w)J�+ɰ�+˄����k��0N�; �
��Y�0qf��X$�X*Z��_��00r�s���u|Uw[mW��|ͤ�
p+�m={U<�E;������!������ƉB�l_l<_ZD��E�0���T��*e�����)!���5ֵ�/�:-���$V���c����L�k�lgzN�'���B���1��j+	��������|G��r�3�����"��4!�v�,�kZY-��I}Rz2Z�V���k��������s{��u[m��Ϥ0�M�?��j5�V�i�"sB��XsU2����ի�^�%���cs�k�u��1�7wT������n~³�0�#�6³��d��P�RS���z�/�� Kh�
Um�~�&����Ω��qnopj���Ag��/])�ڔ��UX䱭vy|�<5I��
&��^�u}IF��s!���ed���`�&HutФq��i<.π_��;0�Z�E!��u錖�C�GP����8���Z��:�l�|d2Xu��c��(S�wgܭ��5�dɼ�Q����iQ���X79Κ�*(
�M n����$��ɵ��oYo�p���{��'>3W�c|����U12�`�8膶F� i�o_H�t���X���VL���U!��]�9�;�]O��YGb�k���WMňk���]� ������ Wꭵֳzׅ�zl�de<�s��xnx�p��y�
a*���s�}n|{󻮧� �I->0�{�V�{�J)��5����|�ex4��?��8&x��A�PZ�"lC�5�ů3t���5"o�BO�#��a�����^/@z�	���<^o\/�c��{�g�VA�~�����������\os|3颓�r�6a��߳[��� Z�= � z�Y�Q��{��Rf׺>������Fp���kV���霃"K��k�n��G���XxYC�a�'��wh<.�[�V��XP"�S�v�F�1s�%�˭�a�\�V@�&��~]b�hi�=�	p�s��~�r�����1�� �O �c���֦��w-�i5��uT�[\WY]�*0��<������]�j���6���e�wYȇÎ\udW�x���i>�®p�=�'?�q~�����-j*�d޻�C�(J /�ԲX�(��M[�]�P��,�.[�tU���!�!�u��`ɽ���:Zk5�0AI�>����F��.����_e��M����e=jYgnb� ,r�=:z	ݝ/c_�iz)�Y-���^���E>Z��*z=i�1�L dg���;2�Ry \d(r��3Z2d���|��Z�����-�<�h��k�~OAY���������\l���:Z۸�Z179{ �j�,\cKu��EK�����\�d�H����q��ߴ�ja4�B����2X�k�����4� �28�x��c�-����tȴ�Y	���N���
�*ìc�\u�d�f�R���eȍ����N7c_]u�0kݻZ}EH�TV�s�c�j��y�u3��O&�9�%~�1��f��jY4�o�� l�MMv,8z�3�?�o�?{��lirU箪.I ��ݭ�%���1���;A������_�O�hG8���E�%@��	��T�o�X��Qc����wUu�0w�X{���̜9�ș33��*Ԁ�Ӹ�^�>�t�w�8^gۤ������I�E����̃�}@�q���k��i���6g&�,w`e}��&�G *��)���
�t�-{�=���$��U���Z/!�09�<���ie��,��	zu��}��8��b=��z��q����D�}��95H׬��mt��]jH�S�.��g�>��Vt��H��%4��ފ���->7�oԦ�W�9���nJ���F-W�o�F�����m��>vC!� ���QH}p��Mץ��}]��[���e�c�<��]\o�呺�O>�A�Z�)o$O�������zT�oO�rK��o������������~���*$�u�.=VMF��%�"*�Ƕ�X3�n'�g��\����#�՞��\y�/1? $+������|s���ƣ?�{x,/ �=��(Yf���%`���9�<�h��qXߟ��b��o��Ξ�K�H�������1�g�w' ���AIڳ�Lt��{���y?ۆrH�)���rX� �u��&�Q�P��Y /f&q�2e��E��6�^}������?����c�H{&T�J W�H�t�p�|4j�I��g�pĳ���M�Ϫ�l7��'�Oe��R�#��iE� �r�o�`�4��~���������<2��d�@��>7%��jS{z�2�N�@<����Z@�+Խ�@�؃�����ZY�<x �=�� y�ܶ���p��>��֋� ��d}M�*]ĩ]� ���4`Z���mu�%�"������x���5{���B���u&cLMi�&o��i���eZ^l���#x���2,�����eޖ����#7*��,�}�R�t��%��}���gPLuL���9�����d�`�I�3���	p��dfE��Z�O�4�������ٸ�l/�5�jJ���������M񠓋�X��d�Ds�.�M�=��B��yFa*��`�l/p�z;^����d:4������z7"�1ϐX'�Er��ڀpj�U{�٣kl�y�+oX�Y���ܴ��zJh*�^c��k޶+5ў���ki����-�8�Q8�We�6!P������J}նb� ���BR\�:���G�y�F���Ǩ:�������>��J�1�V8�V"V�ޞE�P���[	�)���Q�I&��W����m�2�� �
���g�(>�I��ٛ�[�y۳-�3z�8���izϒ�&�4e��S�:.��2o�?��k0��ͤ��o��	p�o`�>�rn��`e��K��/�����Ϥ�m2׀��L����m�k(�iR�]
�'�=���7o2�����N���e.�"G�0�~�N�c�H{Y�[F��ܰ�� ػoX�D+;Y�=��i;��2�C�]4�lG�k�����k_�l�K��Qy�T������U��^:�T�	<WL\)���[^��� �VB���{~��U9��2S����d���V*�MR<���yJ�=;�/�����Z/d���<�Fe�1 �G�J�
M[/rp�G��ӆ:�[�e�A����`�*����{�	�4�=���m1�,��`��!�t�-$K��.�]�st{D���L'�#�0$��4�gl������q���f�s�>y��[��2���|o%+�a)|��A �@
==jħg&0��hz�z�٠�&�=����ķ���RKc��UY3��W�Wv��E�1�eϾy��[����X�C˲�Aw��@=w.ѷw?��x^��ln���iP+[��;�����[�x�߫>p	Q�6�~i�)�-��z��Q���Ql�7�J{������{e�Wʔ�Li��&Es�f*�%@��Z���U��yt�A�?rQ�3�Sr��GҎ��z�2M�j{)=�f,���tSN��9��su����%
fO��@�A��Q.B:�'�J�1�I��A���tV|���[��I�e?ʛ�W9A)4�rκ4�@�7c�<+���ꈞj��ObH���gؼ�1>�\�+��/���)���������ʵt�~����{�d�'uê�+�5��a-�ntڎ�u,�m������A#�m�Ф��a?o|�}�:���i�9���Q��%�޿�GV�d�l����Kd{��e�hyn3���Fɷ�@����<�A�s���^�s	�i�/�� o�K^��jJ�J�S)�cOnz��P��<R��K���P�&
��w�2����8Ya��N�خb9��G�M�V�?JG H���ǔ����{���\���V�k�m��*|�`��O����	z�:O��H{��}��5��ޡ��h�WM>���Z9^�;˒���b�����DM����r���{v �Q��Y�g�������^Ƶ�^�A�!r��C���e�l����L�0���8�����\xfM;P���?���$M\���E����#U���SL���B5Q{�E6Ϊn�{��Ϛ�4,;��T>���"O�{[0���M�~5e���20 N%�{#��"X��m����Dɫ4<G��Q���iE�ߗR�{}iO�����n��f����_�W�ևп-oLC��-��ni���o�]��#�@�T��g��#�lҞ׉�[�s�ost�ي��O�x@?�?��Y�Y�u��%��#�Y5���<\���b�
_c蛷���9�?��(o���귷��}��� ��(p��\<�����Q�m�g/y�NZ����i�v51e�[=��[��*���M�f@�Ҟ<D{�-���=�={N�tc������#��eY��VG��}U9M�2y�_�`U�4��I��r`q�V2��_�[������#�]ozH�|���|~�A�eR�8c��k�N�����sw�L��^ѪͲ?�w3lS��~��59�@)�m kJg����q�G�(�_�� ��T�v�}�ٺ������շCd���A��j&�{�\������9�� ���e�R�/mx^o�^���FM�Z�L}�뺢�l7$1����GFG0��3Gf�VZ�)K���'4)���h2(�"k%�$y��q�����
[�<E�w�=��{�f��y�V�h�	�}��w[����O~&E���7����L���_�^=?����^J+�:�I)7�v=H9k��*3y3�=8�!i�w����3��Tꯦk��V��(��'�K���E�Pm���˪nLc���%垞m�U��i�>PVi��;�`��퐑���tg�w��11D�1����Qܣ=;�lƑ��Q,qI~N�}?J�������l �Ѩfӈ���@���R3�SG�-��2�F��� X�ۖ�%#�fy��sEz*!A	;��j�ת�
HxT�}x���V��W�
p�6�i2t��4�:�h9wIɻ� �G&���ie�){�����5�+���a�.����vw��G�[����'�W��H������ {��X~9�v� ��r�% a;8]���˓>�%��uׄ��3{x�����{}�舎o��2�f ��7{�O�յ��֏���?����_������?��ga���H�m >=ی@*�I91ZȬ�dz�0L�y��(lTe9�K�`P����5�:���m�T����Y����Mo%G��v��vb֊�r=bP��6[�.)�
D�Ҟ�դ�R����&^(��r7�#�{R�M!��>�&��~��U�\֌��s,gl6J��Om��?���lz�<��k���ۻ�#z2�3����>3����mE	��&9l:�}r��J^�Fy J�߮��r�j�${;-�o6��2цL}�ϊ�.#e�:u�8�aGioh�f����`�X��^���U�+S�彴�Rk�U)����O���@H7򤟣���.]�U�i�V���H�z�פ ����Ѳf�F�E��t 0&��=����TĹ���
P1�'�����:�5��&��Ev�����5�����lF���\$��R/�dh�~����yqIn˕{Zf>{ "y�E�L�;��<���k�(W�� �A�5�wO�&�x8��AW�;FQ��vo��)/~�#�mQ�K�����B���d9&�{�Qn�})����v�vm�����lz{�[��ýi���B(b���� Żd�$:�,�D��<y-uX���R�����;Q����`���v{:y��J�.�f�[��� �勭��3�ը��]��(Q�(�h���ȴW�����s��";"�������HP�g���@���p]{��W/��|��T�<���)�k n�S�84j 7��viJ�񠥗ys['��G�<nG�5�sD~X>��ir���Q���m�ȓ\�4�@�񠍇���z��#:xs{�G�BЫԕ�)q]��=0�����R����eO�Ԣ�&�0F3ei'}��aҷ|?��ڡ��<���q�}�u��_��>�GF�����;y�+��]LZ;\J��%Pm���ڳ}�/?K�tB�~-P��;�-5^��
���S��Z�9��5���1��E��սkFb��r[^	��s��9
��j�����R>�B��N��|�¤�i��HC���hW������@�N��'��y��𦴲���d&E��{ˮ ���T����g����a�(�i�o��O6r��f�'���m�F��XV>�v���-����#�c.�cޭ���l�|��E��}���O�a,M��ܗ \�����X[ ���w�uZ�����r��'˗�s������_�/i��YS�u�d�Y?��VֵX�G|��f��pX�~#y���J�'��m�X�K���l�#i���w^M��͏�w�f��. ���rܻ��P*�=���h��P?�W�ܖ�j4�'��-	"� L�O
5����6��1����KO6既4@�;�ڿ��G�F��(H*ON]���?<}�;߹�8i `�b�i�]��N�:�n<׌��W26�)��Ϊ����WK�9^S{
�jk�O��ȴ����_��;��/�h�g�|�.!n_o��ꫯn� 6�퓊�m A����Ij��AAWq��w� x����έ�}�id}����2=|2( `;�{����3�������8n�I}���W�r<�����:���m��xu���7NL�}��xc~�&��l%)}�5��#�4-��$/���$ �EP�TX�m��{��-���� �{�&��:H~��}�T}ʗ�u�Lv*�M�Q�v?��!`��m)�I������I��w���mi|hew��.�տ\v�\�{V��L���˒ʹ)���r�+n�fYx��K�����S<�Dl;O�Ji
����˛"�F�6p>tB
�����z�\�.�~���=�=kDm�,��ގ��G�S�)��I����h�A��k�F�=�"�Ȉ�)9]���B�%��>�� ק�٠��g?�>��:]� ���mh]^������K��^�&Hm Wi�I��e�����P�\V�p�n���]�����׹��N�z��k���io��e7�5�W�?|$s�ݔe����Y�$eJv�q�-{�>�ʿ��H�q�Ї1��Cj0���]���u�����8՟�o��qA�j������)�9[E=�ߒ�W^ye�G��.�Ig�#��'o��������f��7Թ��۩�Ϳ��z�EP�y��5�MG �]�ۉ� ����xvnC����t��"��������5p���r\K{�6�n�dy������?��W��� U}dh��E$�(M`���>\@D�"���}#��~+-v+|�A����6o�bmm�L	�N^�4�9M��,3��g N���+==��d�+�z��!|��	n�V\���4�������_a~2����]>���f	��~[)��y
�����)܆�,QF�^�M��X�u��œ�����I�d���;=%��	2댡��� �^Aomȓ���ɽ����{�����!?��=����i�V��d���=S>ڀ��8(Z\>�	,��J7�/1�� �N	�U W��{����я~t>)�z%�p�mo��K���&���f[�0�-��$��d�_�&��L*���z#�Uy�����]4��{���()y0)�=�k�l.����~��ۿ����3����
qկ�5�_J� �S]�6���	�xZ�S��S�m�2Rѓ�a�
�)�4y�6J���.�{�ij���JNO����������������x���}�|��֎o��M�҃KO�.� H��6�ngz�\�ː ������.A4=}��ߩm�-�׿]~�7Y>ն��3���e�m���z�9�� ��˲�1?���<�@2㤧��5�{\�(Xg�����y�a�	�Ӳ�DM��e�~"�'n~K;�H=�O�Co����ȋ�<U����'[?�ig�w����`N�1��.I�鰯�s��+|�}�ݿ���|�ك������}$���m%7u�KFH�M��)�V��5*h 7�?��5����8��y�`��)`�=��5m2�����'?y���xz��׷0�恵"�v4V�V��$�0%��b5pY	�m���y�g��Fi��sf~4c���jO�KO�=]�\����ܰ�	�D��#�6ϒ�u�:�6Nß��=�Z������:�CzP�v����������8� ˼�tq����������`:m�I˲���ǒ^�VWJ�]\^zs]�&��?�.l�\�������9���`���v;Zn�K���ρo���@�ec�/�w?�Ż�����g��&#�F��"�;T�Aփ��X[�(�Ѡ��}�k_�B�<��Ě�_ٙi��k+[����ܥt)Xk �a�	0�V���F{���M�������4�x���/��������u���;��z%P+ʀ�p� �K;����8�aZ�4�6	�����^��y�e��𔮈�HFË���ԗ~t:�6e�鴜�$/�#b�ac@��������F��~?����us�9�<���-�1A樂���n��<]�Al�Z$p��6�m��f�e,$�ה^2<Jy!8k!	�py��a	�?�Yz��9M^R����c��;����<>����&����m����>���ޘ��{�@����N?���mN�>�v���S��%2o���@=A@��/�ڎ2tM�A@�S��{�������/�7>���s����u� A�3g[��Y?7�����F��)�����?}���?���?=��'�.d	�����<ot`e;dz{ z��i�'\�xp��h���6~�.�d��s��w��f�)���H����$�|v��N���]ҪL{�e��l�7�w�I��vʲO�|j�	$�:��s�K#wO���c*��!�ϳ�m�re�Ҥ�����E -j�s�ƷT �m���9��m���Ӻ���[C�lm�2x���c���;����c1���޹.�g�;oN�&��w(#gI��9_,��=�w���@����G�B�i�?�*�i�$?x�\���w+����f+,�[��{x�@���)�����n��g{2Э��>�����^�/SX��ҡ1o���9�� ����a?_�wo���=�6�)�?����$1$���q.�	|_|�b��)����Klz���_n�!�c9���K�ڻF::`8ʣk G�-�p����ƃ��b��#i �=w�|ϋV�r���7>�Ց�s�~�\ضr��4Cv���=!�:JJN@�#�`���)�l*gX��8nی=^i�)I�9e�|Oi�	=��eϝ*i���N0(���r$��`���O��( �`��E9�����S�|YvHN�n���נ� w�4������p�%���=N9�n��S�}��$�	hl�{����kI�4��2��λ�m��s���#��һgϟC�Aǃ�la��ԗ�?pm|y\�)�&���}�unƮ�|�i�tL�ߙ_�S����[H�;Ov�p_�@Ye��3�=�M&��7=-�� ���K n^o�	._�̷��[�\x*�+����}��L�g�C��^~&�uW@3��=+�Mf�_d�^�>����~�L�:��q�y<K��iU���iV�4�w�wRSF6"�ⵠKqYZY+��R+WQNW� !�!�14�6@V��^4�4<%m��uMp�{x'H`�ʼ�K�>x�����-�R��{�n�ô�)�i{��D�����F���=kdu�������icl�k .�h@��	�ғ�U7�>z��j93 j��Y�i���5�-#�Ӝ�g�}x��3��|�X���=|,����fxd��ӓ���r_0�����;7�y���#���yTRy�{23���l�n�߻�w3���*��l�6�aL�Py D���,��:��i�Ʌ�6g	̻���3/+��{9���\{�ےz"�1?9�$^ʩ��s���:�*P�c?ٳ�)wi�&���y`�=��:��6�hyL���4�8Ҧ�Ҕ���M�~�BS;�l*��-��P.�1i�K����`Ls @e��t��8RΩ�T��T������i:z6����/$�4����s��1sJ8�Jާ؛���Y�$z���-��PѨ���S���r�B/s:2��X�Ӥ�Ə2�� x�q����E;{?9����d^ٿR.�]�3�ږ{�dU)�_�`�s@��>���R��/�m`��#�A!w�Ⱦ��%CZ,x�w��<z���r�<n�7��c xn��g�<َ�ZE�o�O>��&��yʞ�
J#=�[�ɴg��0s�]OOˤ,��$.g�y��� :����wn��Z{�c�W4��<�D�\�2���5�G8%��Y�a�����m�m0)#_[�Չy�`��ES����ިh�G�F(���꒴����*RnRl^Q��W��2X���7��rч���p{&h�-�w��Kz7��t9�N[]O��݀Ļ7���ަ)y:)�N�s9�-�y�� �8���	X�	\���m�_�[��K�����b����� 9�{��V����Od5���N����>x��F8$�m����O�o��٦L�}G�z�_��i��������j���[��-=��KGz)�o������y����E�mz8�y��@϶;F�����m�!j�o%�&:	2�!��c)�GmS���x���#��]+��G+�2a�IO滓.ޣU�O۲��6J��d�soS�ջ�Y�����hC��Z�}�6�Q_��C+����#$�x��_ӠV��W*2Bכ1aV�܋�!?cp�D�0Ӌb�͖�;���K}�N�N����,�(ȋ�����-���KP�An�f�Vn9�C]�t����~ַ񐀀��hm����>�0�n�j��64��O��F�"����U�{|_eh�������;�\�����]�6w�9M�Ǵ�q,yR����t=��3����m{?����z�?�e��e��F9f�m.Ruo�����p}�3�L���f<��[����a'�l||4`�0�)`z�/Z����F��d�Bݝ� ۮق6���l��<��z� ՔG�/�Z_�d�`�����43�=:�6�}��lmdvH?w[�I��O3�m��2���c�+��i�I(�t�lVϷ���(�K���}h��X?��n����s���������ļ9��c"���������N/=9�^\Gz/���{�&�$��E��rˮ4��T0AZ6r  � �eu��������K������e��߀��o���d?ӷ�z�l�}�+�_�g���<ah�y��(��1=���(�~��f�Dy(�O���L� ޲�v�N"~�`Ġ�2���˜3�#Ӊ��3���7���>l��8(m�����<̂9�#�gymO�A�6�k�.+`���r�?l������Z���|��?r��y�����}r�'m ��}�v)������i �i�u������[�~��M�V�5~M��H�t�祴�� Q�>���׮��M��=�y4�I��sG�\���;�ˎwɨ���k������A��@�M���y��� ��������B��{V�4��V��V{/*o+n=c��m�n������R�j%�gԵ`N���������	J��ӻm0�;-�3�E�b��{~Ҩ8l���:-�g@�S�����O��n ��Ѷ,4Y�>cmX�����CVH��+�� o� ��c%	����ӷg���ĳ�d_�m�T.����<��u�W��'O��GH�����;�du����r
�'��ٿ	TS�$x�� �R��]�?��m:-m2��U�ou�rgzLs�A����>��r�ʐ������7&�I�u�=�rM��:_�{js�k������gy����̓}_�|�vWtĞ7Y��XW<��<R��ε|n����6*JE0	�ߡ�kʛ�+�����D���?}OJ��mEm���m�t�Nﬞ���q����;)�<Y7�����l;��3x�pO��_���<l�����7C�u���Y�*����gxp�7���>��%���������iq�ԇQ�l���}v�~�>�-���7x���54�e� �߱a����w������ݶ	Z��� $)9��þI@C@�����1��Gi���1���a![���c��RdPoyR�._\�<! c�8����"�Y+�|\'��6�y����NSe�@S�R����l��A�K�z)�	)_�a?��h(_y�I�6\���|�K�(�J�i� �f{.��l����>rW:�W�m�9c��w#�������v��i ��p�;�����y��N�N�;ʫkh�켿�SǴwa���I��Cv�%��$�#��W�m5Ri���'G��)����{�e���(G�GGeV����JQ�c@O ����7��7�<�������?���pP�/`'E�o�-P���|g{��͠C���p�����wߣWF �� ֪�4�6����w\����������g��O���-�ԫ���m#�O�˸����e�(TN����,g遢~�'��PGe\u�O�N�fn��0=�!ȴn ��7����0�7��a/~� �r�S��%�����J�P/�Cϧ�$��ݓ����~�y���}y|����w��ݭ_s� W^`n��d�5�2�-<(�'cɳ8��(���ܤɎR��#��fK�ۨ٬)}�K��x�Uj~�7~c��t7�����o���t�^B���sRe9���3���E�FS��O�K�ё��i��lyQ���-�$PM�܉X�i����
~R ,۞Hj#��!�Nɏ�m�W�)�#�m�ڂ��(*��� ە�����V���7�؀�<@���kkϭOJ�G^ۿ���9�<x��^��ƍ �@��2�`{�d�������Ώ|�#Y4��;(-�f�+�����;�Dx
�C}�W���dz.=;i��y���E]�3�F��4���S������<si�]���q�bfS���ј'lW��2;�[����Ӗ��,4�@���mz������[�i�A��g�t��w�U�_��?���+��8P�(oMFD�eO�s�D Oǃ?�bSN2��S�4��tv��#`��j�l����֭LI��J�Y0|��o�� j*g^K�rp�G�k��H��>��h�C�ʮ7L�a�
pW *E!&m�<��ƭ�������4J��x�c*���nJ/�ux����QPRk/�����l$���(�R�G���:���@�<���r�����و����R����u�5E����6�S��?����K�T����t�q�m:��~��i�1��\��]�̾���흞,�w�T{h�O��E9O9���1��$s�6=�����F֐�v����20h�j�$�Wz�	��,��ۋ@	��1|D�0�*LA� �k�8���I��k/�� P}�\���AF�ˤ�h�"r<�� �E��߭��|��f��;=�y���d]�	�gh�ʦ2=�/ҕ�]�i]. �Aw��6��N_ޠ��Q�.��S�W��Y�
+ܖV6��L�6E0ux�$$����n��F�y|Z�l�֑F����4�V��UǹM:�w�w�dj��1\\|&j����Ӱ�:s��b������⷏ׁ۔�b�4�"��_)G�o�^.�����AA�j}[�3d���Z����ӌōiq�T���&�r���WeI^������2K�)e9�$8��U�YO�v�����r�G�co�C4H�W�\�PгLޚg�1^�Q�D,�J?6 ��4Vvd���2��"a?M]q�V�|ff���L
u�wU��5(Qh�t�N%��g>s��yf��y��S߻k��J4�y�%�?�t��m`y�4/�Ob�	W��p�3V�
�5l�V��Z�U�&���3���ɤ6:^��#���.:�*�&0�z{�'�X.��ڛ��8o\{�<M/+��S�$�hu��}�����C�C�w8U��N;��W}�����u��t�Ӟ4]�v���.=����ju�V��L��:�|���'&�q�U����yr���l�Sw�,[Y��o��/��m���G���\{���gR��f�P- �bJ\��v�2x�A��?2n��:+Mz��m���+�5щ�-�����.�zw���Փ��k�7~ރ����T��D� �F�N�������M3��]��gQ��R��#�'X0����fqVt��=	��(c�� �=Rv�k SRƧ2��G�ۨ)��R��"�26�a]ZP8Z�M��<]�9	�A^*�3{m��%:.r  f�`z	H'��:�cC<y���FO"����8k�i���y������*��Ծn{.�r���$����y�%���H��S��1��`�^�m�~8��� ���o�Ο����ړih�?�1d:��m��o3#/=�>����6�N{xs�eo����x�,�J_R�5]캥'<���x�%����:�x�S'��:q5���:�Á�ی�����q����{Vg�7�>x|�ݕ��@��;Ҟӽ��]�Y����0o��Z�Ų�t�ěK��T��>�����p�'�Fe6��V�oƛ�9�.��׀�,��V���W�in�v�F�t��"� N>�WO{��ܧ�����J��4�Kp+J�b HJ �������"A둀�&C�-�r.k�8ڋH �@n�����hz�3��e'�tWJm�g����NL�|��0�괌�β�w�CLz�]�bN��1�t+�۠�ir�8~��ʖQ��E�NϞ]�L�����7Bf(+�����v�'�B�1�Ӭ
yb�n���۞3_\�������ʨ'�I���ȲS��X�	��{9�i6�}���1���Lh��b���/����/�tT'�!��
�ʵgw�_��o[�#�����%Xm�}��V-�z����ן��QS�xc�^����6nk��U���*��?�ݪ|T�����ܾ7��K�H'l�����m��߫�i��+D�ڦv'�i׭XYfƆ��'ț���N���}�y��3�l�/4��q;��l����������J�Ķg�_��'�'����&H�ן����:4fȊc�ڸ��yg�	��o/4:�Y�8����ȫ���}r.����	���0�s��<��2e��d;7y���mf}�
����e��	ص��V *���O.r�N���K��>�{���z�@�/hm�tb����5Ƚ���Qk��*��}o�7?��t�s��ī|oU�=p����S�����t���9|��yJ���^ޛ�ٻ~T���o.|���'p�<���?���|o�r,�n&��e}���k�C�E��x�ɛ��К��:8�%�b�Z�,oF��|ۀ��8��`8i�Ә�A���2��[Y�=Ym�c���y�Yz̩����!�jq�9mk��=��}��mO�lcQ;ɌS�L���g��v�����G/���| C��0M/<����5�����ږaB9�l����~�^�����9hq�ٿ�w<�ۋYｏgv:�֖|o}J��o���g�Ә ���8 cT���1�q��A��﹬\�ɓ����m�\�vtZ��k���t����笞9r����t�
�U���g��p4tO��N����d�R�ќmx�0wOh�J�B�t�o�kƐ���5e��#% ��*on�Oc���i������e����#�iH�0���|9��{�]����)���8��4^�B�,�k<k�� ��'ˡ��Ƶ���Z�n�κ�6�r���m�|��n��L}���e%1ߙ��}����D�^� �L�.�u�p	~S^X�k���'�1��홋���>���a��M@�@ۗ�U���:��u~���������p��<�����J9���r7�ƫs������m��~;�LoA���e)|L����P�
u�g(����g�5�?�ҳ�?����taK����64�����&���6��i��H�}[�ކV#�drk���$yH�Q�%�����4 �����<[Y��)��v�|o��U��������R�1�����	b;�f2f�"���v����I`l�&o�L�!��2v�/8�LH���f�[�~4e���0�=����.��5��`*g��@�(	���$0t��1������g������s�ϳ�u���ַ�X�6v_���2��y�^�/��>|we8��qP༩�W�H��5��&�پ+�� �$��+���-�����H{���_����:��z� ��������σ	��"���=J�pD>Z����ջ������,�b�D-�/Z���+�k�'){򯍈	��<���7�R��5�q��.����aEgO��dNkrJ<�h�6�rpP�)7?��3^X���_zF�E��'���W��3Y��[c�@NiL}6eu[��nH�:��"���<J��v"���X�����-ߛ�q���fl�ۉ����eH��<�}Y�I^H��s��2�����m �����y�r5�����fh���K�L��İ�&�^�T�[��J'������'0��Z}T��-u�eo[T���y�,`����dç�9m��Bw>����Qz�uL�!�i���<1�hZ8��=ٺLv#��J�=��=R�V+�6����٫�%LZ1?��q:�	ZR��QA��O0F�앪�$@��%5 x�@c�6 j!�Pe7����h@��l'�������⳹`��g{e��W�J!���6@`�L����ɲ��h2~�h�0��x�3?zsG��)�g>�Y6=�Y�	�O��r�6�����O�e����T��i+�|	Q�{N�<𴹾���w>�9u�S�xd��:�lS�m�헔�&c;�W�������60X�s^O��.��䌖�b� Z���u�!
���QA�>h�kZ9>L �4a�#����$Oהi��Ю�Lsdۭb,�%�>��J��Dǎ.*��&���0������h�J�����N���>EK�@#�\)�`��N����2y��q�޲fZ}=)ԽQ�t��<li7&���+��>���n�P�3��Tn���)f{R:��'_�u�Nc�Ӝ�Jۃ�Iĩ6�'6��g�����϶�)�)mQ�n��K�@��)d�����mS�ɣLϠ���!�a
�iy�>�z��t	s�ƶ�b�����Sh�!uC�s���q�<EP��o����n����4Hg?S^Mp�Q���40a�e'۱�6�;�SF�;�*��p��E-mn�Ɓ��M�O�;H�]ú��?����>��Om 7�X�\�"'0�� h��핵�/�]c���'1����iP5ٔ�|�s��e��|�y��k����6œ��������:��LM�����P6���D�Ӂ�g��ql�7��F��@�4m�CP.XaYר�0uj�O�ts4�B�|;~y/y���:��x'����~���O~�Gg>p�!��%�d�
Ҁ� zёy��M�ɀ;|"���r��2�B�����N�h�v�\�L`D�J@ۀp+��z��3匡5� qս�<����N�7?�OyJpǸo�?�1�6k�2����!)7�u	���V�oʶ5�pˣ�Y�ԕ����U\9o�-���Oڛ��A�G�9˵j?�qp�u%oZ�g{�{���2����3+	,�nM�rZn����m�>�[��BH˱�����?�������r&��-m�C#�����>��G�Y��<ʋ=���M�����3�����Ä����Y�ncđ���	���]�7�u��^H! ��O���k�m���ب3*�L�Ϥ�i���-� `��o��x�ӷ���������H�O`h���_�Y�~�ug�����}��WN�����Vn+��6lzp�NB�/�}ڢ#���t��0��h��T_�'߳A�vl�i�0#�Y�+����>O	²���=':�|���%wkI���Y$���	��m�˼~����.�Z9��M�r �ژ�cpI~q��u��M��������_�?��0.ejZT�2H]��|��G�<c���9�����lS�ܥ��|�<���	�1�-�Ȥ��c�α��o+Ç�.�����K���t/�����̻���ڝ6f�����8.3pi���_�(\ڨ�ФT�3��ڳ��/�������G��	�ٛ�x�,�$�Tz��慶n��w������~��Ʒ�8���?>�$�m���cz���&���	p�)���ꫯn|b���E	������Q�-��Л�k�̋��A��s�r�p�Wj2�I+�4���6-����:��5`O��(�e]\.OWg�Q�{
��x`��.7�����M0��w���S�#�[Uz�	�L�pB��;u��$?9@� �aO�����۰y��e!�Z�ݧ�w�S�1ܗ9e��6�XNѳ�W\�[���Ȝ�J���4A9ۦ�ـ;y���@.��!j_�'�H����f����@��@ז�.l��I�' yD���{�Y=w3^����x`B�TJ��n�dz�`E�b���:�=�zV���^;��o������w��W�zz�嗟�՜@m��,���w�\��Iy��#p��~��'�'������bH����T��H��]�4ʛ��|���J��"�0p��ǆxS������3�|�y<|���'��M2� ����� �c�2��C���(�6:O��r<�i������z�>�����_�m���e�^�Rƿf��}~�N.�s������M��?��y���'�iG
�Sr��N��?7c˙�Y.OO .� ��,�O�����V�ŃT��g;p`mGy��2���dxF�d�y��<�o����-�0&@��h�=� �*;38H]Q�K���l�K$�?�Aix;0(dO�豬�����	�n�y!����`!��0Q����h�Q��f����,L�X�k9{*D���{�����z��^'�ce��- ����򕯜����۷H��,ٛH/ː
;�kP�79m)�F|�K_ڀ��������-�_����g�(�������cy�K���hS�n�4F��������z ^���������H�U�,ۉy$��7���H~��+yĴ�����w����"˲�֧��������Ә��#\*CO����cpŴ�[z�Z�%/���6�3*�����OY�v'� (ny�m�63]��z`+��d�z��s�S�'�:~SO� �G�K�ʧ�A��u��ų*��$�5�68�~��{5�a��19m�z!y0���q��mN>Mz�y��-f�a�=�~r#��Z�V� g <�e���[/��rK��9�[��s��>[�٣���a'��SNN�*]��>l�z`z��6����<�iX�4R{��.io�A��L�JH�Y@���^�@��������x������/A�A��J�K���=���w�`�x����x[�f��:�^�Ϣ}V#0�P'-B��Ye�=o)�|i�3]����tk�{m���ʡ�)���p��p�C*�4R	H������(=_܏������V.�ʛ���qI�.�ǜ��B�4��(��t������}S�j!D	���0'OVéӵ�w{��f�o�g=&�C�&�mϮ��)����t?b]\�9b�z�eyu�9�[����r��T�a~ts�e�"Q>9�͙���0��l5[#�����[��2� G�wu��<�	nE���q����K9�&�=��P]dF�xD^J0�k��w�RI0NNZS-����{�����o W^\�
��P+ZQƗ�xהQ3��_iz;+)��|�3��B����7��}+_�ShC��Q�lJ�h�Р{+�RS������^�)�̋���+%+��v�U;�o�ߊ^�6c��H�[��mGO��%X^������镢ik�G��d;t7�EM����n�)=��N1ϣ� )��e�Ө���A����<b���bp3v����O_k1���P���đ�=�o:�`���0�ˀƱ��EX�Z�r����N��`��l��zP�j��A[���rq�ppf80i!��od���/{z%���1����oO�v�:��v��|�֋C�X`��l���/����ezϒ���.J[�,�sW���w�������`���u����n���GR�ĢѨ�~��~��ۿ��[|�W��I���tZi��Tv����B���Q{�P��9)}�P8.J���g�g��1���ɇ� �J(i�ْ+-�Ֆg	6Y.N�H�zO�U��}\_�{Ε/��Y�� ����Nk�����]s��:�TKgOM��4]z�H���	�َ~O��S�l(W�x��T�0y�{Em�T�E�mڴ�)�9�%o[��?��$뿢Ps�x��-c�dp��0�Z�j�+�c�k����g�g�Y��*-�ZY�<H�@��4�ZX��i@��>����=�Tn�������S$�ϔ?���s�q:�[��Dq\m&-r^x6�:�g,/>P�}��"����hj}8�v�
����i�.�הc/�	`�7��(�<�:�M9{ƪ]���P��qh�<�T�ܶ��k�/~��o��v�qh�f}�A�'p��.Szr�XHy���믟�Vj����gO.�SN�7�7b'L�����Sǐ2/	�rq��n"���.��
�� JN�/Dy��@��O�@c���H���egl��*F�}��\Pؼ�4�SZ+`ݞm�F�3�����R?ػc���CbZQv�;���M�}�i�T��I�.�R7@�t��g��6�b��)��>0�Y/��i��Q>���ɿ�=O�{m���fȆC��[V������4��ͧ&S��k��|\���}�w��N���:y��>eG�xfϭ�E�H��y���zG`���*&��||��E�J���}������`�e9V��0h+_�Ea5bl�^[ѣ�\K�\E�����i�$|���<��4�~�\��+��eN�@�@XY��`��3.�p���/��R�hᙽ�6���Q�E�Q�#�Y��8X�����o��P��+�_�q$jNY����g^&��l��@0��)��b^�f-���cYڽV��&;񀀰��Օ�͞�\tu����׋�D4��(cBY�6��d�Ϻ/6��g���Kk�kh�Lu��Hq�z��zO��`ٱ���rٖ��'���]{	��g�r���f�h!��`���s{��4����� 6�3ۜ}8ue�M}�6
�R��h�h�Z9'�==������k��a�����ϟ�{�jz�.�ܖ�%�m�rJ��@�w��/}i;�E`��X5�a�c%�)(��nA8-%?�k�m��4*a��<�~�������O?��O���e��^¿y��5A~;�-�Ӕ��������}�Ƃ>z$�?�N�"�	D��M,�ێ1�N7y���<�Q�;S���'0������iP�3�a˱>�恟�'/1��:�\y�`����~���g��L�ڥ�V��}����`co��M\W���}��H�=�d�#�kgZ���-xRڹ����90�����f$X�G�˽6������hS��&�9���ݖn;&m���g�8�[#�_��E�]�aJ�M{xpOǼh�pW��|)��m!V��Ɨ�dϰ7C�N*�b��V1���;����)K�4����6�͜W����3V4�����G9���m��8�%�Xx�\��v�e���a;L�h�y����������6�^���c���0�Z;4%���sJz2~@m�4])�f��Z?��?i��M`�x��'\��4���:8-z�L�����]J�k����CО���(��r�2�'�m�{�gN~S�=T�f�K���r0(�m!��$�)g\��e;�7]`������~y�e��+m�����{�3=�~�vQǺ��_9��6E�ur����\�0��V�A{:�(��>{��_���wj^�#� N�����n^[���W-{�^1��L�V�[]M�{�͊��ѝ١�R�ц�=�� �^A)�l��q��kfe�w�y�}��)]m˥�\����K;��W��v4�������ƛg������^���o�+�Vy�=Z�M�&JՀ~�Ŋ�+#��V�tG��l��)^���^���rk�L� y�����)F���D��i���}p�ũO����l�_S��z���Yo�ID���)e���0 �� ���`���~���c��9����g�o�-y�@�ޠ&�'/�Z�ᴓM[���x�V�����$	n�?yM��m�C�D���&0O���W�����#ϑ������F{��Ч�s��N��/f��H�e|��M��ny�wTw@y^{�������m??���N4f��^H�K������VG.ts`����ɻ,�O�G�����hP��3JO[�yꏊ-��%�Lߋ�����V2FXdcg����G��^zp3D`k�w�=��_l�iW��;��@`Ce|�R�������Q��ʴN+��V��l�i��^�1�=5/!���k ����o��g>�����w���Ɨrlb� ��d{���s���W��]/�7yx��K7º��gn�o�t��ƃ��zf�P�{������ j*c�1��f��>\�g�}��~�;�����`���E�,��0ɔ~���
r'�{帄�ٯ��Gb�{`t�n3�){�d�>ӴIJU`V;���M�K�z�����g��~���� ����)]R��V�(-�+E�r�H`Ƕ�@+��m W+�� ���*���G��ZX�L9(�޴�h@�&�4���q���>����IЩ\6��	Y)�v��I~�he�t$hN�׀y -��t�Qfj�#�ۃ��RӋ�t�f̓��Jޤ�_�(��5�����G�޵}5y˼�8(���r��	p��vQ�O��B�I}�m�-�|���=t�D/q�{����	��+M�{���d����+�8��ЅV��pP��:$��~��	������n#�T |-]R�����cb>u>���0��g�m���=�*OuJ풠�Y�� ysE��v��f�9�����������8����?O?��N?���)6���޺畩JW�������[��@h�[�v\�<%��W�B�ё�WeU::`A����&a��V|7�l��x����I���L��^XD��z�xJS�u[�D^%��ۤ�(�+ş���Z)�ij��o����r�a�d]2��@��1�\�<�ԩ��ۘ��ʝ�Z]��&��E���1�U٦��05�-�[�M� �m�6�5�"�\ʥ���{�z�����3`^��M���=��jql�_�j��\�eh}me�[�i}�my������_�g�c=��E]�Bh=kG�t9C���nwC �5��]���=Hޭ��J��0��[ݟ����ki��#����p����Grb~vRD��Nʧ	ߙ�J#ǀ�#
d	�z�>{m���;����g?;}��<����vT�@�@*�1b���MC����-���v@�T�vxx�_�r���?���|��>2��f�f��������o��o7 nCs��e��u׷�$���#ϴ�Уgp˸MN�:/+M�gz~�x�1_�Ȟ@n���X-s�^gxƔ6�n1�i\	�Φ��g���!p�n$.��zҳ�@��D{|g��5n���|&�5X�l�ULf�\�௵��#�y��r-J��v�.�~�~�a
>�ihQ���?��?�4��&�v�texxd}��>�1o�hnV2Ǻ��fKL�0�^�A��n)���O���Cm%p+Ͻt��mnˁB���3�����q)]��z~U�)�U�Z�G�p)��U>�L���ͻ 7�)=_�� {�<�HƵ��a��6Z�:��h2"{D��o���� @*�h��i�,��g�3���������6 h������1��Or9p:�������o����ID\@g^�6�����Ӄ�<������^�اQ�������JY�H$8n�� r��v_y��x���.��ǝ��,A����[�d�J�<��ߊ�>�2,c�( &8h�0��z�;�4ݜyMe�}���B@���G}���b���Q\�.$hˁ����ԯ�@KǼne��m�e;
��nb9\��7������ײ��F�d�V��K��5�I����V/�me�.��n-�m舎y^�:g�[��~����m�]VZ>\g�g &��
��g�{ʓ��kj\�qjZ�Ɩ�����t����O�����}m�l��&���C�<�� 5*��?���:���
�ö`G��U�������f����>n��-=6PT������uˎ�:���]y~2���5Y_�iʗ�����q��Z1�϶���J{�`�@��\�´,/������{	T�xL�_c�2��Rz��Gdy�;]����$�jƪ�v+���tn@��#Y�w����t��p�l�=��{�?���cٳ<S��L^Z�,i���Nh^Z�Zz��k_�R�:jV�I���)̟��Kl�J�W�ۻ{�&!ה��Fה��&~��S�N�5��2g{��DW�#h������;+@�g������f*@5���n幕gU W`W�ʫڌ�l�r���74ͧ��������2mk&��<����=#^�a�� ��,�F>ݖ�1Mŝ
����k��!i���ަ��,�$W�;�z�v�K�l�|��ʨ�U�c��u�ӵxhu���n�g�xF�rA�J�L���g,fXP��	����;�d#?T�Y߉V���L�4 O���:���Ϛ!s��h���2 ��r3�$�M��$�m�;񏼠������~�,�����Q�ktw���o�=��G=���;v�������N�ä_�v\Zϻ�۔�F�O��Kh��>K��ԁ�!�qk�;Q%N�h��(QI�"�ouD[Ťj��n*D�g�X�7�|����}�Z��N�R�H��x`1�@��ڊ̊A�t(����/o�yq�����=���	$�%� ��  �� Wƀ�x�x��nҞ��3�����W^GR���\��D䮞]���Z���F|��Y�)cphmH��tK��>Y��g%�y��|''G��:��I�LpJ�����gy��g��{�4�/8�D֫ՙe#hf��O@�7�h�Oqf!AB��Sֳ�=��c�/�X����m���\e�|�(���s��vgc��Lt :�������Zp���W�~�|��F4�Rxr4�`�1�=�3,9<A ������;��ki�}-"S���n��o�f��õ�)��c�������m!/��^�Š}�88l�ۗyO�e�wM�����s���iL��P�yn��,W�yz��V���9��	��6b�����'�[yy���2����Jq1���v*��l��l��/�-<jed���e�	b�<�D JOaK/��gZ�F���){y����v������<��It)���߫�Ͷ�d2ߝd�魜e#�Z�o�bz��!�~k�f/�)�K�`o��,*�wN�d�t3V�<b���u�4�`��ʷG��R���sd�7�"�l�E:�#���H�s����7����%�Z�.'&(���!�����2�/�(��x[�u�Mͽ2�*+�� 5%ȼ����(hK2yr�Tv]���q��jyZP�jA���ջ>S�YӤ�E�Ҟ����BZک�lm_�����9�6U?��i@��ڧ)pG�h�f�a+�"����&�����ͩ^	n	ʎ�7�%`a��L�����k�g�mA�ʁ��m����[̇@#�=�M��r'�g�f�7�1�K���t8�{�	l��km:������c�w�l���tD�����[d?<����=7�a)������g�km׵8d����J\�_M��w��k�M��wt����F�|��Aa:���m�^J�L{3�9W�x�� �@���ޥw��d]'�nJ�Շ�^�|H�w�����_�kS"�	־���꣐)![q���˿� .���xW#�����{��m�ƾ��� ���1Ԋ=��n�g�vz��@�\��F&�ڋS�+'H�GyoF�=���x��~j�Vߕ��ܚ��B��<���)	4�:�u�]3��-ߟ�J��eNyI���L�m`N�M����O ��s � ���B�&�]�Z��>����{�d�<�dt�+�>��w��,�J��ݓ��3�)����zR��B/�΁��m:��΍�We��������u٦w���	l���6��YХ��Gn�[�(\�ⳓSP��3���7�{ZL�K�T�O@Uq����=k3�C�R;(�}��%�i�	�fک�Z}�P�T^r�?������g�gۂ9V��k�m�*�B(+��������@���S;��o�P�����$��b��}缨����o��֍�I���q�l��
��g���t	��5�d�_�O9@�k����K�5`� ��P�[;�#�9���.�;��.YF湒�̣��Ɠ�oϧ�H��3dٷ2�L�m��+����v˹ ��&0����#�D����z	3��{���{��s������|�)e���������/mu ��\�>>��#��Gp��\�7G����YnK+���.��j����6c=={4M��!�������@���&�|�\�~t��#y�-� �-��@����*�X�P�?��??}����<�S���l���TN�{2���1o%����I���ez�&�%�Zu�D��
H�t�M�� ��3��ƻ�F9@�w� ͭ.��|M��L+�ߌZ�xN���A��T���)��[�{�o��O��bĳ-���|ym��t���59�"����<�8;�<]�֎���g�h|jײ��X��,�d���%�.��l.Ν�H�y��<������ͻ{:f�Z�Y��+�.���QZٌ3�h ��O�z�O�ҿ��*�$���Z
v�(�t|�����o�X��}[y0�ԁW
�����iL}ʗ����ծ�H�.:�B��U���5�k1�i�������ȗ�:.{
rݎ��>����%�9�H��o�*�Lyj x�K�r�8��~0VR�	<��,���{i@o�Hhd��u�@�^�Eu	�H��K���{�2.���9�0��q�� N'[�f{�=��;����S��`�}wJ3mJ���������M�2����3�g���p�� {��)+ɓV'l�����=j[��ݻo7�=�r���] �Km؇�~�a����%t+�(A�4������\d�G���i2�,��ˋ��]Z���i��>�P� :��bV�)��A��R,���������j��V�N ;���P��iFd��=��y�E�>�C�}�u���񠢕G��6`Mʮ�t��͓���4�39���L�}9����K���q�.�w_����&�'^�k{�g��]�x����4��=�ռ���z�zm����XI�����1,/������.��l}e�[;P��O�}���җ��e;
�2-���IߐVvy�O�������sr�>��Pă��g%/	���\��]n����gN���o��e�[���{5�=B���yq!G���6�7C�1�U���� �����Jk�Xq'9�l���ޓ!�r���iDmC���ܺ�S�媳Q�����
4�ܪ���ZX��孖B5�y���.����T�'�:�^�f�s0A@Õ�G:�ӟ�0�p�Ńx����Moy�!���m˗�]�Y6>M��r�����ו��6I��� KYc���)�l_��9�����鹿Y�P���峺&p��R��=�K��.�om��|��ʹZxD��VG��R����nz��G���� 4e�i4���<w[�{��g��9f�d���BwG�/M2��G�����5��'#Ӟk�y\:�K���V�Ǟ_P�^��S��:���i�*@�S8[��F+�{e|��yt�˦�|l�>���!{�k|e�f�N�L#'�l�0��%[�ß3�F���f���3f{u�^�?�`#���|p��ڂ����w�~��x@�h�X�?P�����J^P��3RL�m��o�cR&�P��?gݧ0���Z��h��`f�`ɲ�=n`�m�j�Y�	X:m�l�>n�6��q�E>��2H�'��L�������k 7yp��>?��[=K�:t�'��@���9&���+j������z��p������&}� /�5��8�JSX6~T$�t�O�mn2v\��pܫ7����:aL^\N�qz�ȨcE9e��lT������={}�P��ה�d�}�n`3�1����Ԙ>�g��'�M�o�cj��M���3������o`�<�����s ��`l6A�'���'xn�/�g��ne"�iuj`���HP���k�7�����<��g�N��z�mp�\���,��G��-Nd=j,#��&�����a���^�r*��<���@O�����
��=��?��� (��,Mnyo�fg?َ�.:l�6&���
OPȫ	�����خ U�彴=� f��.�q[Z��V��}U���Z#7A�B�N1u�U^���B�i���PS!
Lꀈ����<
M�k.��e�IEM�0)�f<�"��ޓP ;�d���HM1���h�	��N��*�$�,��}b�6�y��������f�Z�W�24Oa̧�cu������(w�!j���ٓ�ٍ�LA�3����L'���X�T��{r=�R����SK��o`�=?�����[�<l!0S(D^�`��8�A����7n�&彁��������dq¦�m4��|g�#Szn�&gS� M:+�.�����r&�nh�H�� m�����Z�e���i�,����O�yO�%�0U�����e[dY���=|�2N�O�&iv�V1�������ɰM#ҽ2�o���D2�
F�ژ�0��(�P��מ�JS��zq�=�bN�e}<=�)vv�+o�:澽L�4�6(�Z����Ա&`���4��9>�ͼ�o{o��vJ���AV2����$����6�'�0�u�V��;	H��1��.����vpȈ=q��,W+��4P��8�ğv}զ�P��\�l/�Z^-_o^����x����n/EJ��`4� Xf=	�=��2�}<er,K���a>��� �d�����2�#}#ߝ�w4�F�ۊm����}Τ��Mz�6S�BY���d#��m�=�:�كK�δ��M�/���G���|�������wL����3�U�Z�3��/�:Bِ�t:>S�T�N����^�#+O���
di�֗���͘+m}k��`�wXDzG\FO��@
��#^�6�<Z0�{)�L{Ն�\J��{���x�w�1Wы���gӻM�`��6 !����w���:B,�^��A�!�K>�=��`��	`O�⬧e�&��������cK;u�3�O>�3y��J��LG�v曡�ۤ�d��;�33���8/��6h��Z_M^dَؗ���ni^�//�V�# 5���t������k�!�t��|�V�I7�7uP"��x���3���W�M���:�	v�fc����!/�����{�Ӷ'�݈�M�J0+��Sh��1o�w�M����O2�J|���b�H̝ЀR�xE\/|pL��>���[���V�Z��s{�fa����Y�	;�B�	�	�����d`�% 2/���3d����8���=f�N\�E�\����i����7�M�*���h�f�gWy��GK7CiZ�S��d��2,b�yN%Ecfc�ꗊp��2�u(����	l��K��dhY6�J4�*d�d���Mrf�b��ԋ�:����K>��m��)�Oj��Y�=��d'��^��|�L��@=O�mzp�<����Y�Uh �-� 偶�v�\�u�t�����}'{"G�l����iF�Rj�>��.l��|��}d��~>{q�ª�M53������sG��%	�@���>_��-��՗H �1���W	`i�*�+w*-:S�B\/w3Y����Z;�Gi8���B+�uO�p�Pl��]�^���K�)�¡"<�)=/Z9����
goc��U=��S(�ꝣF��Ӳ+j}a*��i��+���g-{�ϷrO�!�u���X̲��_�;:�{$_��M
=��ȳ��NP��de�������^�i�<B�-R'e_�w'Yʴ�����kSYL+ݕ�'�|�`99���l� :]l7���&޻��xf��mg�^����΃ ��l���=�G���&�+�d4��SH=�K���Q�~̶`�W�G~-��+��C���h]���$W4)�Iɯ@n��R�HX�M�y@�:�V�V�ؗ_~��k��k[����[�o=���Q�A��S��j�N{��N��������[��P����W{�r�G���u�����ӛo���WT8>���Ñv���@d��r��G�|�
�
�m���v<o�����H��@NzLG@��K�w��w�x� �ڼ�oi���<���R-��O��]8BG��[��eO@�r�60�ʳҟ��<:�v� aʓ�8����`�aa���	��&�=����ڥ��{���S�S��Z��J��]���g�ڠF��#�=��If��N��+�|�k�;;!��<�٭��8~�ՠm�A�t�נ�<F{E'٤���'=�mͦ~�|]�1e�uwh�0�f��3&�IK{�cY���?Oj���7ڮ�)��nS�+�6%��sŐV���4�yj[^ZG	����_��ӫ���yf���b������4������$���!NO����3rZV��~�������؎�}�7N�q�{�;MQ�ѵ�t���9�O�۞g<�C4����?��h����7�9Ro �k7q�Б� ��G:~�����i�� �Al����;;�<W|q�:N�.+�E�]c�&�6�ta��K<+���5O5k>��9}ʐ�h��=yO�ЀB�uo����cӠ �X�}Ch:"��P+��W�D���Sr�O��O�~��ỏ��َ���3��[/�V�3��Q��������l��-�*�=´/�9]�%y4�e��Y7�,�e�9��J���Szo�=�t�</p�l�ie���c҇G�vu��
L��@�+#N���1�:���b3yq������Q����N�|���������^����A�㎥���+�� O�~Qf�`��a~_�[�\�b��έgT6{�_Q�7��d�['�}+P�O�p��Q�5�q����n*�T3��x\�����'c���>?]O:���/�Mһ������6V��p���Mm�m����W�b�dW|j��X8�'�3��5^�h%'����.�uZ44�@�����������
�f���r��f7�R��܁"ã�����o��k��Oݰj��N�o��ܻw��g��G��f���hzx�C�#;��O}��կ~u۹H����:��6"�˜ �!~�a����hZo������G�B���K吣�i2��m�Gt�</L�z�Y�5����0���T�i$ǆ�I���HRyK��1���o~s�"�_�~���+�n���_"wh,G�.$��<��Ѩ�t}se)���S��)S�VH�������	�-�����=��me �nn��T���݇[X�֮��m��Ɉg>it��'��|>�%P��e���4��2���~�o�o�\����e��Rx=�����ƺ�7��ϷAV/�?՟�X��=�vĀ�,I3,ԡ��.-��_s;dHO�uK�yg^Y����&g-��oy+j�Ĵ��?���e���)�
�L:T�F�S����=|�)���������d�4s��1��;��9x|b���o��!-���v�p�2mַ��I��N���5c�2���C]�s<U�H���ٲ�E��|Vi�{M/���-��=��\�?)���N���:��8�e��K�&�i��8�#�X��1�g.��q�nC��i��	oS��])=��_+�8�i�&*ئhS��-{��Y�%�+�C@��oS�/u`���TL���br�>+��g�Q��ў�k�<�k
���~7 h>p0��ih�ʬk�ؒ�����&^��gY8���6�1�z^P㽣��`3ş'?Ҡ'ȝ�<��y>-�ɲO�����r�ё�9B�w湧C���{���O����Q9j ]:Y3i^l�~x���j3v�}ٻ)]9p�6�_���'g��u����;	fӹ4�7�x�@>߈�Q���L,C/��;�7�����{}��I�TW#�=b��
�I�#�#�I�t�xK�\	�:�W��ӯ|�WΧ�(]�,86�{�M� �-O\_{`:O��:�Gκ�w��UN�sN)]��/�=�n~�'��J�1��f|A��Z���ʼ�}dp����pQD�q�f��-y�϶z���|<8c��?�;�`Z�y�}�-l�V�f��9\^��p+s�)�MWf��d����MF�馕A�tr���x��wU�=u�9=�K ݪ��3|��rF^<�~�"��d�(���+7�kr�eI�K�˺�[�{���ִ(<A@�G ;_ąh�Ë����h�7��|�r���U^�/~�����@�P���A�r�����l�U<b0��!GS+aH M��	$�����j���_��Y(�a�������g�M�ԀHYǤ�s��*&W��a�s=�p��Q���Kڐ|r�Zq9>)q۴l���7E�uY�֩>|�)E��Ie��k��
�M�9���d��Ό���ɺ0�<�Ҟ���,c*2��L]�h2z����t?�m�?�%�p
H���~�2s �!#-�#�?˴��T��^��Y֣�.�پ��d��3.��y��D^��d�����7p��H3���*�V���و�i�Ֆ�;,��/|��ʺ�ti{��p�� ]���ZuQ��\��*˙e�ڧ�Ʒ�E�Ԧ�Vi��'��7�0O��J�l��� K��^��k�_��/���~�X��o�� ����Sr	|��S��zO��׿��p����{ᙷ��TTwE��>�=}��_���{�ox�ݖ簐�MBkS���2gZ�g��L��m��RYƌ'��A#9��Əؙo�� �eM�<�ȰN.��.i���M_$�Hx��{	�2��d���2?��mk�0��f�/�SY�.�g5C�{[�{)�9(j�jD�3�����L�h3ESZ�}�Y�\Зr;��%���ä�X��ֺ_J�yV�����s�o[P&�b/�Zyn� ۬���K}�kӉj�[k�fw�_,7�]���/��!>�;��X��q�Ͻl�m �����^l2?a��ًbp�@
H
�d�W�j2�+`�RL�m%c!2���Jų������@��_}��������+p���!� {�1�����i*�w�w7e���vb	zʃ۱��=e�v:B�+�*���/�?�l���e8=m�s�������14��M�ݖ.���n�\�|�:�iN�w�Vm6���M��ϴK� ���7cڳ[�V 7�~T�>b�X��JOi���>�����j���t�R�~D4��>�p���ɲ�p�{��	�9�͔Ǥ[]s����������;�m�G�3�\6P���as�,ckY��P�Ӿ�8v�-.���ON�^�g�-8�_�̞lN6C��
#�CJ3��qUZvL�.��t����Q�K��I��9}.��mT_�@�:&!m��m���^5�������z��Q�v4�/���	�G?�yE�/������F���E�sVr|�#�O��'N_�җ�r*�����O_����I�l�;��%�ډ<��YṮ8�����\�)��R��R~|��hR�[�{�b��E���_�>��%�vϳS��42y�eYӠ�`�y��,c�Wu�:p1T��I���i� ��I��'����������KO+˘Ϛ�lC�/l�8J.�O���2	g]��e��@�Ϸ{Sy��3։e���޾���^��<��l���?��O�0Ǯ��d\o�<'���{���#�m�e�U5��!�B�׉w�o�i��kS[\j���$�U��bHa���ޝ�2��F=���ՊPݓ�i.DM�H�~k[��˿�˛�P���u�ެ�G�z��XO��w*C�� ׷�ձ��8R�H>$�.�@{=����o`���J4AK����-xL�j d!�K�zqQ�g	����A��ck ����x6����}�s�8���
�O ��3e�i���Զ�@cE^����t�F4�;�<3���)`�/�ǅ7�C���%�q��ʴY�l�,o�� ��괹�K��6�;�.ef�݉���$�O^S.���=^[���^]���ORD����omS���e���?d���o�0y���!k�9�y=��x�6�=w�|��;}�����ַ6�������6e8R��J��,�A��f�y�����'Zv�,$w�`�9��d�Bt�[�&������`���p�F��
<�'=ji�E��z�G�}t]�YH �ˣo�Ȧr����p�=��s[���J�W�ij��\O���Uo��(�,��}*��Ͳ��IN�l��WS�dR؊���_�\�.�]���1�h���c�d�q\��޴�Aҽ~�D`�
�@�_(�,��l�M���|����Y&�?���n�4~7j�'�95�A����a}[�s_�=���-Ą}�z+gKD��~�vb�
f��40L�ɶk�7��~ήl�M�cZ�F��>v���Խ������m���w��p�Z㝏�M�h���59gf�8\�L�z�<gߟlM��ʓ<ad��)3OI�̧��9��o|�[(�׿�����l�[��|&Z=�t۞��%�h��(y��ͤ��ރ�p`{	e���j���!�t0�BԱ�`��@�F[޿N�R�I���ە��Ɏl����1�QPG���)-�{��l[VU���\y�˖L�D�@E�[�D;�W�	�y����@��mp�p�����(rG��A2se�Yz�o��J��Z�c����^�1����۵�Rk��61��w�� �4*�B�i� ��Vj��[����N�ݳ�o�C���yrb��@����Q�W��^%��n�Pn���S�D�˵3X}�:࿆�.R_s>9 _p6�() X�z1N��46�>��w�; A%�!�\�)o�k�w��KP��X�E�^��g��X�����ڝCH�w�[Vr\��]��Ȇ���7�2������&?�s�?gB�j߬�l�����^	S��{W����Vl�6�@{�PƦ )�����/]k~��B�h�h��q�]?��:�]|�Mų���9j3���|�ʙ�줰�z]�G�q�2��( "Ʊ��r<�Ifz�(]�*y��$7�U�C�Xdy���գl������s����J(p�����h,��q�ʸYM�J����|��I)7F฻~+.
�\���+��`�*���(R0K�h@��hB�]�M�]39,r�E&���N�l�B������r�� ׾|̈́�GʥB�~D� ��ޕGv��l�1�=�LZm(0��`��#+��=��)l�Q���+3@�A����U@�*R?��!z^�u��g��˿r��p�eT[�  �f���*��i������1��2�B��j�ýL?D��U��oW0����gH�y����F�E�������X�Y5��t�����Hu�R��JA��.	p����ή?|<d��:�����	~ϗ�cMd>s� ��d(�����gJ<]@�p��)�w�h�8HK9�s2e����}| ��S�G�bvu�����͕�[3�j3-�C���N��^�S��V�/��[p3/oٶ�Xv˳�-���/y�˪�ƍ��u�p.yy+Y�pV�=�u���'�ݚnv�J�G�x���]�Vy�{=�>��Z>��A*����"���ϗ��]���?x�я~t�&3�=Mu�b�&(a(�W�P~z�����J#"ċ[�j�3�c$y�P"���"��oU�W�� ���O"�}��r�%����� \��F�����>� es����D����%�'���vNJ`���i�]��A��~yڬ#�>mY�����û���m���U?�@�V@WR�s�(��υ-{4�տ�+��k��+�ȯ~�;��' ��6��u�꼜�l�]pA 4� ��>�)���ܧ�(c��� ���ʮ,�O���1Ċ�o*u��㲪﬍�w��A�"��N��S�D�B4 }�9��V����哻)�f�ݞ�~��i�2��Ǧǯw���T��Uȍ)+||��	�WX�p%���(,�����\���\�8�c���.�s�\) �
pW!�g���Z���pL I�nQ]���'�Y
k�s �5�sr&�B|Ix	Lk)�#��z�轺/���|�$Ɋ��G��X҄��<���k�5�D�a8�U��P-og9<f��;�G;hK}��T?��0J���l�R~���=k�� 6��Ǹ���Rj���l.Rv��v`R���֕��	~:���Vu�Հ�;A�W��SB��|pa�7��$�9�����[��"�γ|��6�=�j�����N9������2y;���u�b�\�`%���I�W����u�
&.�ܚ�g����\U�\�Ȳ{ۏ���w�}�ϕ�}�ҥ���r,�/(�j+�[�D��d�{��I�>~���[�i�jc��m�y��-rR�*�uζ�>j �C�U?v}�Q%ߪq��_'��o�xW���&�;n�f!oP����Z��{UC2 �,	��Zv�w���Ƞ��k+wM-_�G�w~�w�t�<&ˁ�(�7�Q&N<Sy�V�V��$8�W+�mhu]{��.��8��&}C(�L%�}Tu����/��F�e�Y�_��	�`�XD,��ɟeK�����#]Y�\�v`���)��(�S.R�z{'�uВ�v�O*%��>{օ;��)� v�"c{�E���R�	�@`��T��zwu����}%p*]���F�m��ɳ�w��]}OW7���&�7aݷ�~Q�ml<��ɪH,lwQ�(<��O�L��94��yO���b�yT����t�Bה%�� 0'H���z?Q��e���^����>_s�Ψ�GslD���w���<�Gt��@o��[�o
n�n5L؈�GZʬ\���B)#d���ܵU&�&��0dmu ��� U$��|Ld��'�c�4�*��Ê%fD�y��C�Q���0X��]an�9�J�;���:+�k����gchw_}�
�3���V;���rV]��?VAv\�?��ݻ+��p�f
M�ܥ���R=��o�>�������x����8�K��sYT���,
���N��$�d�-�WT�}>���	�(ΫS����#��<_Y�W���I�O�Y����r�D���nf,��*[���=zͿ�z��^f)��2~4ϙ�=�j�J�\�ҧ�ʹ�ha�$�[�;~�D^�]��>��?���ί��:���FJiV�ˏ��m7V/A]��`�z���m�y/e]�r�z܊f@��>�̨Ӫ��h
�;���wgV&��$�"r�&�\��%ơ0e�_�V��	M�S��+  �IDAT\�����()��$N�,�mR�J#����l7o��uͶp���Y��2��k4�:a�
t�e�70���sK�	�4̗em6�j AB0�?>�[�x7V]/ۥ�����uӵ_�|�<�e�qP��zG}Y��n|$�"���-t��,���8�Q�p�/�)�,Pw_y`����Y?w �{.纷ǌ�Ε�̣��^����|_�G�\'�eL�j
ֶ��y
��b#�~�V(<�;�U,�'P�`�2�
�h��怷U��lOx�+�l��������y���gw���9'�o��*��X�a��T�5/���[��2_��Z�_ͷO�2��kF{���_{� �	
W�p�Ԫ���-%0`���	��'mU�0C�]��Ѯ˿�˿ܖ�>��o W ��Ȑ�sF��,�r��\�1��i��$?,ۏ<$4Tv,)���|+JN5�|�%���U��7��G�� ��(N��>%/�9&���C��pki5��2ACݳ�ƙ���?RX��>F|i�+��f��<r��~�^�Y��������v`�� n=t����y��G��l�mdQ���N����+���彪�*�w�d�_i|B����-'H�2�@p�J)[��j�u����B����xާ�q���z�ͳ�\1Ie��T�W�o��c/m���ѵ��dGG<��<���z�h&��}�3�Y����̿�ߢ�p��qS]{S,�N���#r�X	�j��Zs�������o��ߙ��>x~�cS�|g�������[��[�UV�8�O��k��O�}����P��U_%�p�[܊I*��:�0W�-2�h�?��N9�h�|���d��"Dl�b�!-�p��@v�{��}�qc	�ќ���ߕ����>R����j[�{������q �� .D�`U��t�?����7���T���i�Χo#�R���J�'�ں��n��1��tޑV�|��O��;@�`�d|��)6-.D l��x;��:�_�-�E��<h��~���y=]�r,g���X��\���/-��������1]p�/��~�q=G����*�@\%/D��nPW���W|Օ/U�
���G�r�R������Y�r UR���K>� �+Z��� �$��x������"�r�@�]>������J`�ov��ϙ��R(��V�G���#�>�*;a�L�*��=f��|��R6��zh�PX<_�ɍ��n/S�z�Z��U�G��^��M0S���ʘ�R�l���T���z?  0������,dD��>���g%����^���q���Ғ��n�r��R��4�+|-�=�\=r���5�B��#e����ļ̶H����'�u���u�ڢ{�j��Í�Wϥ�Y��x�U����w���ΐ�s5:���U����	~+>�Rު��fg�Y,���3�{3����l?�%rK���P59:������14��/l�tj�c �{����E���r�EF+��cw�{�'z���gq4.+E �&�?����*n�nD@n'a�?�`�MZ��P�����Y����ꝕR�-�3N�.����V�Ya�)d����l��B���x/��w.?���jϸ�bi���Ϟo�+��k�\T�rd#�X	m�	n=���zp|x9]�۳�9������
�5���������"���Jg�&ݦ��}���2v ���# �c�j�*-ï�>H��e�����m��K��=D}\y��r���	r�{%]R�7�P�JN仫�T�����: WUl��P[�����t��[>��Q%�-��<�A.;u�ݣ�t�H�,��XCsy�'��`�����z���<68�D^ԋ���F~)pW�R���{GDy�O<~Z�x�T2O���� \�:���}ZBH%��v=�}���Ni����+S��w�*%lG�4�U׹��yY���	��H˹+�����ڏ����M�xt��*�G�A�YX���Ю�U��*���(tsz6潞՘u�E4�����7�72KϢ��:�����8��}��j$��еa���P�t!��͏�^~`3]�gG�b��=��KF���j���H���z�T��i$[�<��
�b�Q[� w�f�������;:^�����h�+p˹ﺯ%(E2Љ#:(?)bZv w�f�9� ����/�v��X�z�N+�M'M5A�����*�,�����}�}"8��	�m`Zc�\�W�kW� 6h�����	� O܁<L��n~��;�`t}Đ����1�pI_m2Y�]�jsS�'�C�)O�8%x;~֮�dZ>}L����u���*;�sTc���7Ҭ �����q�n��jn'p���?A��v�8����G飾#z�G��Wӗ(;D���������� \�^����Z���v�u��i���EW��2�1�f3��u�Mp{N>�~�Vy��M�Rɟsq�M��N�̙�i��޻B�|N 7�B{�{�r@�3`S�t�-�o�^�����ͫ��t W�V �k_��&����i˅�%�@�~U��^�`�",�*/7�w���&���k��\��q���6����n@�a��2~5�f�`���1�
�`�x���X1�u��{8���rP�Og5��>��Np��mGy�m��]�,���7;a���SXVLؕ�jv��Ϩ�����2��v��o_ea�r��J�xyV)�`��P3�KY�LWSw�� �TlE��j�6w寀���l?����V�'M��ލ�E��)d��v�O�p���H	��a�_K��H�zm;[w�jR�V�y��u_Q�*�x(������f�C�?�oQ�mF�sS�'�0��a�����U��P%�RHw�l6�;����H01Ymu ¯���o������������\�e����peI�����I�v�T���I9�rW���u������ގi�up@;T��r�w��c��j��3>�X��� X�f[T��`�a���=����y�F��o�ڦBV������|wZ�� dຢ5��[�C��L�t�O��r3yu֒�*�P�S����aķ���o���t�� ��K���S�^�s�U��_y`i��M6��#����D@A�E^���-2D��ߵ����\"m�d��ɨ���{�e*y���y��~�ь����mt.N�#����,�M��j�oU�j,T
��͹����1{�����'���������pc�L�d��F�̫���h��3#�*�qb)���	_���7��`>,��))�>�@ ˣ����~��<�Z�{T�$���&K�"b��@�qv��b�֨���Ȓ[C�_���ႆ%{��NKW&��Z�{�?��>)l���e�S��c{)e�˘����9.'J��n����17e�aG���~c%���	)����~�`�����ԁش󞮜٧~�R`�z��.�(-~�!+,zN
����j>��D(Aʇ�I�I�U�pʲ��0���f�����Jxy$�Na��ܔ�'��
xUc+ǞσM)����:�a�Kt�%���)��!��9� ��A��>�s����--W�4z=�:Ϯ�B��uW;p��ᵒ����vXs���[�f
�^�0@�9ԁ��3��ݹf�����~B[��@ߴ�KG�\�V�������f,���V4�"��1�;�o�V�uO�E�芁����j9��K�,U�H 
��#����>v��}hc���w!�%���"�Hu&��)}$��UJ���Nh#0��?��%l|����z5^�l㑖\={��re�w��c�;��p]@�VE��>z^cN�J�f�r�Uh����ï%Us3�n���t�U��);��`.��g�LF����	�\�<���Q���P����xW_qĶ�[�@( �/����9�N�wFB�S*�=k�����m�>�(�#p�uI�Q����s����Ob�bh���F��l`F��ĸ�k�r�Eg�vu�k���1QY�;J�#��y����	�o����#*~wI�V���ũW�X-[W�J�ZQ�������ڑ�U��i����M+�"��p��f�R�[jNL��'�MA��
dʝ�ct5Y��\{]���L��t_=#.z�,̿�˿|���W������CLӣx;�R7a��z��]��K�����:&X�ξ���m�^L?}�}W2 w��ϗ�3�����I�x��0�|/���It�~���O �j7&�wf�=��_~��ӯ�%���]1�U!Wչ�
<S���E;98���{��*\]���]?~=t��P���>��X]��w������%S��>����j�ww@���ڬ�y�{���ҁUW^��@Z���|��1���U�zxI ��U�����w�s��#��5����K��׼w��9@���ќྦྷ��&�H�����[nl�$�{3�@��M���&�M�������o�s#yu'v/���0t��(�&�}�0}�y��)ˬ�p%p��83ú��MieA�j(�җ�t
��%��Ъ=+p��T�*�{���MX
��r�k��k��Xoq5pk��[�8�,7t̬#+�����K�X6�E�%xuЃ���b�~�댷��7D�� M��戴"�,��C�yd����5���Jp�,�X�=2�Z����w@��4�S�{����F �A��۴"�*���@��WJՖ�*#���~p��"E��_��j�?�WlH"_�I���b��:%n�g���aU������'ٶ9�����?�����tc�2���9�+
F܊�_�k��	�Q}8��c�¿QT�QPj�Po�=�E�c��T8+e��۩��v�'�T�4�m ����6�+z |�DQؓ���^�}߄ ��E���z�v"�>�����p�P0bT��K�t:�VVT	0-� .|R#�G�]�9/��Q�����7�)_amvӷ ��#�?��������KQ2B�>jgN���lY�s�Eo?��v�\i��,��A)�SX�}�)-���bE��<�S��R�	��PB�]Z���)�����+��kX;���Y�#�]	���Lx$�+`Kٳޯ�e|t�T)��y'�.�,/���/�+��	�U��?��qոQPFF�*M�_�ӽ��� �Zm���;g`���V]��CX E(��{�qҤ�%�Ss�=��-���
��q�y�u���dg�Q)ٶ��9�>��N���8V��7Lܔ:��
�Ao=��#��op��U�>�Å��"�M)�k?���BbTLZ�j���D�F��X1+	)��y��B/Iװ���{Y�?��o~�q�,U��"� �c0��I���lX�4�ur!�:�l���"�.�����V\�a�V`� �gĕ��Q%@I�w�� O�G�
�
�?��s[I(�dɲ5@H��q,F(e[W��{�5/eU��@O�H^���;���΢�i����C������Y�V�y{}���1�G�7����9ǘ�
�E|B����⒤<t���c��nW+4���#�z��_��JF�|��TR���;^��0���Wr@}�k�%������/�+/��u����<�n���ь\��>���qY����/r_ϥ(y�A�K>fcj/U��RJW��z>����~�������tZz���������=�K�LN6oiØ����XX"�*��,��{X~�o?���7��@�'%V�ϭ>�~׻�~�W~e�շ,�5�B  2
.�y}�$���o_������Wu��/����vm����Z\�]m`������U
eg�3k���d�l%�����x����O2.)X6n�OD� Ra�n%�M���� �w����#˙�Nזdr�9��z���U �:d_{��q=���4��f\�Gn	jw�J�ƺ����5/����Z�#������s��*�J�����jN��j�U������^����^�]|Dʭ��X]�rAxHYpe���<��@}����;��C���[<�^x����q�.�|��A�_h$��u��R�җ ���"�nT7�T�+t�[�\Nt�W������g�����'�	z*a��h�;U 8��@M��,@�ʴ�K�!<$F�k06��� �ϼ�g����{O�M���Ii��Wn��~�����4|���f��Epb�������|�+x�����w\�}�w�duV����e씥���-2���W�r��8��FY{d��G W�N���J}4�OK("�;�[�X�(�*%AㄱLx)"����_��fD0�|��>��l�%��|*�Z�J����*0T���l����O�l����J�U�U_X��[�l��O=yR�������m�`4���M����>��Ӹ��Yn��ݽ��;�����z������R���¢guM��?��:���e���2�����Y�F�H{8ج����T�m�����wp�u wW�F4�InP�qS)Y��^��N�x��)�K�f���{T�]r��bE�ZH[1��V�T�|�'�З���nb.l8� 	)ߨ���(T���h����1:iᚼ�ߏ��vپ_�Mq		$� �,@Xn�zYJ&D�T&��h�T���p�/~��r�/�'(�4!��T�'Le�6��%�'�u�(��9��@�̒�� ��cmɠ�j�ȧ?jwYᗧ|t_ W�u��E4>4N%���ַ��=��X
w������G�R:�� \��0!<��=Z��%���%�%�����n ���_)�X���G�d����)�\x��+���f�xMaTWҧ�O�.����=>�+!�F�P�
VI���2��{5��W#���>J��޷$���R<��7J�*|r���s 3q�56���
Lf_�e�2T%��B��FW��3��*߮?��q��+�u=�!��D�3���
;���MS5g~Z(����w�/y���y���,��C&LB>��)P��T��U��Y �����z	�a	(d v�����Uz�%��_��p}�ŭ�r}'��!a���ש����9 Y߲��%�����>��\��?��i�.B�}�; x�UEe�Ji�S{�H����+p+a�mȁՑɾ�u��+
W��C
��,aG~�.�H|`��D	Q�%$ �j�q�/�w=���e��ae���%���uaY-O����ܿ��b��yׇ��������R.K�K}�!����T���c�Si�&���M��o��t]���c�Sf|�S&�6O�an�O��o�y�*@q ]mZ��#�LW~���~�[���˒z�R�ݗ�x�ƃ��X�c��a36�:>]�
�W׺~�q@Z�~o�y���g%p�G=ER=��&2��c8[�39�)`޿�_�j��4��ݴ�3�[��f�{D \��]��Nc�)j'?���MMZ	-�kc�U�ӷ=��p��ǏO.�i���@������ݷ�АP�<��a��_�{ܪA�4g���_��W7�[Yne��o��rS�ĩ��sӆ7-�{<��c�/�<: ���"Na{��{���5�8#�����
k�,6>ژ�eF�� =@�_�Rm��	�G]EnK�� ��eO]VA�/��G�37	�6U���T��Z�{�{r��Z��X\�CY�e���傢����o�5PsWiqEѼ��A�Gi���Ǜ����C�L���l�#�����㟊��T�*w���H���7�0R n�J��5�n9A�m�7.yoW߹�����������G�vy���iD ��Ζ���cHJ�ƴo0�x~�ue��si�7�4Q5����읹�y�N��ԸG/1��s�W�F��9��8U��5�p�NVMVś!����ᛚ)֝n� �3L�}� 4\�Q:��#MY>���
�^��V`�R�)��S�$�e� <;��r�a��i�e�����k�v�MUޕq^���!��\3OR4�O�I�7���Kʉ��S��ڏ%�P�/c2wu��� ����1�F`�������2�*�H/��"�k
�J���j}M~l d�jh�룾� ���]V���X �-���B��]�X�	��k���#��r��} ���k&݇V���\���+�'( �C�*��poPG7��:���!�������~ZG�])-U�z����p���5<��ڀMx�O��3�����@�_����mSʜJ�)}�=�����I�|*m?}' ���+�'�}�`G;H�K@l;-�ջ'����y����E�<р=����A��/�����&:,K�{)��Pࠞ��a�Ģ���`?F�Ɗ� �}��͊P���6��ڀ�A8�Y��U95�d�������:G�( 0�:���I��φڸ�xYG��&��U�҅k% 3��*F�髼=M�<�d_�~��ʒ��el��vtM�W.M�ߊ��ռ�%P�X` ���\����y�� m�ɋ���T�FώSx�Np[)��~)?x��'����W�tO�R�76 �����IķF.�����Ԃ�����Ն��aū��\~�j��Gm��o��?�����y��q��K	Ї#�+7�s��e��Ӫ~=<J�^�5Qe��4�������t'/��\�(��2�d��@�ʓ3�<}���A��$�8Y������(� \�Np�m���x�'��q�W9���/`��W�����b9�e�2�U-(�%��G#�R~�,�����뛎�a��
J�D��_�g��>��i`Ӣ�`$�t�V^����(W1Yi;�~�'70�6�8�O�q��+�����!n3-�c2	h��lx�h��d��{�/�r$����Y�"ܟD�R��P���@�>Ӹ��r��3����?�'��Ə���:�(7�vmY��yA��ȭ_w�owͩ�Ŏ|<��8��ښ�%pJ���7�7��O0��vE=��3� �9��MD����\�6�~�<�x�=W0s��0F�E'��.�qa��ZɌpzc��H+|co~Ј�T�f
x��w�;<ɬ*�*r��[�OԊ�u��i��8����DV3өe��=#/�3�Q�tu��#r��`Ǘ�Y"��Fl&cC��,��U@nB�,�s@�� H���-�"���B�����񷍡W�xR���wT�oUì�"�r���DJ��k��6�`��RD�(Yt��w{�ICm��Ĳ�X��zW�܇��d�;o3����m9z��o���])��s����U�bTFQ�21� $E��T.)'�C-E(06��"����/m>�(i�O�P(||��R�M���g�z5�V�ɶ���p����)�YO �H�0�'�W���98��hٟ��3cZ�檝f ��_����s�1a���y7V�g����l�@v��Y�Y�ꚏ�N���~g��;�hR� BE�#��UU�{,�`��pb�\ �]���0`D �Mj.�H��ݕ�%��Z:�^i$�?,��_��_m~�򿕅H Ru��e�Qy�e9�*C;�B��q:K���~�MU�c����?��镯]������-3��,Ԫ��,�G���'j·I(JGe�=��%�:Cj�� l����l~��:���7�um�i�i͡o�/ԗ6=]e���/���qz]�N���+4,[cm��]? �|�D�a)O�C������b����7R*F�u��;ٍ���4�,��?G�V>ÀK�aa%�+�CJ+
<J��0�,�9&�*_\ �̯tE�xoU�L�)��w�E>=�e���x�+��{����o��z��*����6z��m��Ra����ַw��ө|V��U����Ϭ"#F�`��ic�=p��dȕ���.
�D<C_Rr��כwV�>;�ǲ�o��6U�ج%0K�Yqz���������sl�9B��<K�n��雍T�G����|�pSp���W�&�l��~U}F��
~z���A��=G�[�Q���C}c���HJ���|y�D�y q�pF���*���^9�*����׽o��w��8I���f�,���՝�<>��'���I�(u�[� ��W��{0�����k��i��n�sY����8�#��B9r�x^+��+g�% W�J��j{�3�1(2����*-��Mc(�4�D����0�-��9�[iG�}�ѵK'�}�{�0eEV�Q�7�u)�qV�|���=����w�ҿ�4���3%xϻ;)7����jN��e��Zm��t��@��ii^��� �����H�P�?������ww�����J�Ң�����T�aX��CQ1Y��L��w�m,C� �(?6-���1�*]N�*=KYj ����2&=��yD
�U�SOb�z����� e��؛�硲�r������nb���4���K�T�r:��X�J#`LU�{X��u"�#���yT��#0�
��wԞU>�.�ں �:�T�@���j��1���^���LW�A������`݅琇�KY����q� `��������M_K��z�G+�$�2��ڶK��7�<�2���*�x3��a"<6:�Q��>�� ;<��	�ď���ܽD|��V�Y�]����\iS�d)�Ki��NĘ\M��X��ey�{�F�*��g�~��gi/�+��)3P�a�7 �j��O�[�%Y	Ǵ�hu�U#�+x�[�\�!IX��-t]9�ML^w��a�RL����>���n�V�[�>,��&U�W(�wߔ�̩7���y6P�"`8���<��]+/W*<#A:jV��%�'��s<2'ީ_9w^� �#ᅔ��w r%9�"�&�p�G>���6]QF�|�����io�t|����ب^�.�����
��[cB��Æ}�� m~��\���/��� >���B���o���t����}��Z�	��|>�[������Y�@H1�TpO�<v77��!\�M���������;�[��̀���O��y1�h�0'>�q�8��q/e�J?U��Z����� nE���f<���<��%+��B'�NS��dt�t��R-��`�g܊��Mx3�4�J ��K���r���}h[�ڀ�SOoB�Ȫw�{�`�*�m��"��%H��}���ݢ%� 1��gP&���vF=�Zj�>��8�[EE�EQֹ'�oo�e�¨=)��1O�ʋ��o�����-aG�!���M�ld�£�t wD�9^�_*e�\���GO_����c\���M_Y��e��y/�����
��8W_T�����O����\aA�u��� �ऺj���?{i�V�
t3WN�2���Q�6,>����~O�P�kT����zV2kf�����Qw6�[��^u�g_W�k?�Ǖ������y�b��j� �i�+��Q�i��|K�mu|��u
�
��`>lZm�Q�K��*Gg4Y�e���΀�S
��(�n�nO�B�';�җ�9�F V��+_��ƸҴ�K�q]��S�ŵ�Ryy�Ni��N&�[��dv o/U
E:��y��IY ���pe�dsi*0�;�ٰÆ&g�sg/�R�YDV'��J� k3����\9�A,�q�����c1�G�/�Gᤴ�I�4��t�9���꾷[v:�<`+��>K �e��̿+O��Z�O8��ԇl(�96�^.��)P�� �H�|y�p��:�o6�9P�"�d�u
E�&{i�G�#<���l%������Go���9�b��J�+���_��x]���&F,�3FL�ց	rI��^�c#4{:�թ�#�[��;A{p�
����?x��A+���d��h�V%�|���u2���LF��k�&���'�����|&5p�{�Qd���Ձ�a!��6vi��%@@S�[B]I����w�|�@05d���|me����}�� �Ӗ�V���IE��n ����u�˸�ӵ{�0��s����� �F�� ��I`S	J�Ʈj|�d��%�>��Y���\x  ��`��_<Y�X��JX��hx?$�b��V�u`�*�w
��h��W�;˖SYJvK,ᾰ�;":
�����8�/~�Q�w?&�1 �!m����f 7���8�����xϨ��}����e����'BIEQQ���������;|�9��}w�ЇR��>\��#�1����
T���]���q-医d�Ï*v��m>s�Z�g��S �g�����*�o&��O��j_U��"+V���f
��F�
�V�g��[M��1>`=���46���抙Ъ���i���v�<�q� ���Q��W�dU������:�=ޗc K>�\�������Ge)Ϻ̬II0�rr.",1 �ѭ:,y�>�FH{��ĕ�s K������+(Ut�J8̄R`���X��f�)���P����i�'/���Ѐ��X�N��h��=���w?�v��� ��U��z' ��c������F��̫�K��F��Mc�������o���ON��D(9z�:�v���x�JQ��j��c��)��ܪ~{�>�G~�'<ۏ9�޽J]�nB�|8'��*��L���i�07RTF��Q��fW/�*R=�1=.�ܹp��8��a73K1X!�q`��7�?~��&-O��X�~(��{G3 ����h��u��}ܔ[�j?��˻�������R[	�T:�Ř�0SԨ'`V�@����)]��= ��3��h�>}�̧��c���	��(y��ǪR�gnf�оb��	�Θ���@��M���y��.�^�x�2~|�))>���֧�A�cO\��c�1�_�����*��ST�������OU^����r�{�[�Lp�帚`�u@�+�oj杬�x<��U���G�32����I��y�ۚ��j��ے��]��V)2�Pf��u���bW�l��zګX��7��?��2D݄i�U�Y�V'�
u���i���/��f��	�	0{�n"��rƗ zde1=�{��6Oƿ*8H��A.��������*��Ax��\6d <4�������^=�	��t���S�k|Ҳ�(�ҏRE@�b[ދɩGv	�g5� Bc"����6���)CU��*��i>S�]5����/��'���:ϧ2R��R�GuN�ȭ�w{����w�{;uN�&�LRz�Gߦ%���,�؃��R��w��*�i�.�^~��u6~��w*��H &"�=B3�1���&]Z��(<l��l�\`e'Ǡ�����
��1�X����Gw�����n:>�UF��ȇ_4��֕o��*e)B3���>��M1˛E]���+�X���R5��/�NrY?�'1�LW�J�da����U�/E3r�̹!��>Ľ��؆�FuBؤ���P�G �:��۬g�v��V���c��|���r��Zc ]"Wx���L���s��
W����R6R漍������VE�z�G�\�/�ѕ\0<ȿp$�|}�V>�Y'�V���|�JW�N`T��7���&�IK��y8�	��:N��\���� ��Z�	}��R~3�=��wG!T��͉ �����6���^�T����ږ���<�է,w��
�:��SO'�J�c�d9���Y|��DB�4��Ӳ�|~�j��~���U����ǀ��J�UM��qO���۵�o>�1<��i��V�_QЪ���
ԽU����Q;x�+�YU�\��:��VK��T'����+��R�5 ����Xn}��J9��8�<��>�n��r�+�t�<,Lԁ��W��}}���w�e�S��@��	v ����b�ˣ,�jO]�%��O��E��La��+A�l��0���~;���G�$=]�]�/���E�X3U�W�e^�z6�Xu�?��2 �%���DY4�ף(��Wu�1�c#7~r-�RbG>��{o"LG���N��3�#������^?���G��y�B��?��+��2��\��; _��EC�����y�6�(�[�Ǘ�A�=g�uJ��}�1�f�M�c�N�?�^���-+��'��e�"ܻ����uĀ�L3�娴�,���cE���	,����/cv�넕��S�s����*�边rP��-�] $�{���+�Rx�W�P5VΘ  7@;ϋܯ�vH�{j���!��`�c�fy��LRu�*�g�������O�ܼ�@>Ǟ��U>T��u<�,����J,��%˶U;P .��	�e�MiT���6�
I>�Җ�\�q0�i{�Ì�u�|�}mNzd��y�Q�(����lH$z>�߻�ߵ�M�+m�ʤ+r�c�~��vÎ>N�	"��h~yg�Wi���MCA7�~Z��9σR�.�8��k��2aE�`��V���$φ������˗�фd���	�[0�1�w�Qg8{��2�=�}��r��6,���C%� ���l�"�=��W���������s��3zϧ�Xqp���������~n����A� lEn��͑��|�s>�)7FWyG��ݬep�0A����3�ޕ�㇌�x��l�һ_"V[�<_
���%���+9�||�k��u���=�30[)�#�������D�x�	y�k�Μ�7�oX$�l�&Qd�~2W+}D�Dt��#.�ތ�������.��#㨎:�SG��NY�F2Ra.�����[Gk�O��J��wu�ԃ���\������n�����jmI�n�����jy�o�Xf�]�������Q�a>�V ʩ6RH+19�Yӆ�OEn�c�b-A���:��\
���޴)\px_��$r�g;B�0�]��q�E�{�~��i��2�`eN:�f�W�`5��G��說b�fJnRU���>W8N�{�����e�	U�N |��ɇ(#>>x�G_�<>�F�p�'A挪~�:>���R�����h���=�X�vd���ǚ��=�1�r��׸�?��sdtwY���r�6m�=ぱ���jYo?��n��x��s��ts+�=�Z��sy*p��|O�P�U��� �W�:9�4k�n�d�Xp�R0{a
�J�t�rD)�sC�
u��=e������Tui+���|o2Agￍɘ�3�r��1�����Yzu�u��w5�ϖ�pDR(t�sWh6f)�orW?��V[�5�|��|d�����	`�%�\�N0�1������@��	���������6*�0�����i+a�.D��V�����~�_�X<<��+�GۊP�R����n�W���Vi�'\������e��{���gd�
CxC��G<�+ZY�������P�>��||瘾	_�����ч@�?F��}���T��\�P�9��J�~/�Лp+�=J;������S��}�(/�ʲu�Y:�l�8��v��</�Y�ՆrZ}�*�t�0^�������y�ua����L޻Ԅ�'��i�J'��M��-Ei9q��F�Lv������o�F�!������ңz�W�z�W�Q��Y1�,G�������F�䛙��d+`��Y;x�҅���e���v���;̳j'��FL0A����>�(K��SQ��2��j4�\Qqk��I
�
�vu=<T�80��.yyD��]1H�/u<v��+l���!��!!y��,�����-��@	pD�����m��,S�~'B��݆�ť�͖�7!�p�逊�{��\Z��˳�Y��W��2��w�WoR�,ˬ�� n����d�oʒ������錷�.�i��]�Δ��FZ�39�?Z��W�ocBV�g�;�R�\6���˲�hH����H#�oT��񌥍c8ݲ)k����u�W������3;��:����,�71wo�ǣq,r��|�-�d2=��=�����+r�&�כ��ܦ��E,ͺx���X��L��&S���J��"�n�_#w�=���+ۆ~�~�1�}�������V⮎��U}���n,��3WH��V�8���n��ʏ����<=�'�N�p���u�?*�F�]�ٯ��\Rn����ځ�������x����]��ڑ1�
nU�YYgm��3r\Ϩ�ݙ�J>7M7�MY�Y�ex���7��-��e�@h	�V�`��r��P}
��Q�.`�aT���rNʮ~����\V��Q{d�u����uaiNB&'�� �' ��4�����0٤�g|��<X
s��e]�����7�Oe�k����j >��xy���v����9��z��'_��ʰ�v��*�$rp����|�x;��E��oUX칗��(��x����8�t,"`П�C�vذ��[�ϭ
Y�VyT`3on���߈ߍ�d�;��x�o`��ۺ�9�;��EQ坬X0Q��'|=t��!�p�����#W壏(�~���y�{6�[\�<�#�_�����ue7˖��{�_�������|:�_-��}+��\�g���+yT�%^�	9��a�*�9ꈪ*��1��Э�se�Q&f�c���+��Z�̳��i>��U[^�W���Z�|�<䗃,����v�{�?�<ܒ>�nU}��&VS�Wy�L����B5-�	 C|�H�J�%��jGU��[�q�TH�_��v��X��n��e~r���7e&��c/SMa�<��Kn}f	�����,-�����e��"]��}/#�=݇�vJr�xƅ[�91���.Z���嘞���#�+�\pE�'a����{T�C� Y6)��-QD���#�`��'e��!������}�1��R��ާ�UΛ֧��ԥ=؍�\ٔ�'&��Ɉ���Օ/�_�ȕze�:%uu��,�#mw�"�Ҙ.I^��oo'T�T���<k��w�EX̔�*ϕ���� ����(p�����;�� 6K�O�ǑؑN�~о��¿�kW�N�I OYneq&蹾u��_<��ukʊ�P�ͥ���$`CZW��Vuv0���yҸ53�p3��e��>X�3���u_��^a7�>��ƺ����=,��X�+U��w���.�͕ǎ�Ϗ���n�v��-v/!�p��T>��=j���ӳ�^�O��sz*OXo���h����~��+A�-m���}�ٸ�`���W�y�hx��&VY}�p�ʂ�[�P�j����s���a�T�`/8�gn�.A{��H�TiS1�@u'��i�,繴�E�{q�\�gR�Nr&�˝�C�cԝ�8�	`��޹�P����\���3�@�M�%&d�3�ʕ���G���]�<�Y�g�����K�������J��D]i�Ȯ$! ��jȋ��r�r}��ܖ> ���� ����ύ����������

rk�-ަ^�U �t<r���>.���1_�t���Y��6qE�[�1���[�+��(c�稏k_a ̻����< �x]�;��6�xN�*^#J��
�u�%��l�"N*!�\re(�P���6������	覯�Q�z�c�,`�0��t�AI�8b|ms��7�D��_�m#�V�����G���SO�,��W�2�@�N(8���3eqU�W��նY�?�4j��fߌ����]�͕qp6��
�g�]�}�����Ŝ<������W�]f9v�}��&U���_=Ȣ�0p��-Z"1G	�g�~}I^��~�VK�+�(��\p��jXNU^��#F�Dl�˲%� �"�D~hˢ�eLm�K�/	w����)������~�bB�q_SڔMs� �|ΝKS�>�H���*����*�>�����s�^���h�o�=��R䡧<����(��P��9�Ͼ�~b�i��WSJ�[)�,�F�?/�:���:�Ϭ,����������2羴����"�2��}]����\X�>6�|�ɫ�y�Ϝ6��O:uq� E`$c�o���j�����UAn�3�SBV�������|���J��������}� p��L���ʵ��l�s��A����D���Q���(��O��e�;(��]�܀����4C�e9D>W�b΁Na��D:�eg_�F`	�"0!��e�0��WZ�tP��(C�y���4"�*����L�S2 ��dy\a߼�\!�q�4G���+��I"{�ܝ�� ���2�u�7�+|[??���O^�ɩ�r	��[�����\3.s�ߣ�Ud�{�綏�K��QԖ(8~"$���=��ӏ�@�S�16wm �ɧ6`'��.D$}���f������>�ߕxw��5U}�qP=�5�������l��Q��=�����F
X��e�wm��w５i����	8sL����z�Ǩη��z���L�k�=*X�v�HU��2���;��/����{� +f��Jˬڲ*k�6V��g�.Y��w��*UyЮ��o}�|��{���2�R�J�N]���2�@��D]O�u��:�<��u N_N�Z"@��!h��o��X�X"�g�2슩0g\��:z��F�L���JC<M���}ӊ�#�k�����j| ��n6�Qf�%@�uv�� 1���	@0v��sg���%����U��W�YW�q�p�c\��^u/���O��,��x���ҍ���??XE��@.�I���u�o潃�T�p?q�\�ix�u�mW�w�}�^*�t���+J��<9�WU�
��67veյ��#���,�j�ռ�1�㭻?�{t��;����z�ǌwU��u:ɬ��}'�X����^��O��g����ʍ0}>�r�ۅ�@%`u���گ��F90���Y�Չ<�ގ��Zҿ�˅ �����{��N4]�����F0VV�L0d?�f*��C� o[��'�<	(��?!+�6ǁ�G�N� ��6Ⱦ��L���_Ok.�s @T-o
 �])`�辠n����۷]����o������7�:�C�å���YWZ�}:��3��u��V�G9UV���5�r+p�����W?�s?����j4'v�[<A]�N��Ϝ.F�I73���e�)��Yj_VE8���:���Ly|x�טq��c��Eq�p��
�tszD����������>��mF\�D�h ��k<h����z_d�]:���T�z�M*�����9�Vd�S����գ��ݫrU��kUٲ�9]��x���׻�D�u����j@u��*��y�{@m��Zea�o�u`+�>�h��mZ��?�H�p��Bv��3}%��>~_�Nc]��|���>��sĢ%���˿l!	߬�m�Ҟ�����u�r���(�y�����T����������o.�����F����FBwY�~�q~��T�A�2H_� �X�q�-���++�$�i��V�c���E�� �澻D�]X�|��U[��s��n���>^QL�����R�o�ʊ�<�G�������V���;�}���/ʖ+��LDL���e�������jG�,�r�e�ћ��	ʥr�]LJ�>�;�9�$��M�i�;����~�t�(��Z֭�co�U
䪜�Q�O�F��j�Jvs�k���@num����;�0*���*�%��Z�wrG4�Y�|��3洶&�JM��f}*!���-�����ʲ��������=	��P��!aeؘ��J��R�$���mo�v�*�@Ri8H�b�Ri&�)G7~Gu��� |�MK`2,ʡ<�u��M��v��{�\a�e6��eJ�bM��X�G>�W�)����pSʱ��e>���۞yݟ��;* ,�*(R_�����%�>�ϥ���(��
�SN�o����{��ޭ���pF�HR�&e�շ�ӏ�β�~��/D� ډ�]/g�vY���4y���>#5�;��W�Vy�\cXu�%�����䋗���U�g r��f�Q�<���zt2p/��9��Z�a#����*�r�^�����)�k�(�2�I~�8��Y�
�q&��@�d�|3T�����Z5����7�j;��Z�Y�t��I?�Xl�$�~�[�/��r�h�{������R	SYq�8L_*%������D�ƘoP�z��ƭ�l�R�����;7g��)�.я�_��=�G�`IW��/���f����OiO6o�Ĩ�d��7�Ҕ.7�UL��r_�h?���3o{�d����|�9
57�y�X���
mpS�򪀤[�*� �\����%+�������$E�q���g��18�˹Ę�_>�\iu0�n:AB����%��w�m���;�{�l�I\�
Q��������Q�3`t.p���
�᝜s��C�sU۟3��V���g������J�0a��S��g�~U���KM�k��#i*W~�.5Q��v�>!yn�n.�f�`8�e�s�G�`�"?j4�ȭD�����e !!)���?��NG�V>�|w���I��F�Jef��+��H�Q$ ��_�|��>�:�u\�U%�`X.Uo|������{�������H;郋�\<��-+/ut�+3m0�������c�V{����Ǌ�K��>F�a?"�2�f�K�e��OUcȿl���V�,�2��Tc�%F��Ɔ��c��] ��(�{xਭ<r��?Uύ # G^j�D]�����♮{����{���#�0��^)��Y}wRG�c�&����3��i������un�|󞗫����ޑc�*c�W��*� �b,��s��嗚�*��A�OFg
Y�\#�tWp�:��WL!�QQ7��~�ӊ2��,�*����!&(�����%�NJ�+�!1D=��˚ k�I �)���ґm��7R��Xpe�§��h \�3�ͭ�r|�2}��2�Ɓ����m�yC�;�+�#˞��Ͼ�gX�V�d�R[���|͎{=��tV����j��Z���[���f1��c����	X�< W� cJ�+�Y��:��7���ɉez�J�\O��zK)���s���
K)d�w�Z]].M�ܬ�e'3V�� �2�cYi�y��'%���Ag�ߪ:����rZ�K�����)��G��i�f$�*w���wm������.�^��N٬ޱgL�{	~3]'[V���z�f���n�y9��
5x#�:s�}��7D2�Q�Ug8��6��X���by>ՠ��U�ѳ����M*Y3��(K�@(�&�	�դ�h�>�D�p�p���,���XYmi�N��C^����_Ľ�W�w��#��|�?달�(]>sS�|K�ٌ���pv���0�}-��F:��|�W˓���.��휋n��)S'����z��V��:�1��ݥ����)3~;�מeU��L
�,��Cw��-�eS�H�Ѹ��%�h� �DQ���_��x�D�Pw?�ND��f���j�սj;�����w&?��(g*���\i�u�H�xr�Y���ˉ=���2t`��=��z�\��*��]?wne�TJ��v��_�9)��w� ��g��v����P5X�#�֌r���U��r�IGU@�ӎ�:Е�w��'K�gD�p��$n���Ś	�I����Y��Q^\ �ۯ�뛥υj�+�v�6���J���ծ�T��k�pX�g�p���s���3�ɩtl:"j«w_�B>���o؄���eO�˲'+. (����]����k��4k�����b���6�uY?��.9�3���WWm��4?�� �z���; ��RO6���+�E�A�¸�mp۔�du_Yz�}��9�x]1g�!�/QD�rxy�o�Jά���7�/�yǊpY���8�6�:d]����������%q�䎞=���>���R�^��e��P�o�sW�pk�]y8TY�P'�;괽,��N_Ͻe�6��>�:���Y9f푀6�~�����������6%�m�c��o~��^�! W��-X�b#�o�ra.�*ФK�"&��E)g�K5Yf>�'��0�:��\� ��o?�35��"�Mn�]���"ߟ}�~��[ ˞��*��\}����O����,��i���տ���V4���i������ͽ��q�� �:dy_W~�� ��8|鷫_���j\u��zȏ�����V�����6�����9��}�t�4+>�z8��,ۗ"���g (!�|u�����ΕX�3i���fc#w�l�ņ\�duaLk�r�o:dlzY�b)��K������z$GTɟ4H��I`��:��Us��#��yd�G 2���[Q�3]7~��U�ڋo*�[��
�u�tZ��#�;�&�9yd^�����t~����]H�7�:�+'�w~|�B��#����ɟy��d�������7���}�s��k� L
 @.�E��IZ����Oe�{pW`��*�P�|P�n%a��"rǿ�깥�eL�P.Y"X�N6vuT���.սJ�z{�"+���\�] n�Z-�j<�����G�~��/��)����F��c�>3�6L ���7^�X��>�}����
���^Qpf���x-`E}�9(��>Vɥ���ʋ>X��OW[������>Yp���כu�4���PYU�:��X�^p�����}�ݥ��_r�@wc��'i]Yt���B{��p���+������oŋ�����_���׾��S���7�ݬ��'�Oʕ�*/�_��	�F����W����u�f;w�F�c��P��{��y<��*�|�E�Z+��%�F3+��6������غ&8�#mD�Y�g��{+�҆�RU��mv�6/��?��m�Z����2��S�pĺ�K�~l+V01`|���˜՘M��Ѹ�#T�*��×�q*�9��r>u�p��b�θ��#o�����f%�V��{��	���ዪ{���B�HG{J!����Ri����`U����<��-SU�U�-w�7 ���y����=V�N�q��ZsO��U���J�qVܐ4/���\pe�#	���Ǖ:y[����f��(�����x�����غ�	��}�+E��W��L[�wJ��x����V_����[��e3��������o6����0�N�U�}��/�#��v�
�*��q�a���R�f�zݤO�yfU�h-�{@n�{4�sh�����c�}�]����{"g*��L&4�Y��t������S+1�o��W�7sb�����q�'&����#YA�% %l	��&&o��yۏ@G�,�;���:���=� șr*YɠyF����|�u���1��I��S��|`�z���O}��ɉ],窟9�W��g<�lι�g<�I�|f�a���ʃu���� �b����-����8 Z�XW�]���Dz��.��T�9 ��߈�;�q⧱)���Z�.�e����g�k���ޮ0��ຏy���'���Yi�/�+�p=�����[��ȭҥ,S�5_9qPsN��-���Q��g��ϗ����|�3W_��W7�Ǭ{�v�2��_�ە���fUg�n���v�y֦]�+~T��׵[��C��[��v�����*~˲��rM-��D�nfq巊�g\�[�
�v﯄}%P��
`Te� Ŋb1K�����F�������������O���p��<��c�����W�>`��eO��`	�kV�ˢ�ʚK�g˼�=�Ee��D�(�m�V�,#�Ҿ��97XTK���b)�9�Ш�x�=���S����%��Emuڼr��픺��[[�v��� � Ve�Q�*!xu]mm�c�]�} 0���z,[�H�8�O2B�ۘq�b|�A!���9>V6%y�����t����h^�M�ӽ��R���u�� I����XQ[�8�Σt��ꋝm�ߴOZ����@���I9��7"?m����F��C�>W���e��T��rW b$��K�W⟄��XiŢ��?�Se��)� � �g?��͝H��nbl&�f���Z�F��6pP�}�~؝��˽�Ja��K>�
OU��xx���?���L�ɱ)��Qxϩd�dW��J����B�` 贌Qx�=�s�w��e�w�����qp ��/}i��˒�UVY���'�Ј����W\K�lN�z��r��5���۪�;e'�{ ~1t} '�憐�4���+�B2yO��R�9f~"o+Z��.���/K��'Z���,S2Oܧ�b��DL�o�)@,!�;��^7�����ٯU;S�mE╗7@�b��:�K�	���c��^N6q��:��,��ۈ�z��;�&)�6�[������ �������jS��u))Ǣ+t�sח���E�$��o�k~���)����S��ʐ��h�j���dŷr��ő�*� +m��͕i\l�
��k�����U�G��E��?�����M�=�k�=����ɿ+��y���V��Ly�v� z滂�.E뮍h	�^�|�U����f�H�vR����9���Q�NK�r�gWֽ�{�	�*�[=�Vz|�b�9)GBb���;��]���",��s���	���+�Guѧ:��3�pk�חLS�U���_�C�Se�J����=�%F�=�C�VD �/~�Pβ9p�zW�쳭���d�r�C�&QV�f�o���)-�_���1�R�z?�����,�P*}35��?+f�N�k� ��%����F΍5#>̘ �T��矹���ͤ�Ay'}���"��U�y��{����֕8����!��-���\�2�9�+$�]��=¼m����(�5�Dy�,^�c�4�p>�i:������g�q���!:���3~���c�n7a��߷I��4��sʛ~�	8*-0�k�ϲ��l`��l%o}���&��r����H[��li�3�T�N1`��6�/&ᣏ[���[G|I��^g��� \<�A�y��:y`A�&n�u��e��Ju� ���x�P�<^�*-���|��1��fc���'�R*�VL���]�|�>�}D���c�+W���R�p��b�j��B��XAI�r���}���c~�Os��U�
 �
�L�s?�?�8X�i+"�T��G`���,��江��ʤGߠ/ `]�U�>��7w� o�E���m�����p=R�LN����<�����V�E^??p��rq�p�K��3����j^��^�K��?�!�xd&�+�p)�Y��������{�Ͷ^�5�,���_E�#x`6^�JC���k� >��{i���z5(�*A�y�;�LU��m���7����Z~���&� �>4��R�)�,Jb����e�]����x�	t�p�b���7�|��>��Ӆ�[��$cNW/��V�Ŏ9���ʃ>���>`�Y��9�s����Ǎ�]D�c �7��iK.P+�:�����{��ޫ�F�Q]��x������?s�)'�e }����8%�r�����9QU��(}̎����?O]	#��u��tM���U}��J���1�Qs�J�+��rFD�����9�q�N�A�u�4s;������T�B���1(�+�P�F��'_��.��ZW�
���n\�XM7����ۜ��b���Ko��ë��R�.]���!�;��6�gRepӵ;/���'����������V�:U���R��33 4K�	�)Dr3�L��T�=bʗ���r��3��ѳX�|9R�\��]����`B��8��%������������C0��S�|7��_�Z��f]+]�譞4f�8���X0E�z���?x��NP�xU�����':��yo?�1&�h�pŒ���{oe@��E�V{����
r+��u���u��A��-~�y/�7��U���ܽ��C,i��K2B�V���"���QX�+ ��"��-���k�K��Vc��{�rAD���V�=�7#Z��3��hE����bn���u+8#�5+c7�]���v\2SPFJjE����z���{���O0�9A����p��~Ը����*p�jGe}rPu�{�5Җf�/E�v�ߝ�2�j�W
BW��A�bΌe�7-�|�M;U���˭]�(� a�7L�`��" ,	'�>v2��n�ʺD*�K{dy��n�[xgs�S��n������� �S5�체��pƚG��gf@�|�� <��o�\�� ��ڨm�@��ܭ��X�Ͻ4*��@�7��a���A~��͂d^}����}�_]c3�@u'�VdΈw*ow�p��k>�+�7�+e��>��si�ueH�3�g+@9�����۾Y�\}���)��k�;��*�I���A�*�b���*ѩ��ɂt�&�[��9�F���i<{��N�봨KPe��������Ue��@T�3)�si1�ʓ���`!�f���K�	��("v��
��-u���|�{!��bq�G�K�!�F��v�}�k�hy�֮/:�)s��%�a=� �X��0K�hy;f�^�����7� �gK�<�� ���٠�5Q�զL}�����@���ܙ)<#�ˏW�)Y��n�����˜��]' � ������#0�Ph��E���׀�N�L7k���^^w=�<hV���k�go���{�h�(�^��/�wm>�w#E�r/����ʵ䲲�U�Qa�;��O�����'\K=�O���*����?_����~mU#�ʰ���R��pSZ�,��wU���L���J3cP�����Xh�X������wl���
���|G�6���=�/@%�UX|4W�P�IF�>b��#ƟmJ�Ф�?�O���]ݢ�&�tݻ��WH��?���)�YGDx(���w)��͊��"��4Y���iäs�e��7�w�h�k�rU'|a]�a>� ���c4J���>v�����X
f���<�~{]V \N�����h������n"�ViV����۪C��Ka��8�K#�[��]��J�U�Q��;�>��}�ӟ����ۿ����'-��
Wi��g�{T�*���4��&z]B��&e߬�wO�+�F�~U�K���g�W� BȤ��ǧczu��V����~k�I��r#�*���t,C���������^x�-�0�hֶ�>#�����
0j�s(�qZ:H�V��Z����X�E�/��(Χ@+��p@���V<G_�$�C@&��i�"�̡(W�ϥ���ފ�~���]}��2�m(�>���s��8�@lQ��V��lM��n4�2|	���%�J�f�%�Ǌ��t�8a������]7�3���I���E0y=r�5���'���F�w}�9�>V@���g��t�m���Bf.ϥNK�jr���3ճ�|N���;�w�A����������_��W��E	1�L�ʈ��uA�9��a��f��!�����?��|�O��x����%(��rV��3RFZx�ϊ0����;�sCh>���(�8s��N�߿���R���Bi���F��/s��Ӿ!�� �}�rݿ��V����ڣ���V�_�^�ͫ?�����/��I�3�4�KP��>���X�?��_���?�~�b�e��^�����<�W�7X暲��*�WQ*%�� ���{�ڛ	n��̏Uй�~d�۫%%ߜ��=��ۺ��չ��Ǯ?�Iȏ|�#������At]��y-��g�y��n�q`����ė��1�?� ['\,�z���?���>�?��ҡ?�я>��gW=K� X�G�pE�7�����������lH�w�O����ǷL:j��>�C,PF�?� !Ju�)~�bL�} 3��7p��񧮕��������:蠳顟dv�A?�t-��ק?��?�%�;S8Q́��U��! �U�@7�%�k��og�A��6˸��妀�n"�+�v|�^�|���s�;�����H:��!�u�=���X�|:�e>�2{���������5<>Yzٌ(��si9����nH�=�ѵ�:	Ez1_ �o,t�������I�
 �������w�e����SK��f�_5Q1����:5��oN��`�����n�h���{sT�K��*�}��+/�\KPJ�P?��}���V	���?���At6 ���.Li��ڃ �"��C�&��ZK^��	ty�_��5���(S��(�EQb����rn<كΣ�Oup�
�pEq��<��_?�!�þ��f;:��tХ � � >"��D�	$i�;�8pЛC��sP?yH?!��5]�}���cV��c�uLQ�!�]X|<c��P�Q0Wed���o����&[|�=m�u�A�G�=��/]"�\P��k�@
䧑)4���H�娊1{���{��?�ԧ>�'�r/P�����p3��fN%c#�o>K�#;��WrM9 �å�z�57$��zĖ'���0r���f���At> ���.D~��=y�]/%�b#M� ���<�;�!]�G9eL��%��� ��;?w[��P�e�l\�FG�*��<<J�%�?���?����b�J߳ӣ:��t ܃� e�[�3�D�<���e�݊��y<M}㳛�\?��'?a�?K,����Ң��_@-�D�Q�y�8(.���9��" �nྴ �-�=`�~��b����!dX��G9 �A]��{�A�J��'�W.Oc�<a��؛M��,��=��J�.eF}�����v"�< W��{\R�ź݀���EA�8lࠇCX^_}���ԺR� 9�L}�I}���QHr�A�O�=�V�|/���_ W��tOgg��-'��{I�S��u⿋E��<\��C(�;���o����~�{�;����#m�����Ol']��Xտlf:���!V]N������\=ru�D��z��(;�[ƃHפ�h^��d5Ï>蠃Χct�IL��x�����f�A z`wҋ8+��=���z��B|y��p�h	 ����[��K�T���(�I=P�����d+}tM��:Z���!���s-�����~��i��~��y��E�H~��Ꚕ=/�eEi��p�A��p:�B�E_��H�}�Aŏ��z x�<�;�8!MD����A��#�����fG� ��~��h���pJ.&۽��n���3���`�p�6�uH@TJ�)���&O��<'@���O!t��h�!]?m9蠛�p:�B� �w�����e����J\��a�D������{��!,�l�/������e�����3��O^z������Gt��T	�pE��kÙ����0�QXQh�oߴ�<Ǖ堃:��{�A"�@�����|�;7K>u��ė�� #6�!�ܵ�eLvi{8��n�X�V��R�

���ࢀ���T+�1���}��s�݁�����+/�Va �<��˦B�V{$]`VZ���99����:��{�A"�Er$�w������P X���˝�' ��Cn��O����L$������z���ǀ"\Y\�q��R��~&��A��PW.�fn�kKX8��Ƅ����~�R+�o\�-	���s�A���tЅ��c��cXl��*�:`��+���<2`�q��G# ����7�3�S�O@�~����K���;��-�@��!B�A�O�Z_|�ŭ�p����⇻�D�����L�ҧ��Y�qk>t��� �t!�<b�o"r�ؗ�%��xFD~|���#�� )n(��۰�i7�۞y۶�-�$���� .��DNP8}�����}"�1�z����a���"N�S�	��M��Ƃ��*bCy2F:蠛�p:�Bt�}��tX��Mcn����~
@I�;]Ƿ�7���xO,A�%��+,��q�~��g���r_z����3�t?���F�e,�쾻�>qb�ڛ��1� ;`�G���r"+.}�ʧo6E!��Vt�	;蠛��-:�B��#*ː�N���ܚ��M _�j��+ߘ�a����*����Bĝ��_�������귔6&��X���P@��W��b]�b�>1.��A� o!��$B_:蠃nF�=�Od��B#ʳ���JLL�ұ�0b��%T�,D<s��+1"�F_�j"�o\H8rY�4F �n����ͅ=<��5A}!���GVY���WN7���Ϝ���{+�>d�Ѿ��s�A݌�x�A"'#�����@�M_�Hyހ�
�����'�G� 9Xa9����'�ܫ�����n ������d2,�򣟙�rMa3���QS�(�=���p:�@����Ӧ}$(3^���S�'^z%\���`��wO����!�� H<F�o�p��8���,n&��D�Ò�p��� R���DO����jǆD��||���c.t��� �t!�x�P�$��"� VV�� ���#R<M	R|r�a���#zCX��H�E��� �%�����S} ��6V�M��g�x���#?)�Pm"?F���5G�e�.��ݍ @�+Nt��� �t!ª�o��Ǿu�����,z}p	u���ګ� =���!�
Eí���#WQF8 �S�8@}��	�/ Ex)BG�������8�LsV��o���N1nuosS��E]������#���!)6��p�A݌�{�A$�s ��_zy�*�� �ŀ����<}u�yb��F��n�:���7w' .*a�P�|#�\����.
� ��z׻^_Ay��W~��I�T�m ��'_�w_9Y�5��� �p��� ��W����~>���p:�B���I��V�V[�en$��c��������r_g��~bG��"�!�PD?E�[��El.�o��������-�O]��\���a�67�k�*�bs<���O�;��~�괹������:�ft ܃� n$�~|�������n;�%���"��U�]�>[|a��(��7���	n@��c����ۂd���P��dr��9ɒ%׊���Z3y*�&Wňs�)����(u���jQuzVӰ����Zg�ڊT�o0���t��G֏!XP��.���x��V_W׍d�ys!u�8d,���A�͋>ǧ���'��B8��&��-Z,Pm�"�0���.j^�?�S/�g�{�C����v��8e�6�e�p�@`�+rl�Ϻ�yab�ɋm#����E�r�3�yO�.��"���*��a"pC���L�[O_��mv�]e,��w_E�@9�!���YR���r2��!�������+��_�X~W6��C:����u�FśI�!"��߅4��0�!L�/J|@� X�|�n�t3̇<���,��Yl�q{��@��f��՛P�����G	pԍ������go9�Q|G��(��M�oB���J�Oj\�z|��!Gn��wE�<�?��H�,�h��!r������J"|����zS��5�~������("�X��ƈ����(\����.�4��qhE,淪ׇ<$k��D��0^���N$�aO�/�,�ܨ�tq[�ɶk����]&�ӛ����V|m��%��/c�����o۔���cd
@��Mmf?|��7r*6>��� ��B��8�`���b´D��0���F���ȴ��va�]	#�ֶ��"��iB�E�;��]�.L�Gu�m�=\JV��r�'p���{t/DÙD������k��~����'��ӳ��y���!������y�R?
!ܞ�&�̝D΋/���'�x�X�	d��C�ʸ^�.N�׽���jo�M�J<~^V��а�r�8�Y��!K���G�L�^Z���ٽ���Ç��P�~�!���򁽜�J����!Gn��(#���m��[^����X[�H�-�jf��jL��Y�	f}��3ā�=��>��[�j��P,3	ZJ���h��&�)�)NB?|���c�⎱B��4�5����;�_"���*r���ldB8��&D��]5���ɰ^���H|�k�If�-��9�����VR^�@�d��WU #��Kf^��8_�$�=�K�0��I�-S�ܻ���gy=��m��
E ����q�*
a"8m�r�ܫ�=�I݊TQ����e^����ɠ�����mk*/�Eஶ�FaSw�븥	�/^K�5҇2����	�����1jo�o��G��0��B�������̷o��,p�M��g��3����/�?�@lz=t�gL&�|JLZ9�bb��"�8�|�����(�����%F�Q�i�*CQ�>M����A�����a"�1!���1�\�D-"������F���6{램��=P�=G�x�2��̭PV�(�ybۗ�DA��Ջ�d��y뱗��9o$t[@}�D.�pl��.QB8��&!KW<��t$�Eo}�7.l���:�6��Y\'"h~�;� ��Q���!j�f�Ө��{��A���}�� C+�'�xy����v�*�������xI�;f(3,hBd��j|C�!L�S-dd��V���;(@k5U�?���OF
�!G���E�zW}���FvnG���i�[�ާ��e'�lHw�c9�Y�b���ex�b��k����u,�0��0�pj�B���D�H!H���x��,�t�{O b��`%%J������@�7�A��ٳg{f�>�ʧ\����DK�3��>�|hk�üpk#�����ѣG5몍�b��J���E>��>�O�<)�4��3u�'<!��Ȋ�Dp<�5�^{���N�ů���'S��m
�wޝͱg���-�a>|c��W�\�8�<��y��g���'��FN�g�{D6����o���I���e��M�u��p�B��+z�>��?.�V��ϟ�a )G	a"pC���dk�˅2i�p2@7\���G��`r�c�[�Ha~�w���"1Kf�ZK��X(���j�pv~VP�����u�ð7v�P�H�f"q{��,%)|�62uͪ|ɯe+=J
7�#��a"��ݻ�]�
�E���2=>��
��f�XP9"�R,��D�̲����2�V�6�3�w�;���{��D�/l,�u|��2����n>�YaWN�%D�ae�nOy��L�!	c}�F���Z��B8��&��i���t+�/�{�II�T�'���F�^�ƕg��z��֔<D���#iJԀ�&w��>�Y�MD�З�K�sNX���F�i s����T���垕��-�յ���~C���D xT?�~�4���ux	b� ��KF����zӒwy��Ta><�Z\.ΫXq��
X�&$�uؼ���u)U胏���\68����R6��$C������������-�g!ܚ�&�%J��I�J�J��G�Z �����%Jǭo.�,�9�����ͣ�l�C��q6B�����BS�7�	@�����O�7�QVrhS��4z}�އ�e��`��7c=��"7�@�~��wu�<����Gc]�f����%�?��C��F���:o2k��n�t��S�B=��dۚ�0/���4�'ؑ}�͌C��������m�7��#7���.e.N��%[���~V��h�oO_�J4�a�?�"���;��Dy������7%"�&��l,�����Lj�U.D�^׶|q=�mͽbHF^BV�c���^�|���u�k9�i��ab�L�ō�U�T�pr̉��T�Ѥ#,�x����b%�9��f���DF��R��Ȓy�L��<Ͽ+���fx��
	�o����\�\}��O��:��^�I��u��;���˭��U����>Ɨ�p����ab�9E�H��aAC�C���O"w���}ءc�0/�h�
϶D�P���:��0�V�m_Ȣ*&����xWk�&�>`�,�(eIæ��jq9��߳!ܚ�&�m.��cN?~��ֳ~�	_0�^���P�we�� 4}���������_��8f�}�ܳ�4���lb�Bـ,�$R�'��ϊ�8�5-ؼ����Rڢ��K�����5�p��B��C�h����Ƈ��]�u
�
)�㋠��g�U_\�R6����,|� ֊��/�̮DT���Ax^m��e�ٷ)�^J	.·��ӽ��������7F�nMn���b�E���=��d����8O���	�oԾ�1rGq�=���ᾠ���ms�D.^�Xƅ~�E~Ԡ2f���ZJ��RGl�\����pyn8<$����Dx�M?�d����"hf}{t����k1�uq^�R*"����|cC�&b�7>�XS� !�?5E��oei]�2V�k��RJBc(�Z��[��d�u������b��!ܞ�&�3t��r]3q�Ǹ�"���?�6��=�
Z$��}p+8Ǜ�ʦd��Q���eÂ�i=P��{��L��{�r*C��nqq?k���@��\69��q�a:"pC���C�\\^�Y��G��}����{W5"ȅ��ƣ4���K������*��`O5-�	�-�En�������?�B)^�}�ͅ��+��'�؃�ᤖ�z]md|�`���=�����qdeaB\���s��O�������!�G�rdJ�o��{��6�4+b"�߃���yS+���R}�$r���4<�[��C�^]��z��6dm�M�kc�j9��m���={v�?W��`��D��0!��=?_�h�R�O&���/x�g���r�3�mNNNO�{W���u���.x���C[7�0�q�9}�s��������7��7�kF�3���z���
��������ANcD[�B��!L�g�\�0]��BgX��J���!��{����a1\w���x����ٻ!���pH�b�������[�x�_��P�5퐥W�2�?諾!��D��0��g��<��g�|(�g�0���x�B�zw�b�M~�)�Ͱ7�����1�w����3��h�ca�>�!R�r7�M방�glJ�#	6�4�	�ڐ�������'7��Q��bȑ&Ǜx���]So.�j�>#v�5*v��֒��\�T��I�^�RD�G�}���I�R��D�ļ�m�[��eߡXz�����כ��7@d�C���x��{6_Z�����%b��LF��1-�B���Ɛ�&K��m.�C������O���q�k��߿;  Z�y������˘h �ύ3JӐ�(��9���,pZ�����z�r0�Ǐ�=����YU�(=���Q���i��{��j/�����o�"X٨��V�dm��m����y���ln2�!LCn���M����hҽn�U�"��4���e�F�n�6a�M7L��|�2��.P���y�qj��tԗv���l!h�#�>�P�[=��~�Vw[�bw�H�C���&��)��/	T���|"�����^:���u1����e�|�5����{���)�C�S��Z�!�b՗CW��{�V���gmn��X��ud�7!"�}胻0�nOn���
��;T�邉���ۨ���G�C��a^n�d�w�,�d�6��o�	��f�Ͻ\�m��n4��(�jX¹O��oN|�f��3�׽pC���D��M7kw/S�jI�1�{G՗E�2D��	��(c`SB��Q����p{������p��DK��������]�bm��$�3��ކ0�!̀7		��"{Gm.5|1UӬ��d��CMF�*�n�?���c~���]�{k����J�%N�����m���Ko#6��"^=^%��o���+��&3��D��0m�[�ͥqL���G�mm��z�m*��n��6c��ܷ����(���YS�M����a^|��b�ş�u�r-�c��ᖌnSR�#��d�Y�����X�bQ�H�dtW'�X��b9����� �Ǜ�|�!ج84	nv������b+�����I�R���fo�&�]�s�li'���c[�B8��&��?G�,��H�Qwi&Z_7�;�ih|.����>x�,�n�T�Mη��j6��������E8me��2�Z�'���n*"�?m��8RB�����]�c#�[�|�ϋ��x"pC�wEhGz*���-��x�Ҕ������Z����rj:�Z���͏MJI����P_Y��M"�Z�};��b	������?s�������l��,9�\_�|/�w�B8��&�-�$Fu��6��IE��a{�-MJ䩩el�x~��Ó'O���zțT�"�yq�B���㮠8).s����qo,"��Rn�*�k�x�5WK�k]eFl^K#�z����F3���lonǓ1���"w\얫�^�	�� K+$Q�Y<�+�^�ګ�}��Au\����dll���=޼~3<{��f�ȸz�pA+(IqO[?�o�N���퇗�x�;��6�|a��S�Ě��ru��q�C�!�?�\E!LL-QX-���kI���z��]�,r�^G���\w[��ŦHx�S��оy��d����k�=��M�иk(�d~��h�gv��x���B�%Y�=��u��RKO��#�r�W{��BD=�	!En3�G��"j���r����O<��������^�����/_������A��Q��v1��w#�x��(M`�ӗ����:�Z[=�P�mN^��.�Q/_Pl%n)k�Y�K�m������g{���y	��q�:��U-5�s�誱Le'J��E��k�y���3��?�� �t��q��\ՊG�66���3µ/��'0�����U�{�OTe��lP���0�[��,"�p{"pC��=�s��L��z\e/^�(�PZ)I���@����ӂ���>�a^7���{℘m���l~xI
�������6�y�hkۦ8�d�5�PwZp��}�o6�!LC��a"|�+���e1�'#�{7�����o�¨2�C=�U�>��}:��ufQ�]���G�f+�Z9�KvX�~�����yn=�)#����uN]��Ɍx�;��RD�7��nOn3@YA9�|�f�/�	fd�;^s�`�q�o��*�G�juzR7%�=*?+�m��:N<p=�۾����48 L6�� ��ъ/��*Q`�2�ء|_lmb��q!GnÑ�.��q$)��Ő��Uw��Λ��i�%ӣ���9�u��C����u��⡸�\�6`�<�sd ��gp���u������E��U��3�%��b/�K=���O�{w�8"pC���;₠�D��ǝ�V����=�x���P�(̋��bGi�g�;�=o����P�C8�~�r����7���k�}�%D�}+x�&46D��t�*
a4��@"����[\/[`$��[oxq�����+�i��B�	޶���?���5��@���oV��oGe�Ƥm�3�$3���r��ֳ��!O��&����9��V�x�%��'��g�XXA��XP�9��#�1A I�����W���Rʇ<�C����m���>��6�B�~lP8�i�۸yi�ۍ�����#7��8��q�����4���؄����V����'O���&'o�v^�FS�@c���@�A=$Z��G�&3�hé��C�ڍ(q�Z.1?Y���I��}�b�����ʅ�#+b�G�4~��d\��"��G�q��՜��'�/]	\<tC(C@��ؐ�� r;0��[{nKۈ��'"~�
�Y P�b����	5���%c´dEa"��ѻ��� T���B��AOS�jq���,��()�+��N�g~ںK�g�g5�.��p<�u�����X��'��_����vQ��ߗ]���{���V��!Gn�Q#�1�5�.p<>�S��aƂ��N����
��q�κ��n���.n�K{�1?����ؿG�\�4���o^=^��{9B���u��&U�4�^ p��0�p{"pC��-�m-��t�(@pl݊bJB�ks���1���$�l@D��Őw�;.l�d�-�B�ڥ�L1����c����z#!��5�z��do�m%�p{"pC��<��g���~��G�.z��P�
Kvo~��D npN�N�ث��r����,��;�w�����o��F�>��b�7\O&C���w��T������������c��S���r]�K!�ۓ-C���zWu�5�����.^�)��!�����3L��Xnp��ѵg^y��"ZONk��X,�}�[+)^Gf8���דUوx�$Pu�[��}�'2�VL�fXJ�N˟���'7�ps~��1�r��]�d�X��y׾TD�ߒݛ��T�XV���H�"`��;|~��\�O.���ݿ7��n������;�Tm�v�YZ�8Q��{���k�����O��Gn'�!OV�&�]�x����!����M�("rh.#;�
1��Cmv�X/�U�:�9�f8 �K�*���Y�v��g�>h��jl �ޓ�o�sxL}j��T��/^��5���fTs���D�c6k-�Nشu�U�.�74oN�gp<�s�8�ya^��/�����ZY�pi0<�ſ{�	�aO���CA��6)l0E���y���a~������+ï{�<�+!���a"ڲ�Ժh�#|��\��>݌O�?Qqh�ñ�oj��D�~�Ղ�Ki�y���-�nڃ1��L}@�*�~=�Q'�����M��S��uw��&.�p{"pC�D	Bď)=s�S��D^H̪�O��]�\�\���F+^n��oPl�NNk�Pm��������y�� ��gq��`���j'�y��^�uױ	a"pC��:uOK�.h}H �ˊ���%����zn��ŝ<�J�f�P�1��&j9٬�^}w�H���)	1S|�����'׹�u���P[��>���a:"pC�?^$���x�2�H��nV���'v�[�Ǟ�ķڀ]���o�u������.���Yݐ pՠ�&4��{���}H $��8TG��m=p9U�:w������e�u�z�)�xZ�p<�!̄OB"ksH��t#1�������J�<���U�U֝�n�c{���=A�亗/_��
�y��M6�n�����̧rmr}��,'����#�������U���'7��p1�#z������d3�&�f����*?����*{�x�����;lx'}k'�"�]v���]���gJ��I/���e(D;Dװ�/������Oe�Ј�QD��0�@�Xt�9�x����]�����%���8�)§?���;a�E�e���Ov �x��<�'�������v�*<k��K������ի��q[�'�!LBn3�@�G�O7*"g�a�l�ӪW˭ȑp���"VBw5��Ӓ���y�������I����d�rL}w��5�Mc�����=����Y�7�*mQ#�>k9�p��7����Dx��-�<��6ALG�9�"r�S����Ѐ�d���XQ\T�����2}J���ojm%�'���V�Q��c$3��.T�|�6���
�f^�D��S�{�]��������5����!LCn����0 ��7�q��g0�W���������|��a��~�������"z=z4|���=[8�>����M/ա�������Ђ[Qm�v����B�S߼p��x�ז�<���a"���(���#N݊����K8&Ղ�"����/��ĭ��%Nݗ�x؞�P����F��!��>�lj|x��8� R���f�5ָ��~�z�}�.�Um���E�����0�p<�!�@��\����~��ǈ�bv�)��>��j���>���ZZ����>*�I����'��b��m;����Il������h�֓���#�ٰHЪ�E�2�rnB���f�,VZ��nZA������r}�7����ڙ�i8��:�z��Wi�2����vm�h�/'����qx}�j���Џ�1�ڤ�����c�5\=�w�\.�rd���\�!On3��xh*�/h���1͛�D���u�����͇l��\�L��\���7��܈��b�6�A�~����G+�ֽ�}P���ml|̳�?>("��x"pC���~V���ON��6�̭}���lO��#q"3n�Uv��nL�}��q7pmz�Hٴ�������1����u�5c��n���j����H�̕�Ū��jO��R���q�Ű/d�$D�����!q�//9h�ꍺ����B_����<��¶�ŭ����q�����x�76a!Onq#S��ܟ��˶D��ή����6;A�'�����{�e$j���!����O��Ļ��\����JT�u|�.n�v����U��2����F�׽�f��Is
�<���9Eh���F͏P�����J�x��!��ߓ����յ�B,��HF�?���&�6�\�~��׫}@0�}L��6J���$��!7�`���Z����i�;�g�Yٶ��œ��L__|ӎ����M��B����*�0���0?����^�S1�߽���Fױ��+�ds���˿<�#�3�.���a������T��]V��f��!�C�������7����}�g�Q�!v��wB�&��"BhdH^��{��ɍ1�4����1k7<d������qD��0mM�7�
�����'�u�g?� &{ۗC�m��rq=����F$>��P=/�+����~p#n�J�Z�Y�.�kl����'��X�:�����$��_6����B�=�!� G��%�eO�-Qh��L�-�{nLX2b%5?�,���]���y���P��P����cJT��d������⡿����<'���]�]�;���Z�z[/g����Dŝk��#�¼$%�p{"pC�-T��h��,�"�{V�&��{e��v�ڇ���;�콛���>������B鉐����LKK��U(#` �6%d_و��V��z�fЇ�����q�{jsٴ��U�C���D��0{�Ywv_m�	��sy�8~\I�á#��Nlnn0��wؗc�1$,����#?�@�~��B��U��@�"|����J����óg�����.W5�z�>����n�s�x"pC��C�K
�������d�7�뾸��(Y��z ��J��U�L�c�r���Ly?�!񣌭y��?^�8����p<h�>q�p+@��V�IL���!7��h���ԅM;Ũŏ����\��ݷ>�����Gֶ�v�OY���������*��"~���� �cs�D�?�PE,פ��RK��u�FE���+0���QwO{N(�8f�0��2��8d��cmf���_�}O3��>���.t���vb_k�������Ԏ�mk��������]��A3�ó��KSx=�7�)`��ĵZ�m����'7�p�/����v��v1�uғ�s��&k+Xh��ܻ��L�2����l��w���ꅻ���jS��T�Q�Ac��0l�8]��>tMz���s�CP��#7��h-�|��^�n�e�6C�@�6YJ���9������W��*�=qm?�?q[��v(�{���;S����\F���[3�F�|/x�ov(I��j��N��&,���aB�5Ul��d�SR����y����Ξ��i���������l��,76#��q�^z�^jo��f[�\��l����`��iM׽�����w!�?����D��Q[G�A+j\0	���{�<}�����ͪ�].j}ei[\�e���'�~�Z���%�e��
�B)���7N`�c�]������\�x=ͧ��B���D�x��E,�i1cd��۹�4��h��ɚȳEmg~�wŠ��zI�4�w[_����j���\�P�!̑���*�O�<�����ŋ��X�0/^.@̽.כ=E�}g@�!6W���0TG/[q�n!���U�DTѩ�l�����3=��J�Q+;�5rK)2@���S����	�A$�La���;u�^�6-�fJ�{��A��e@@�b��Tl\���e�W�mN��};nt../��3��i���ƅ�#7���=�2wn�U���.���b�&��J&��l��1y�n�t�fD"F�t@&�iX�&ϩ&wy����x����>�ה�`�������q+!���|�O�뺎���`��!7��p��"���^w�Me�RRey<kT�{�ok߼}s#���<N%n�f��ի2�����|�ƨu]��ѣ{9(�s��>��j���M���bۦ�K�R3O)��s���	D�;2[�7 �p�!L��6e�"s�uv,����,��}��m� E���-�t����!��῿����^��>K"�f�6��H����S�=zT��g���f���`hq�߇v�B�=��2��pC�jq�)�;�ή���4����χ� x��%!ꂆ,,׏��n��A�p�MƏ����N}���µH<נ#KKM�g{���r<uAe+�����q�ٴ�p<��2�`B�4�ظN��U�IC���V�!nUwK=�^���Ò����������w���������?.v^�����Wexoi:#�n'%Em�p�U����ڸ�T�5��ۉQ���A���7ʒ���dU�R��)K
!LCnq��dk��Za�>�M��H��c��Ԃ*q#q���nF���ͬ{����������@Rn9��f�}�1�d9�vO�0?^.���E�$�~� d��63�{���_߭�n�g�v���DP'�Xт�L+�9���<���!�����w��<�H��mN>��ᣏ>*�epِ����m�A�L#����z�ӓ��Y�����v��_oĂ�F�j�w�-+���ހF͵~��77���a"��b$q���>���.��2ň�i�]�z�WS��G�������b��	\�[�W=�WǺ*��m�?�G��2���%ۯ�qg��a^�X�'���R�����6:L���;��4���G�b٬�0�!L�O1>Ё�T�Z�t�q65|oTa����9.p�G�=���������{�:�w�= ��C#{��v������ImJ�5n)槵��T��?A㟾xU�t��zeoe�w���>���Y�gj��e���D��0!��)�-d_A=.��[��dv�~�k%���M�süP7[����py=��f$��n=N�V��
X��e���(g�U?|��)?�:f|�� (�zL�+��6W����$���J�|#KY��!�nOn��@:r���4#!N�գY	��p�P^��B�\��ĺ(�n��������ɝ��A,1+�����.'�X�G��$+���[��#z�)j���3NB���D��27^�G���3��|(��D�vW�ت�S�V��:
u;���6w~�P�p�{�>�
�'����\������߸�a�c^B��VP�PG�7)���`�^�;��!7���1��\�
�%�夾V#_��H��1?���S7�_�����"��w�ŏ���F}���]�yG�u|o�5�7�G{m6����v�Cm �7��/P[��HpM㏭�O�!܎�&�.ǌn��&�e����h�����, v�Ӎ��gq3.D=�2�/�5�XG1����j&�4lnd|C_ܦ�2ߨRc͵NF^���=o]��I������0�!L��(pc��p�L=����u��%�.u���I���@��'3�F�}� ^E�l����M���{'�2���=׫ۃ�_��Z��l��%"V7�'�hK�|�B8��&b\䮼Q�E�����iA���8��k<xP�#�ۊ���!���2�d�b�����m��!�Rư����
���㒠�*=r�c���k_����@c)�1��4��0�!L��_�ŋ/~>ފ`Ѣ()>�ȏ$i&�I<��§�-���"�i�}�2�����=��V�`�%�gߌxV�,|}�f�i�����n��}ӵx�:)��B��������%�+�{�ר��6����n,7���a*Zش�Q��ϭ.�坞�VSxM�:��c��H�������a^<sGÑ�q�.Zok��g|���Q��M�/�H�>{���Y�P�h����;b:�ѿ�:�{Q�%n�o��)y�&���a>��_��7���(b��L�p/͒�Y�/���{����?��]�&�L�g}�ץ!-�	�i7��P��M�Gp$�nN4����Z�6Lmv7��>������Zj�	���J-�2�ʰ�gIؾ|����0�����a"pC���f����=-~�������L�bH�C����
�Nn_Fqr�u�t�#pٌH�
j-)1i��|��7� ����b$����;g���b��e�c}9�zL�����E�R�D���6�p{"pC�2yx\��E�^\]��J=&q�]������|M��n��h��|����~�#k�-S��xicB���_�����ě� "zD��� �*7@�*>���(e!��ll���z��i�ۂ.���\����nOn�W�5�{.N����ѝ�{�$���P�b���;/3o"c�x^2w�NSNr��{��pK*�,]��U]�dU���Hʵ�C\����qL�����{9D61!LGn3��G��,�G���/Mj�t,��>D����y���O��_��c|��L≛1�ʭ���fG�%X��u�@}��(����s���F��->��%J���V?�q�zm���#7��`��"�$#-d�Hq��u��/hq�0�C}T/B�&�V0�y�����	5����g���� ������"��N�Q���-R��<��ͧoV�#�|�o\���x"pC��Ct�)&d��3�,v��ڼ����!����_.��4}A}p�.�G�0�Lx��z[�s�������}A�Pߙ��>��T���B\u=��G�#o�'7�e�2���+h(��=��'7��`���l�gm�"��)I^{��D���n�j�a��Z�G����w�Xa�Oi��u�f4�0�`���̔5P��%(�q$>�@J�*6lP�l0ǫ��-5����^��,��q�A�Z��9�i��a&�������"�/GẾ�ﰷh��c���QG��n������$�� �mØ>O��=���L���цC�(U �NV��P�]����#�y=���!ܞ�f����v�+ ���kry���CQ�/ޫta�>PZB-����={m.��>��@�0��<��wJ��%'*Z��j��2�*Cb�����/x�����ɓ'u�C;��:���D��0���"D��Y��}d�X%�bI�������2�e^ɬR;�z����(�tL�w�7@�WD�>W1��b�s �,:�MFp+&��r}R]�z����Z�<�WD�^/Q+7]Ӟ�%��!On3�fpy�{�����ؒl-���Ziva�����l6�d�XPC[k����j��y��`ljD��ȑu_�dW��>z���R����\mv�ŋ�����TױoP�3Sr��D��0!n������z^�W,�vG��@���d��A{�0?�_S�JF�������__���_�\7�y�	��m��%#����ZC�b�&���\�
[���n�F����|J����!Gn3�vB��I�	��Z���{�&��2�E�cne��A�} �Fl�JY�\bJCY����ժ�Y�|d�j�w�o�/"|��Y6��T"�'�	/A"�<�=�&�ǪCJ=�0)�!L�(e�[uym����yw=MHz��Hu�g�_�W��Qv���!A"�C�@��1�,�^�%V�����a���;���JS���f�0/my�[��jR���+�v�O6�&�M�6��5��C�� V�˱&���7ID-S�1d���V���P�>��>��߽D޷���L�].���NW�=61��^���Wógϊ_��/��L-n?<��e@���5���jY2�4��A=��Y�^��G���#7�`�*G��u3�}@����nq��ӏ9��0��/>��1����^GK��A �C6�-g9Ԥ�~�ĭ⤍�IϾ��V#\���^��B��}2�!On��Ģ��op�(�Y��2�JG�O2k��B��J Q��M���>�m2���b��*<n�J�7$���6�f���D��0!�T�0eA�����P�ZMGH�+������ R=�G�κ�~y���}qY�55yǽot�p��<�u6!n�[64�f�g��:�a:"pC���y3�gjD���y�,�^����e9��\/<�g��f�m2@�P��S�2 �\���&VlX?y��T�>���/��һ�JFC���f�������f��=�����7��Qq�ߐ <ɺ2��HA��lD��	�,��6k��o��+�\�൙a�q�)S��)װ�[�"/i
!Gn���n�:[�U; 2�X&'����H��oh�,���߽b"+/D-�P�ZxÙ@0!j��]D� |'<���m�$p5�Y1T̩�&NmC�_�.V���oOa��	a:"pC�.df�4��?��9~&����>v}yݵ��7���]b���V�Mg�di}R�g��L�X��p���G�������<��c�k]�b/F6�����7���aBX��԰��N.r�1��	I��͵����ˋڹ�"+��e�G٪�l� y��D�D���v̽��[ճ�a~�H��q�L�sQJ<����-�kܛ������#7�	9t�O�pFɁ7����x�zor���5e���{����1���:�ww�c����]q�Jܲ�t�o ��,�ŝ#e�����1%n!LGn��;�]� p��mzW5��?�7�����fm��������-ʏ�E��3���Q�~1��2�n�{�����e��~b�u���Z�#7� �zzrZ�|��O���1�>��s}��Z�pw����Д+��~@�z���k<��{?>��ӯ�����c<�Rv�����p�x�ѥiPqT��b�ת�!�&a!LOn�&E��b�L��*Y(��3�x�z>�������D��馿{M����ϭ�^G��u���Kl���7�<������?{��^�!���TAlO�t%h<xP�u��U�)w��D��Ƅp<�!� ���m��w�@r�)ރX"c(A��}��)̋O�C��?*MH53��f3�S����w��x�l��S�(���"ti s��i�G�:l�ab�5�n��!�������4�7��-.	���V�v<�6�+��PV�3����|P�������d�Y{���J�x�·tx�!��m��)��{e��Џ1>k���p7ϲ�A�����}�6��h��s��`[�B�Ӊ�a"\`z�U�G��ďw�Bl����>��i��y���{�������eݔx9�{{��B�Fl�8c^��� ������ᄸiBV�/��W��W��f��%�^�٬�p<YC�/���~�G�zm_+r=S�q�[S	���5������f�_6&�(�7*�%���.������V���i���C�e�x#:2�n�cB���2�a��{��ay�Np���oC�8r�01��)��Q_I֕cmčOKB,)$��q��A����xm��F}�[|y�A+��Sƽ�R�P��z��}{},�Pn'g�
�c�V�L/Uhi-�|P��������'�|R05؜�����^BG��Ĵ�"d������K��NG���.����>w~�"J��L/lZ��"p�\�lzv��jY.���NϪ�%�������_�1y�M����F��@���&��c���E��������O7�i�U� DKʰ����]�ר$A�	���P���2U��	�-����:�����n�[�[.��cy�~7c(U��n��>|��g_���r��S��I��Ai;ٌ�5&>�����As��d��#7��Nh_���DMD�4!����qev���ѣr��j,���pbB��z*F����a�XVk1^G��>�|��Z�zMh�������ȯa�vk�d|ٸ�PZ����՚]}t���M)J����k|�[Eᛊa<S̄D�����Є���K�8C��YwI�vV����1�2��k��CFK��j;��P��C��Z�0�G�덅���x���4Ҽ?�p�!L��Z� 8��񼼇E�x�>�C��=��l��_o^WG��ݳ��j��;BL�����5��"*��ϕ<��į=jdݧ��-�f��gp���|��Π��'7��p�َ�l��O�?��g��AS�K��En��{Fܺ�N��M2�i���6��m_���맿��o��w�ݘ&�o1b�ZNch&�,�7*^�䍥)A
a:"pC����m���#p�D�����%j9�t�\N5�i���3|wF �Ǜ����{�K�4��cgQ6=�Zl�����yF�o{"�g�A���Ǻ��O-��@�a��C<��̿z�/J��~��o��B8��&�l������=D�����D��
��յ��g��v��/�ʶV{�{��%�[[�I�J��ڭ��x�]��av�\O���!P� ���1�&����=��|�����ٳ����C���&�P&����U���ڋ�E�J�!�3�m�>�����F��1�L?���]7��y7��+$@U��l�b������?������� �)�E1��2��Җ�tD��0���������"GG4YW�R�p��c�׭����c��ϲ���T����pzvZ���4e�LjV�; ��f��O�;Ԙ�BL�m����c��2��)T[k6ӆ��/;��JZ8JB�=�!L��37����'V����E��"�5���Ìn�<�����2rzL:�wa5
��k[�ۊXď2y�&�%�]Yy#`)K7��Xf2�[~ᰁ8�FP6��5�2�ӓ�e,�a!B8��&�����W���W����1� Ҭ���(^���F���|C��e���..Y��L�j��Y���z�3�����_�~����w��|0��'?)������n����<Z����k苀]\{\�1!On�#<_�zUnO�<)��$�Ts'����G�Yl�B�|T�F���3���/����x=f9�^n������z/��:��;T���O�b����O>���F@�;�6�lrhR��)Orb�4D��0�[�G����1-h��o���G�Rߧ{�D9e���1"�������شs k��T9�>;-�e	�]�$;ݻm\������Q�~�Xf�\�,��R"�	t��"b��q��l���@P��w$6a!On��F5�Z��t?T]��-��z�6�MuP`l+�M-]�����ҭ�-B�6]���T�3��Q�d�߼�v�K!p�1̏�X�~�psm��ȕ��ͧ�y6��s+�4�q}{6?�(!On�c9U��H����|[����2�T�ˑ5vqo\讶��!ğ�swP;)�Β�g�RD�N�0�d���T�[��z�}h-�R�p����r��c\���e4��X��r���W2� �݉���B8��&�g�K����D�Dl����%2;,|�窗A��ъ�v����xA����z�`�8�7mcY;�#��g�}��ȗ���S2�x����F�:xe�_��X#r�Y�X`}M�ٸ�0�!LVa����拝;/��2�?{'>��ruw0��r���J��]'�G-&&�]\���m-�ۃ��q"n�3�sI������-XmX.�eKݽ�ͩ�O��X����ktb��k���ĸ�i��{��u�K�%�|��s�܈�� P%x��	����?#pK��ŵ�F;�Χh9��!ӎ����s]�\À�5�p�^�ph�"X�c~(��Dr�x"pC�/Q��Ƣ'�0-�����K���Ͷ���6ۣ�do�����"^|Z��̳���~)B
�;��-�&��@㘞g���8/pR��\J(A�9e�_�|YK��	�x"pC��V�r|�'�>�,嚠L͡ѯ��X���˾����\��=fd^��$k/�#���).�{��ĸ/~���Ǹ��6<����|g���b�ϳA���M�a��C�'7��p�ô"�T��X�J����V�.�VW "�퉼C���Ccz#~���>��K�q���جx�<����<�UF@��/ʦU�Bx䒥gb���4PO]�v���r��u�d�u��%7��h��Y�U��?��7�a��J-�j>�Q��k>��d�Q_|�Af�4��7��nX}����U9�>b��FxSb�m�*5`��b���ߗ�jm��%˫��/�����ݘ���!G��&��i�@QH5��a��d#��7Z,M�Y�S�G6����,_臗���5
'�����N�mtQKI�V���"�zk��6�����~�ʗ�℆2w�!Gn���ZД�Q&�6��u���B�"	a�����u� �� ����5�W�Ϸ%>+9��oD������į��7���)�D3]���zI��c�C�#7�	�ZK25tX���1�Z]es����^���Du����ѥ�3�Mw����	��r2��˓e��!���d������/j������֞�y6�悍.|F���UXG�����,"��==G�&�-p��R�Ǭ�:�a7�,���Ͱ���e���Oe4o[�@ݮ�n�C��Ф�0/.n�7��t3���ڐ���^��2�z����[q�0�p4�!L��@	[�U-f8$(CKǵD,K8ʔ�Q�	����#��ꈟ~P��"��\���Z��u|�){�6�G�����&�w��(��q��4�Q��I�b�U�F(S� (W�ߝ����B����x�/en���3YZ�4>��U��L� �x~��uA�2|�.p=����ʻHiuse����Hk���dщ	�b>*���oR���3����C@<;L�Y�8"pC�?�t;(�  ��J��g�~䉗&� ǚ�'��^�P?����������?T��\-���7�;�6$J�d;H|�C�g`��rͲ�9;=�~֌in��G;��w��P�tD��0!�\�b��129,zB���ǭ�����`�r����B���=3+U`���b�^Q2���l�J>�.��� p#�=�tO���U6�׫,��������Eu���4�w����!ܞ�&�m���kn5������F���?}�@Q}5��d�uk���װ�닛#�׻��j=q��z�<l�2����a���9#�i��a"Z��ry���U����}�gm�N���	G��A}A�"j(%���:�*n��M2S�V?�l��z�^�ufp���~�wN�7���<m��m7���w�����E�E��p<�!LeC�Z\-n�!��TR;��G��OlqR�L��������z�-"�X?]����Ѭ�\�[uas��:�����j��X��eDL&��z/��^��+!�i��a"�!��޼}3,ί���[_�NNKvQ��M�϶W��~�	)B�n@l�9��ޛ���� ���e\�r���k��6q��؉{?����y2��p�9U�T��z�az��ݶ����!LCn3��$�a,���!xE�?�����F�?3����Zh�ʓqo� 7�k��z?[G&��t=����{?�{##�7Nhe(�������Zm�r�{s�HF7���a"\|ptI��3�j����u�����B�U6�'�\��
��<$J��QʭǱ���FJݷ�ooLǊ'���H]�t='�x`�Em�h�6t�z�Nj~��붡4q�x"pC��
T/�B�kr9�dѣ�����/�؃id�uF����x^�\���/\�*��� ��v'� ����>(>lR��9]!��`߸��u�jʌ�����fQ!LCnAfO����p������5|M+޴$J���m�|�E�/.X[���.��fJ5��,��%nR5��;��C_t]���ի��G̲��Lx�}�����r���n��B�'7��8T#���I���,W$�>[��Q����B�γ���oBN�Nˍ	vz��L�����!���Ƶ0/%c��ϳ��D3߬
���>�7=��7,��#7��84||1l�
BFc[U���$�pK���Y=��H&w~<#�L};�����r=lVc<��:[�W���2�4,������K�a�_{�W�����A��r��R����dwۉ������x"pC�?^t��8�<�}/�T	!J�JF�m�|ԫ�����O�d�u�^���cZ�_��XKa=�wF����n���vm�ͣG���C�SbR������L;��=4"�p<�!LDk��A�Ѷ\o:�,�^O&���ж�?ü�DFFO�-����&��I�lLظ\^\��oPT�{vo۝O�,q�'^O�8)���.��-�*Bױjo���!���C8��&�m�Z/S�-�ڔ�����y��S��<�ӭ��7;��@����|���[���u���Z��Z�F3wZdo��Җ �D1S��b-��FE"1�׸E�v+d��u!����Dx��S�6��W�&��i_��ܓ1�����	��{AY���n>�WxyvrX�y�dwח{5��w�]Zl"�i�&N�KF�X�z�7<\��!���a"괲���֣���.k�[�|�ouT�	(ol�AI�q-�n-��f��̵���[�F�Æ��1|��7��})�4�����67���� (-B�"�)K��Z�)򓟜Ƅ0�!LD8õ��3��=t鵺m��="�q����G[&Bv��=��MEd��.����g���|E���ů�vr�6�8�(���eC�LFS!'54��{���7���#7�p�{����(2>>�^���w�����Nx&[������S����ŵǪo�ڍPbݗ����:��W���!�6��wL��y1>�!LCns��!>��Ű�d����\���bǢ�ȅdo�w@<���f��j�r��J��J�
	(��3���vjZy}b��̽��c&p�QiA}#���7�}?��4@H S�B�=�!�@[���Tf��Y�0��)Vm���*D���Ѐ���f����p��__�ox&������ĺ�V�x�.����}r}s��v�����Y��x"pC�?�D�j��	H��17xfG�s�nZq�?���̜�a�ضv`.p��D+�BܷZת7��ee2!u��Q��q�.�وiN B�'7�����n���i=/ی�O��Ϫ�lP��5{������>n��>�>o@�*A��}�봭��:ib�qn��Ϣ���ǵ�n���D�1��*uS�4�zX!rtlMG��9,�X
a�H@}i��%���&G�������r{Sn���_+�����+����S	��O�L{9�^����D��0�Q�gw��K�>B<~��N<"�Ǒ���@'���;ޙ�h��g����V�"^>఼�~G�~M6x��7F�oExr������-�ĈѼ����u㽔6�{C���D�zw�xia��[)3K��D��p^��=S[����Q-��u��C�]Ć,mɺ�����7�й5\�^�G�tz��~�gf=��nZt��^�^��SS���+��>Gc}�7@�%K�	!ܞ�&�k���z��l���P���gt�gO�^��7�E�/��{�lnq �5���Ǜ5�l�~|�c�x�Ҙ�ߛ0?^vpȪ��	���՞՛� �_S�;��n���Ĵ�[2�:i�ud�8����y�'��z��?>�=6C?�E��E6�u��K7��w鳹!3���	�ܾ�2�]�g['-�1Ui�����mP�(���0�ſ;>ʹm@!܎�&�����{4�����O_�<c?}�=u���c8D;0"���>@͂�����M[0��j��s�#bS���-�M{��@Ul؜z�
�x�vE����K|LsNfB8��&�Ŋ� |NON��j�H� ������=&���w4f��1B������|j��q�M1�m��72��G���]���[�\�ʾk��&�$�f3�@�3��4D��0�z���6W�R��8�8�b�cR��R��E8̏��"P|�ǡѬ�a��~%,B�㶡���3��-G�ڤ,�]Q|ܲon��cey���1�l�ÇKI�o�C�����D�'�١�5�޽ͽ�ñ�S��5������ywN�e|ډg\��{#��)�mSR���D�E�_�daK���d�:�zg)	U�GW�
�B�A)R�x"pC�	?n�B(��q�9enZ�w�]@y���1f�5��T \��-�x��b
�>���jpY����A��Z�
��R�p6���zd3�q�����FBW�j~rB8��f ��ƘB&��Nu�e}���cUY\����N�ە�q�Z��*�K����]�� ��q� {����Z{�)���	emI����hs���?���ǅ�(�0�!� vO,T�*K�r�iu�d��}A���ΫW�j6H�z�	����������Ų�_��e3�ӱ�fg�~赞�M�/lD���!T�1�|6מ�|/���{M.��O:�|����0�%��!7��!�#��{��+?�\+)2C^��b��R��z\G��Iщ���~D�7�gpEkV7�ˆ�}�z=����lo�@苋[\䒹��;��OS�Y�	��?y�N�^66\�"��x"pC�J�P!l=�Wj+���]�k�2�����>�]��0��0]�^n���撩u�7�G<+��H|��;~�á���]���9�c��YT����q��� l�׻�J^��f�WY�F��D-�z�#�����Z���Tg��Ex]�7����c���������~���2X��n
5����ͰW�˵N� �mS||s�8"pC������,��E�P��>��,BW���z�gm�B�1�N;_cyo��1svzV��[j�jk�6c�n ξ�$�c�ٖ(h򙲸�7�ia����4�M�o�r=�p<�!L�[9����f~��x]Md��z��z4�=�(W�/�(���zMe)-��YzI�.�=�w��l/ ��!���A��h��w!Z����`��¼>�}�9ݡ쁆���#7���Qz�\�-������Q���zM�{qr����?�/t<]b���ެ̠���n���R����_62Xą���R�r�^�L��������x����Q�x�ַ^˹�C���&��)h>�X��2�� ��꼖uX;< �Û ����b/�14��C\)?�hb�uּ��3��L_����f��^�.X�ʮ��Zǫ��1y߾y�fx{���gI�Π��!7��h����������,�5��G��=���n��R��ZV�C���|�X�:��bXo��q�b���N%�a|�����`��Ln?��M�#�B��~����60�_����Jf_׻nlz^�zY�gt�(q?Je�!On�"���ն�!�׍���/�y��E�	��%�_>7�/ڼ���n�O�pq������v��bB�GYA�ّ����8�Q�p�.�}�)�-�8�$�+�޸�M���w�V7�W'9�m�;B8��&�]�}���Y}|�;,����7���C�qQ�m�2�mHp��A�,�DA��q�n>�C�ɳ�^����~ P��կz�Z�k��O��&T��{�`�>h�����z]���#7�x�{��l��~oF���fس����~�x]ߔ�^�:& ��	�gϞ�F2=��#o0�	W���R#Oʹ`��Y����m�x\�
~�a�f��]�u)s!ܞ�&��?�=�[ !d��u����:�~��U=4�*%
�@�R:BY�������j���~'gY�I��<��B)��~��H9my{^���a��q�Aԭ�\ �ZF$kcC)��Y�%�i��a"���.n�񠈗����ru�g!�
\�F~�Y���r,���	��'>r�m"�5׋�������D`�׸�Ln7\t*&r=P���[^t�$�͍ǎ�j�f�]�z�x"pC�����%	�qA�X��*��Z��ѣ���mY�V8uh,��*&�Z n�@1�cX{��2ry�mF�g綄��TC?�k��mu]SJ�Z[�F��*7��n��nɻɅz�����'7�@�R�Y-��Ӻ�S��3�,��'ĭDYC��OƧ\�����i5|�s���EшD�~��nr���i2�_W�~�V?qQ�Ԑ��"�	��Pw/t=+sO�Qn���� xX���[�aہ��if=��g���"�vWS���'+����8�vӁW��Ѭ^��f��%l*�g�6�^���-�n�XQJ�͊ۊA[v�FU�+{O�a;-�p{"pC��t_��]�\��yM��"�pe��/ӳH�.#{��B�3�.Py�g��'��F��qjp�*{�U���>�/^��(E��u�4E�=��غE�^��(1��S�q�tD��0��v�.�P>�ճ{�}�^��čDX��s\ gQ�O*�Z�Q����uҔ�;����nS7�/�����c�d����)Å�6e�ˮ�'�V�cP◍.�|=ϰ/eI�>�i��aB��V�2�s��Y;fړ�i�1DS�hZC(�Q;-�O=�>�Q�;��5�t��0Fs��e��(d�����{!{V?̏g��&NM$���Z����I��s����3�γ�!S�A!LGn�"���ek�����
_PY�� z�u������ic�quw�t���y+|����E�w�~K\L�E�lq=n���o�/|b���ϟ?�N<�w������B8��&�����wF��y[��N�Zt��ʢ�3?�L������Z��B����p�����ի��⼈(�s�����S���I�d۽�?��~mx_�xQ��I�
	!LCn�"�u����Rx�R�����$cG��#��N϶N�ᆃB�1V��Ʃ)��:v���ZLD�����9�}������k�W���
�.L���m7�\��������\��8.�BV����e��DD��01�e�QL�,b4��x�6�	2�mÒ�&�^��n}'{��{&S�����0��kr��`��%*�|P�T�Iy���N���wpG�q6�z��	u�z��,�Dm���ʟ��=#{˿W��a*"pC��-��^B�W��ي#-�Zu��)�vj�OA"�治�X*>�J|����)���-�2����ĺ/��C�9m!Kۖ���? �����;e�8�0�!LD���i��k-���p~v^J��\��.�cM�1
}qb2��-Y��nbJC�cS�sqb�]��� z�
"§�`�6%����K���mq'�R��+UP�V�� �0�!L��o*!���V2BJ���Z@%�x�n-���>` B���G�e(L�#Fd �O�=7/[a��^�ꬿw�^��jp���0?d[��X%Ė���?�@3����u�+�?��q�<�Z�c�4�ِ�l��D��0��Y�y��xqqS��_�K��>�&�n��Z$����˗/���B����2.��Ğ�$A���"L����y����c��/�}�zsK�<��Xmksو�����=צ��n%�)[�/��/���F&����a"���������ĪJ��¨�2��rhuR�h(�k$��n&�!ez��9|ȠS���*.t���$ZJ,we4"��L��)cp�L�O?Ƙ�(I`0�l(����p�æ�ѣG�w]����U)5�4��gs!Gn��������_��S���8�b�ѽ���Z�M'e�� HH)�#�L�k�D���;3��V��[e눉:�%r[_T��r_\�7}��f�?�����r���b�Ou��Z�`�5؎�Ě���qK
b��O��	a:"pC��q�[zW�;�P��Z�ͣΏ����W�G&Y`�������z�WZ��0+d���Y�T<$f+wU@�p�x�|��<MJ�p�hHc��˅>|��_��׿�r���fF�]����d�i&�T��t��굂랑ݢx���M��!�p�!L�V26d�8��]b�-�<#�NCR���W�������/?�䓯�0+� Y1~Y1�D���)v�a2��X�̬�'dq��2���(�a�K]���@I	��Q g�6����l���#��|%�p;"pC�F�={VDL��5"��Q�֣l-�4*	j����I��kxY��dE��Ǹ}1ޞJ�
j2u��P!3K�է�����0���{��shl�M��}��R��j���d:w<ؼ�;���ݠz�0^6��̤7���aZ�*��9J��(�.Y`�s�U��M��&p|���HyBTg�����_��O9�\*�du�Q���=��U���dk��4�	X�k�K�;B9�V�X�3���ؒ�G�r�¿^�R\4��L�8"pC��q�*N
���ԧ��b;)&�	2~d�h:sq���}�Ls��㗪B�ʩ���M���l��(?A	��4�w68Ļ����7~Η�q�ܑ�[y�	1ц�f�z_m��I��ŞU��O�@�L�6���a"pC���������韾E�S���ryqCMG�x��Q���B�7��3D��tu�>�����_��OG�E��	�(ח�5�4�I�J�J����_2ݎ����%Ν����/ƿ���׻W5��⮱\��i6-�j
D㜢&4�v������O)JG��Č�v)q��G�&3�H�d��f?��F�>�]�p��P�=}Q����������?���(����`cC��[M�ͯ�q��iJZ�8'�/�g��?��?��7�|S3��x�̵I9�`C#��]�z�eJ���jwB8��&f(+	cR���`�#đ��m������ml��1��4�,��rX-W�VS�
;�L���c&K������o�zw��ǏK�ʃ�	��k��.���]�Q�7�u���Ű\,�wC�W��O~򓔢�p$�!L��5���*>	 -�Z �ZDǽ�auT�T=��q�����G�tf�㗣���ɓ'O�qr�� 3瓮J�v}UkuB�,�%r|$��3j0K#������ʵ̠]��ۈ�y|qq�^�K�Q��/���ϒ�BG���0�l\�⁫����d���s��)���x�:^���Y,��g~5�"|:�W�W_�˿�˗=:����ZN��y�|�x��^�y]j.q��s�u�����i^�9e|����������s�>�w�Q�W1�I�n�+(��F
A�R"6:ltqJa��گ�����D��0�bx�%4q\����R&3�qN�<��#D�P�-����;�3s�Jc&�#h:�ڜ(k��؈%�[��C��G�z�d��1&K	Q�G����JC��O9 (�dvU�2J��>w�@�r-S�@6W�Wy��~���D��0���q�z:
�/^�xQ�+�Z[�SѤ��=Y��ۯ�{5��n���秣P��2�4b�C��)7��T�q��e�)5�.�l��񻑬�3��J��N�	�o��vP)vndgqZL�s@Am6u��{ST�DD��0�:h�k��`[k�~����2��9�6�z�#�$�z���������td>�n���g��}����T1�Xj3#�#aZj.7C�(�z�\��%�$nW��4JH��K���o��oO�����g���]�����������%��8~����{���T�(�W�tB�H������oVB������H�B>�&]ќ�#L�f��^l�J�w��esɼ_"�7��Ͱ�����GF ud7k�t��8Q&O1W�u�L�&��Q?�y	X:�)?�D�n|>Y����܂����������\�^�L#,����'7�/��~,�ez��c���h�B���f�ŋkeg0s���������)�k,������I�:=��)�Mbj|n=��<|�p�c�ٽ��e	e�c���	�"`��D�2��၊�1��ju����/�x}�����~����������-q����k=5�fL2,�o^�{6�n'B���f`/+-xjD�X���Z�-x�R�G#
G����M�������v�ѣG�c���;�穄�6�ȎB�6aE}�S�ZE�w�^���;��&p�;�/��/���=y����Y�X������*��65�4%
�!�a""pC��qq��n��w�j�Lݕ"�("~�5�# �x\��ϝ��j���C�������j����~�;��g�3��L)�Z[�pL��X��|d�(K0�	�������k� i��/���g�����M�~��D��w@Hs��_6�x%����>�a"�}MS}k&    IEND�B`�PK
     w�O\�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     w�O\��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK
     w�O\acO��� �� /   images/90a26a0e-dc54-4725-bfe3-cfd4e64c35ea.png�PNG

   IHDR  �     ���Q   	pHYs       O%��  ��IDATx��i�^�y��;�g�g��HQ�dɲeɱ�Tn���P$�4h�E��Pn[$�Aq�~hj�E�k�h�[�7�se'��Y)��8�<<�|�;������h�EG�5�wA8����k|�3?��%I�K��K��K���Ox�\�7�N�8���j>����V+�$�lvuu�T*��g��]ڥ]ڥ]ڥ]��"��h4D��<???22���R�T�Oq �*��~��K��K��˝]2�"���Q�x����'��L��T�]ڥ]ڥ]���.�f3�ɢ���~�k���=�`&�l�٦���.��.��.wp�����$����������{��h��d2�\ޜ�T�]ڥ]ڥ]��.�lV��j�X�������_|����E����r�����m��.��.��.�rgQwH���O|�z��ʒ��;B/˺�6�o�vi�vi�v�����k%I���VWW[Icxx��K�����٦���.��.��.��.(yyyumyllljj���������G�A�Z)Km��.��.��.���)�Bam=���{��m4��w��ڲ~��K��K����������ŵZML�d�jm=����K��K��K�|p��~6��V�ٌ��_\\���iS�vi�vi�vi�N)�����|!��D��\.72<���E�6�o�vi�vi�v���b�(2���<;����W.���f�^�T*==}m��.��.��.��*��I���Wj�b��l6k��������.��.��.��+������W�^���.
���>y�o|�h4n���V�o�4~�/[��R0g�(���d0���N.�O��[�{Qn���3˻���6;~���*�;��M��7�dޡN�oӾ݆ow��->�Ռ�������{�?i��N/?b=�)�X/�ϕ3q�'�Ul�k+Ջ�����c��o$��g��l�z�!���AƗ��-�@�E��Y��_H�� �p�큔��r��[��?���O�~{��v��˝T��/�{�ܹ��v����~��'>�i�̅�����w"��n*�/,,�����l�R�׫ժ��1*�Z�������	����z>�'������F��g+h���R����	��Wq�9F�����H��4C�T+p!&򫸁f�i7���0[����)�e�mru��~�������I��_X!@C���ԙ3g���jkkk�j_�.��ED!�V.]�$Z><<�[��[���_���Se�M�bH����p�rs���,-��XZZZ^^�����e�%�C\�X
��n&�k.�-4�ij'�&�ɓ��x=�g�nJ�M��d����#_�N�Ӌ�j"�/�Ʀ�,#���56����;k˝Wn��j���*���Է]�埣@�D���^z���|e}��ѣ죒k����H����������ޡ����~��_�������؊�mK4I��h������G�5��������r�[�%_�8�ԑe��9�����ԋ�.dÖ��p2x5��5hj����V&q�旭כ�Z�aqq9�A�A�a�G)���F^�vD�!G������i
�-T�	}�5�<�s��3�{Đ�q۲J�Be�JQ����k�����ɂ���� ���$�0�x�~3���`z�tbt���v�O�|���7~0�Y�I[�;��_����_|��C�FFF���k׮E��~7߃C��D����ܜ�%O�>����uS�#�B�D��@��נ쎎��/�rY5՚�U�+�uH����J��0._�|����|�3�s>�R�hE)9M6�Z��(� �;F=��A��i}(����g��/��&`F㩠.�F�7����l�3gtt�Z�z�bFÃ�7��:Ư�4�jAð�PMl1���4�4p+;z����y���V#��>kӺ��i[-�*U8$c��*��;�f����7�ʭtZ��&^��7�#˿d}O��j�ۋ�.�2<<�w��m۶�<yrl�6шٙ������P}�!��!�p����{L�ľ}����)r����( �f���uuuU|р}�
j��M�|k�V�R���+W���?���sقZ����r��t����
�K�?.ݸ��	�U嵵�Q}�	>&������4���x�"�E��K��z���7dh�D���Zx���& �9N��X8�oJ�Y
�d����.����/�1^-��D�ƪb 6�i�A��4qM?0�4�g<P�4�4K7k�˭�����Mߧ-A�%7e6=�j6�W�{&��M`�$
��4Tڏ��o0�VMm�K�[M�o�x�y�s��;0d��Z�w_�M���_FGG�=*Y�ҥK:hG���sB�_D�Dn�8>��OF^�y�'&'':De��9ʍx�yA٪ T�_E���c�G+P��Cl=�8����"��f�;x�����E����� -3<�S��Aio%�j#��զ�3��[5����	Uf�ɛ"�aW��'�_��8C���
�����ދ��u��30�
��~�|񠴩�su�
|����(XO`��!v�_��(bgH���o;��ln%˚.�F�op�&Ϸ��y��G�ǆ@��5V�,)|~+��Z�ċ� �b�%F���Ӽ)\��|�V�S���kz�z�ȕ��EA�]�o�`�7�rn$��Z�[q��6n�%ܪܪ}����o�y�˿�"�!"��u�ԩ���kg�G	;f�u��������,�"���9���
�3�X
gԌd�����n>���?]L"Q���4�I/�^o�?�
m��!~�]�	$o��i�S��^�]�?����6�1�'���|Z�B�%i�M�`|��;���o�. 	�2󢾿L��(�b��#ˊ�c<===�W��/�v$�)�%\��P�AѲ1k�A-�+��W/����#DH��J]럪	�����ʶ�݉�z�Y�1;;��`��K���n���MD2`��`������;;�`�T_�Se� I`$�Q��-���a����R�S�#��13�.v��
x&>��44��R� ����a����As�fH���Q<�nG��I|�-J���.��p��kgG�� ¡f���o2�كu�W
̱V�a�lj�86��4Sȶ
D�Hg�!N�Z=6Z��jU�	��- �,5�2sd�wU8��u��%cC��Q8lV�:�E����e6��,���������bv@}ů�U+�)Wߨ]ܾ��>$o�y��OZ �� n�N��Q�T{l�(���3�H�{���T�7��o�w���6*=&)�0ht�Jq��	癚���c	ʣA��u�����Y0Ih>�s��6	LiYJ+�υq���e4B�3Z�\���R�"��{�?�|�C�z~�B��l51�Y ���`JhS������`k�Ԁ�54ۄ){X:[U��A�i�	H3Nik�@��M���dsT �GA
����el�P�
ĐX�,o��|�l�@�)#k�F���ig!	&	v�g9�	~�Y0x@`�- ��.cK��`l%Q��HV�\oE��P�u6wQ�5	nv�pٳ�&��6T�6��+v^ҌZ��f����V�	2�5zØUY"J�c�a�D���:8���'=a�Ҩ�<�9�,&T����gA�L���F�_�&^
�	��+�M��eK��m+@;��#c�@![��#?���"5��0I)���1Lr�=΄�4C���4h�Kd�ϴ�3-�eS�^�Xѿ���|�iZ�>~���w�_Y\|��}�Qq�#����R}�з�L	����k��}�
��MJ��=-7rq0���4yEn��3on� k}�a6��y����~�Lj���ȅ�5i'�ML�x��^��ȟh<]C\��@g����������%~`@�?3U�pB�����v��Z�Ф4��/i�0���Ԡ�5z� AF�v0ňA�:�\jB�T$�,"�wh�}�JL��$��&���v&�KF)_��6��Mz�����x��4�5ob�1�F3���`l�RZb���1
�&�$�� MVfYl�P�@ZPk�rY/i�L�7�������i�6��\/맩��+�� :�M<]�����[jt�!P�Ns�!�ubbB�B����r�σ��1�F�`�L!֯�(0vpb`�TPzS��.C���*�#�R���jV������{$,n� $g��/d5��g'm���;@�l�����B1�i�7���?Jz��r�����n�U]�YA�Ű�pӫqx��T��lp855%�������l�5�����$e<��2Ae�V�M�aB�'-���O|V��ˢ����Oeql��F9z��޽{��nIU?����������mQ}#����3)�-��0��W�r�@��$��80)��:����Ks �M�Be
��e��I��h�ť}�,b�g h��	vnp�55+ �H|����Yev~N�L�h��%}���HυSa�:�W�R�#��׎
��!;z�S��������4�po�x�6�>�����k�Sr�OscF�o�p��Lk
��W"3���P�<��)3�����lį�$��h���DS���81�D����C��fE!�3���0�	�F�.4��.fQ`AlA6��i�n���"�AI`�5v����F,�ܵ�&z ��2x�H�D���<�.k�_��E�zS&D(	&KցY��´N+<:�H���k��0F0�(�S��F��;����I���L	ci|b[`ۦ���>�4�^��l@K��ull_6��ҤZuPä�a��r�Z�}���K�x�C��y���.ol+M^m��!�
-�l�P�e�	π���%[)�}��X��`���hH��� �̙3��]'O���OzfffW�]|r۲~+h ᡌҟ�!}m�A�U�t�S�V����Tc����{-�}��A�թ���HX�"����T�T���^+��H��B�5��Pjq}����PG�ayyՇ����������*�{���jը��#|@�� DY<d�a��8*����o$?33v��� r� È2Q8�B���T����a&�Y��9�k&��Z��q�r�`6f�[�k�>��w�U�5��r!_Ѓ��3J���(�迖K��Q|�qG���'�[K��� 팲��L��7f��K���B���w�8�m���)z��s����F�x/3�F��4����-�c�&E���i���p~B}mMq�����'�.�'� 6��C�Q�4�^�$�^l��fc�����ezH�"G��*�yj�(�^/7I���y� rͤU�UQcf0�*I]Ma��k��L�θ:�\!��ޠ�Q���	�]�f�2��QR�tJ,U��#��9��B��Y�`mmS�6>!�S,��wjY {0+|��?�J��l��=-�{⦦����o�X0¦iE�$��_�����CX~��_ͫ�xn�����#�>����
�ST�)�Co�JE�{M�i6�Z�G��� j�[A���Y*V%M�M��K2��)
a ���� �4XSI#�i��*G)�$��E�K63Jya�<uq@5&�$��柛b�쀯�VZ�<i�VF�
�5��֘ɩ��-�]�W_}����B����0wF�YXKcJ�z�uY�7;�nB����;���z~	�F���;���6N#�~�7��Fh�gr3޸�*C}�v�}#%9cBU�D��v�h¡�M_3&t���(i�B���Bg���F�����qC��v
Q}���Ɂ� � �r�I�b S��3`�imz�4E1���L���̻;	�f+����>w7H��PG�Y)��!�h����f�!@M�������QAh�i�i��3R���^h0D`�Q�~t}vF���X(v�-N���/b���Dj3�eG��'���J&�6���N"���1oB�-o�n�V�|����j��gsF��`�Ң�'[YYA��穩)tW d�,�:}f�`�씆�O���d��]�f��`�R�]��Ck�3�9N����V�+B�B�d�W5F��D���zƗ�l4B��5�����A �bg{�{�W�1#b8�/���Y^-�yr�6�b�F��|3��Ѧ۠��ɀ��7�l1>
O5�d}��B���i��<�6I��J)t���6
ܿ�-Ie�0._%CG�`�I����=y��	B_3����	���\Q*�8H2�J\�"C5�[Ğ ��Ĥ�8F(�����ڔ#G�t��	]R�ۥ�iq���)=���I��T~$�`pio!�4�Ɇ��i��9$���x 
%|�%pp�����%d7R�lh>@%���G�.E)��`�C$!�P����M�)���W��ݛr�d��mI�ް�Fq��E:�$JC��\*WkU	�j%�h��'�Ф�
���Q���A}Et�w�2;�h[˜����rZ�l*n#`q�����0 �Y=wwuL&!Á��EA%�ɬiŬ=��Ʌ|(x�՚q-@����F3e,��5�ӛ�/:�@���Z���<�"�`�QꐚKZn��L։R͌a��q�V#�~� >�Q1�L�fG�͐:J�q��2�}-3�2��CY���<\�;ƿ�����*��by�����7(�՚��-[�\�z5�:(�W�u�]��=�@\3Aa�h%����&[ޚ�K��
j�X/��1_�+�������OS6f>�z�>$�qt�� ���2+�Y.�8�^���S9lJ����B��M���&$o{0���-����KC���8a0��k����0�Xe��N���Φ��}���&��U���Fq͂c��N�	!�F_Ө��6���u�t�>��,8z��	Mc��j�-��n�zS�f�G6�������1J�� dxx������G����ؕ_�:F�'��F7�Ϗ�L�V�E�^iA�ʞq��g��8�yWW���)�=�G�ӳ��Z�0'f��f�j+�j&e�MR.�QpB6�����n��s�\����ϫ&���;آ+i��d;P�gDp3lE�#�� JHҞ�ŭ�$��ȅC�]��hy�#B�Z)���c�f�@�& ����
�A� z�S&2��	��!�Y0�#ܛ}�j�^��-�U_h�F���7���"�t[�T���F��D�4B�7Ö	�q�Ol������d:0:��Of�`��E�ǆ8i"B�����}3e��>��/��`�U�b������A3L�f�Eg�ࡡ�fp�`�x6��}�_�FgƋ㍘��Z��ئc�B���t�),�FH�[�r�5N����Ȉ��^z�'����S���J$��r�-FN*�+�'z�/�(AL7U0��� y2�5���k��.Ax��s�v�n�R��*0��~,v���� ����a�#cN0�D���i�J�����! %R���CZ
���	u �6r�sX��z��S<%Y(S��������,�k�� `-��|F�Yj[r��Y\92�T����/i��;S�(8(�q���[!�¸�l&�451S����~��t�h�����)�f�]�h���YdB�&�����=t~�����OP�{HC"婚CӢ�y:�%�|���`I��Z��Nc^&�ӏ�euu�G9�!m�%(��fN�WV��7��_�r�V�V�����m3t�t}��G�s>9q�)=ѝ��8p� �ɉ�y@��8� �ଞ�+�u&�k�j�l������NON�M���8�t�0���h]��M��aiaQ��Z��י���ܴ֧��3�u�mt�!���5�q�X�g�i�����յeR���G�)�S���ag�UAc�x��E����Q$NW6��I�g���Ȫ����A����IK$���}�)A������*am�;;D�:�:�whd�`(7L�r (V���onv�1 (蓷�zk߾}&�$!?<͖�~�$r%H�8��F��(�}β3�? !���������(��˕�u�i��ϕ��{�ꍚҦOL^uTad��$'�厹�Y������|p?�![���"D�5��;vLNNj�ǎ���]��- ���я~��ŋX%�Oql1���	��F���d55���uyqIk2?;7<8���/�s�W��ǻ��<Wם�&H�!��O�������e�*M��j��JU�V�"qMԝ�ҥK:Z��n����x��R�8;=#�\��w���ejeԩ����|672沪�Fe�P�Z]e̍�����|������!�ӓs�w���*k�F-�Bd��B�����t� ����IRh�`;��!�Ö�&�* �˫+	���=t�Ъ/l�ɓ���33s�>�Q�UZ��9�W^yE8G�9�Ī�g|5���h�3� X�a����}Ҙ��r�#�:�a��^�xK/�)�<nٲe��T�àԝ����O��Je@��84qͷQo�4ְi��O>8yll,�+\D������:0�����3����Ҫԇ�\Q`Q*���������T�a&Δ������j�q�u��f�޺:��	�5�\	����e�O �ܿ�~�z���B��Y�Nf�(����sϡ�9��������3?�3�l>q�J�6���j߱��?Q��G��DF�'D��)o�����R�9����Kt}(jҟ��+�ަ�S6��"���L�<�@(Hi袣����$(�t	�yϞ=:�ݾ I3}�Q0�#�q�'�A�@=�c�7B�j5�������Wl�+xYf�#�1��A*��jA5I+�ʨ;aL��JLC�����5NMYDH5I �������t�H��E?m۶M킺�C�
hb��\�\�[����_���p%����A_��4�ɩIU�b�6RP��a�e�R�[n��F�]��C!�"~�W�Y��QC=j� �"@��߃�L���f� �v4�|�)�d	MF�;����+������۱�"�� � 4�D*0MP�Ԙ���e�ʺ\���'@p�^��d�z��Ǒz5AH>�3��� �A��kG�hEu��y`�#h�TS��˗9�8|i��@� �Ĩ4�*@9�
j����7��9ݵk�рxhq�N�vY5a����
�C��}��_=j%5k��&[�\<�����W㉄�`�:u*����Ύ�J�(L0�_�v6]cX�E��b�E�ew*��+�Aӧ ������▙3`Pԑ轸X"6Y%wZ�� �/��"`��q�ϟ�L5N���V$�>͛�6
z A?	P��!�F6�$!9���W�gන�	qi��9���9�����b�50��.T�މ�0����kvms�%�>,i�<6�=����y ��Y$?��m1������Z@���D;a�hdL�o�k�}�-W��ܗ�ih� �lH�aᑑGӹTD���)����H��S�X9:0
������\���8x$�)���`ZL1�͒�<-c����s���*_0_(�:Ŝ��Yƻ�����x�{�<Y�ZH~���Z�0����j �>%��)rj��J��/�9S�B<���Üy�VM���QAs']��߈s�'�P�V@k��hA.\� l_�g�^�>���b8Q-k�Nk�%6�X|L�X@�(s>]DBSP� DUNk��`rMh����LB{#d0�f3DW�b &��]�
�+��&]�����z�)Z(�.Bg��I*$-��� j8"-A�ZLA�F~��9@key�,o������	}��������'�
�5_!P�� '
��iUhq���۷O�/�$��c��'r��ѵ�'n����<*"�S���<p���D�7��λi�H���6i�@��7��r�ԔF��
UK�S���8W��z@[P�����^�^���T�Z�'N��Vb�<���Y
�2���x�^t]jV����;xƘ�x�1F>R)7��)=XF�bHEJ���_b.J���)�Q���g5H
y�q>�n�M{��-���p���G ҡ��C�jS�b���Th-��,�9X�4�J�3l#Ds<xP<���{��Ĥ>�)��=]4�o���Ju��M�`�`0�������T>�V���M�$��Q*s���$��dC&Z6���$�n@D�8���jB+�1���GH��ڏIX�>	���Y�����x#�a���?uu�@�؉��ʁrkT�;B�Dt�o�5Bs���b�^�+�!I��z@|'����G�>��C� D0,r?vkB��/^W�� � �x�Cxb������(�?>>��
M}�컐t�t��^w����
��U�H��5�-[��V���R�
� Lk�D�����l%vG�*�����������!p_��n��B�YO�`A�?�.T>��|��_�uRۂ�E/�љ3g���&�H�U�0�h;DTHP��S#��ARQS�]��^PY���%Vw�2�Lj��� �=�9�h��ף�<yR0F����V͔�=L�Z.�Ba�y�\ޗ�b��Ѣ�CA�5'B���h2>�E�B��Z�t�t:G_�	�C��A���D3�Z��!	�z������%��dJ�V˥%KG"p�>:<o��v�ܩ�jR8^0���ə��@�?ࠡye jJk���Zp �c���~�;$��}�c8W���
�� _m���9����h�sô�25�]��	:+��Dc�ه6L�ō݄�E�e��Y=�C�	� �$�����b4��;�V��۶�G�S�$jn"f��w��?�>�N3-��O�M?��΅̲&�o�$�����~���!�.� �[�7�1�n3����ޑ3t��5�����>4I%�A��yE���N�QC�Ex@���PZ�%� 
 ��:Ջ��`�W0X�g�#gX$y��]�s�BRt���GP��" ��D��`�й�/^�(R�f5Cd3�"�@)ʪ���Qբ�6���;�iF��)��F� W҅}��~�[Z��ϕ#LH#�!�h0����<@�����^��d=!��	D��<���d�����f8  =���l|��
d���6Y�|���e_���bI�T����E�QS	&a:UZ���C�v�BT�����_�R� TN˔L�f2��)��Ȟ�>�,8 ���Ҩ�!��'hHh��������W�g�G�c���{���q�����м��٣qj�G�QMq6p�� ���H��m��]F���t��l��_p�����ն��j͹4f�-�Z��L�-��Ϻ�E�GA���`�^���H/Ѭ@�5�
I�Te�����Kj%��1��tK��eǼjH}=�䡑�y��0��q�aa�}�;Pj�Vu�=`�ł%�����(�$�"	��ԥ~`:S���C�������(!#$�{�w�.!�yᘸ���D������ ��^�3>���cׯ��ެ�Nnۮ�O����
�������J�GA�������!����Ռ�ߴ�$��C�?�`���qOʅ�z��y>�R��C�!�Fejg�%�0��L���Sx&��y��a�֣`���(�DmC�����`}�s���N�s��d���jFE$��#T^��8������/.-���YA#9}����gj�0�R�Q�^�z&+̕6,5렿XГo۶��C�!����W��kA��GO��=��"�`*fA��0��(5bx�@E�^4O+��S��s�5l:[�-ؼ�r�J>����@H���4f�Q/p!�c-:s,����5�u`���4;�3l\����"q�<v��#�<��oDj,�R�jz�TG�bjV?�i��h����'~L���Է��Z	������+,_�4\�V5��ջ�S�蜀&Ry�E��W$?��]�&��Zp�{���
e�Ơ^��1�"kh���h���d P��j�$�b�!��H�Ԧ�V��3Ї�͔-��JfC�>
��X������ٳg�|��LH��ꔉ)G"�����2=5HM2~�����
@��v*	�x�hy]�8k�Μ9���V���?�V������| Ն�@ ��
-�Y��J0�0^�2�y���Ë���k��.
-U�3f��ß�!���aP��2î�C�,�L���VH�2�j��7	 �>B�#[b��;��v:K��\6�J̇������9��g��,ٛ�I�Ix���޹�4uOB"6{	�h�&�|m�t"B5B�F
�1ƫb? b�<=�0N\��%,Y�$��3�r ,����ό�̂v&�iEg[#��3�(�3�o�� y��|��F^ra'͆)'X�
Ӆ�4ͻ�Kg+Q���9PXnm�5�I'�L�F x�0b͹s�"կ0���r�!��
UX�Zئ5_2!��zB	�T�1D��F�`س��B �H����Y�s��5ȆVO�xD�o���1�G�9Ix@c:�?@_�'�5<(=��B�����Opi0yLJ���=R�5��6QC�}�P!����*ШDߠ:xZ`�������bT��ƥ�C����0}+�<�^&z�UM;���zB�1���5�(��aQ�|D{
�S4�8U�?���Xj�[ESsG�7�����
�&��w<K��(��V���]0��W����������}чCC�+���6W�[;�΂�jj9�"Z14�h����ͣ��aI��k�.�/��$�1}8���ʦ�`��������JGZ���$H�$!�@8U��9�����[�!����_'���)��f�����x��GeC����M^Pu4����l�v�� ��%|T�"o��yh�!���K/�Ō�����a��wi�1�;p�J�@o,����ߧ����gbd�c��[��M�6`41]�&��VE���D�:!�ѱ�AH�i����<���P�<(?�Uq�F����qp�F�&T���q�kc�	G���y�"2�VYc�s�v��'�$\�)���M7�
w-���ݻ3$�j�dY$�LuԵ�����p���B�	J��h�s��Tx���p��p����YF}(D'�m,�S_/.i��O3\�{�~�+	%��,J�[���L5�,l+j��u�vdC�y�7�_��1���~1r��!t������Z>��e̝�6�S5��	�ז�F��p��T�A0����_���d��ԋ�ꅫ�Y|�a\�>�>G߃��lB�R�ST|�[�҃�%E������z'�VHp�\���0��ǘ����ݻ���f�;���l�e�_Ոv�S@~��I<-P�aˇp�(�ҳ�<��oH�&6��G��x��^�U�jV�g;���A���$:_Qh9�x}���}>.����D�-�ǃr^���?��S��z�Q���B_IL�:�Բ�i$b�<PE�M�k���@�� <�9���g/
��u12���O���P9�!�L�%P��
]s�$h�p	�`"��M���J�a7m�z��D��`�ʙ����.���[!��Q��j6ܔ�����ѱ#G��y�TCZ�Y�R�DV�d�"0�u��Ly��X��MK|��MLG�EAΤR�G��A�2ק����N�"Y�g��iC 솞_`��1��z�_"O�kr1y�!r'~N�2�J��$d� ������r��
���j��K�C�0z����O�wӇΫAl�.���{�����D�*S����ƫM\]�U��ލ�j�s��ؾcj��JU ��&5�V VUa+�$(�F�PMB�^����UV/���??D���	��w�]k~��	Lш�q�R��bp~�ax��-K�P0F��4u��;������S#�p04��ىr��B����������"�.P9h��чd f��.ˆj+3!�!f~U�ڊB�C�(����p��9Ri^�X%���5r��(�����gQh�~r�������V�L_�N��A	��y�����}���8%Q�3!�.*�U/�!����Jj:hb�h0�wq��bO�,Fj��`�V�:>����P%�Q���ჵՀ5-J`b5��Hi���I�w��t�E~��6H=k=	$S��N�ډ�Я�Tl�^�!��u��*���Ϟ=+�A/E��eS}����0Z
��F�������
�	ډ�v�)�A͚����Y]�s�&�x�4C*��`f@�i"�h��V���
�A4�BJ����K�.�qf�`m�E��|���>|} ou�x�7oE�6Os�Ɔ�D/��O>���/k���(���)�5{���U�]�}yg� %�+��Fw�8u`+`�7[8�/����7~�^+��s��(�q!6A'
�c���7�*�wQH�L]Q��ꯄǻmxV_a �5�ޜ:s]:1�^\su�PBb�б�6���<�u����P���݇�}�Y�o�(�� t���S�Z�ܷo��VFd#H!�L8o뙻��R��ٽ��G#����n �ra.a
4�R�$b��xhy�R�x�8qqNa�O4�Jg[�E/�)�W���!v ���jk$lA����~i"0g07�Ν;5/�P�"%	��߄�g�t^xV@6s�T�dnny�nXq3$�!� z�LH�������kRD�A�$'> �-�aW_Yn�ϐ�
�U���"��c�1�����-�:`_'RNS��@+,Lz��)1�A���8v� �@Z2w	>����s�=�������U���x^�{ZO�9�e�dx\j7�+�SO=�uFD��fy��8-�_�Ns�XD���~q���{�%P�б�WQbA��Ks�7�d�6���
 Ԉ�QܭV ��.�P����j�C��za����;|��&�
jD�Ÿ�#m�F2����>�(�t��$�2<|5e��~�G�ja�r�|�:���]�7�~�P?~\o08�BQ���Ӄ��	�{��
��	� �\,���P^��ͳ�0�j06j��P>94��]�兂
�S����~��g����ؽX�A��E�D	7�L��Y��Ӗ$ujt���ꘟ���T-	��ӟ�u ! �3��ZH�S��ux���ML �3y�3��Eu6�H��f�"�7�Q���>���D���@^Ĕ@���:[�l��؋<�4c�d\�\�9�Uk���st��ׅ,���¼'�DoXi"M���A蛙���C"O0`��6Dx�O`�m!5~��y�����Z7MD���	@�c3F�G�s4�<
�FCX̄�u*£Ԥ���Oxl�� VJ��B�PG��S#�y����԰U_(�L55av²U�Ќ�ϙH|A6\pNGVF#�V�Hzx�f�����Ă S�3>�u+\��{�EZ,j�I.#u��z/�T����#G���A�p�U��W5%6I��@���z�:h5$�j��W��zHl
GL=��S�.�}TY�h~s���%L�9vq���פy-��KTS4���C�D����]��ꫯ���µp��w�P^�����&	���BsD�������O���E٣���`R���s���'6ˌ�84ZD�WM��M�������@����PÈ��`��ׂl������"�����\�B���i��#9��W�*ig_�u �L���ӟ�4*�!~�]U�����x��rA��vQn���UG��VVA)�!��*����eص(uQ�&:"����8���d���O�m�z�G�<
x��?C�q���h�M��=��~#\Og�VT �R�:��H�7/IF�/�����G���:�	��d�!
�n�x8[	��.b��@��Fe,���d܎��ZE�,��5�ʒ-�2jR�����]'AXպ�?bب7���Ԭj�L�Vl��D��;~4q�@x��v�a�'��?�h���>G#��!&"�i�§�	焲/0|��,�.PV���a�,19!+��VyM8q���7�{r!"�(7��Qd^+�K6.�Zl���^�اAԷ"~�FU�/VI4�xD�YXX=�8�a��z�"��p�ЮX7��:E�Z�Y�@�'80��� �B>��A⇴&��d������ȫ�Рh`b� �	ay�U�xv�؁�V$D���F��h	�{���b5T<�~�W/j�\q��L�R�����T����f`�4l��o�c5��Ϛ���lWZ<:Yp���k�WNv.�(�w2���{ｸ�E�I�� �P�FQ�Qi^Z
US��;���u���h
� �сa�j8��X>Q, �!.M TA�"#!7�b5�����"�.�qL�;2
h�4G�I�@�[59���S�jň �K�#�K!ô�f�5$��4I(����jh�)�H�o=�0�m.�o�	L�-�؏�V����=�7N�n������P�b��8��c�̟����f~t�QjO��D�7}b8����rQȞ�za����J$��GV��#A��:Yqi�\%>���N]�g�կP�\H[�Y�L�OB�<�]�(�|�V<��hAߪG�����A=���B[rlA;�,\�W���W�.(\&1�"�
�N����p��4©�G����H4/���r*��)��y�������ç�� v�C�Mɑꋑ �0��ƍ��@�_���	��x8ja�R+��#��p- �Z.�tU�rT�7yc���@L~Rx��r@�5<ځ�R�$�c��!�Z[��-����n`S5H)l�S��hJ᫘�eD(���	"a^��ߨֹ�Sʘ%j��4�B�y	̸;�/�V#�z/`8p��ިm"�n�'�U�Ȭ;�>���@B�q5@@G����>>[#<~��Ș~�tPbk��կ�rM�ԩSh��C�}��!�DT��;I1s>�z�jh��o�1�R9{挺�Ep�3>y�}����E��5�:���kջ�E��;x�1f��@/"�8v�6(�6tj>���Z]YɈ_��[n4�<ύcʪg84/qi�&ǆ��e�zL-���q{����6W�C���/��#�������\O]0�����E���p�	��� h�"�Yv�v�uFmS�b����3.'�DG r��P5���s��֛i����g�{z��R,�vy/�M#���o��or���3`3˙�?�6(8
����^��=:[�YT�F!�����U-�������V��8���	?�S�<� ����U��Eea�djXѢc�WM�ttO�>��s�����;vN\���ơ=n��#l�2�bD5�4¦D^�^�P�਌�."c&�L| ���^c��@�����8;�������!Unb�	��j�~T�>�s��(D=a�7F^j��D�>K.����>>�H03q�hz#/��-h�l�w%>1"x�Ų�[���a0�]�N!<�P��Dԑ2>Y�6W�T#xN�16��}L��MQ�5}%h����"��K2�bى&�r����[��0�����Q_��@��z_/���G��T��}�x��K-���qA�j���G
L�3g#��qQ,͔xwM\k���Q�UM�.�ہ���Ka�"?�0�nn^Ά���M�9RkZ+����B.�L����ṡ��S�Bkxj�N�>���:x8����s���?t��+���u01U����U_�Q#�\{-�NZ.�Eԣx)[�_�DW�
pNI0L,>�$��{����i�Ʀ�ش5�cn���qLpB� ��I�z�`k+��+���N�RG!uu��x�D�^"�B�T�so��='j�BI�7�WhO+dHL�q��r闹��69	�/`y�X0�--
�"���F+	Y�ҞE��M'
�#��|I��VBb����X�Q[������m8۝oIH4m1�8��J�N�ΐ9<���xarD�$��E��}:}͗D�9��WH	��������� �#��Z���	Rīe5���r��v$Ql��p�7�@�tu��BH;v}�"� \��F�a}?s�
O��H"����l����<ffMb�g\�!�x�U�=�9�/�^��O=c����x����a�@���OI�
̚@V��}�Qag͝tI�� tA ��&������2���y��'�0'�q
�K�Gգ]�O�6������n�;Z�jJ+�jJ����k�5Ќ�VU��Ĉ8�����>�|�p��.��Q�E3�s~���|*_�U��z�\yƚ�O�ʚ�v\À5�0��.Pѯ8vhx�������a'ĀC�h��8k�R����W_��{�!�/Fa��G	V��XxP<+a �>�&r�&��@���o�� O���k�3f�ٵ�z���)��eՄ��G��aL���>�1�����V��0�yX(R��9���f�°�0�Z�zj*�*w�Z�s*`�l�)Q��Vt3Y����T��^y�����G�Õ���f適;���U��6x׮������߈��(�����/�T�n2o;xj�
�%��K>��y�O�G�5�4����<W#�	��#1N�'�#�
�!��P{�j}"�G���o t�x~A!�c��O�/8�\.:<N7�m���4H}�,
�ۦ�P��˪jl����82Z�	w!fXю
a�0�� >w,��##��~=\��/����}G�1}	�pg�􌃍1_�������ٳ�)yA_e-"�Z��vr*x�����2yq��xz�#?��CT�LJ��pH��d|�bDU�������� e�h��P�C�h}��P���HWI��ЌD�Ը*k�Lۄ��[-��C!��^z	5F��R�L���E#-��
S=��SN�2���(� J�~��d�Gd�CS�!� �$vT5M����{ p���EQ�,�o��W�1A�V�C *�0���Wq(��I2;�?� @%8�K5?�`^��|�������֐�z�i"x"��@ �?t�ZV����&��.���P�_�)�5�fZ�]��Q��J���@n�:�5W8�p|�Y�J���<��ک�|�#ٌ;�8�a�gT�G����N�O`�U�Ad�0̱c�H�AL��f�M!/l���k�HX�ݻw��J-j<�Q:��(��*h\�yީ�R_������|�5�-#������,h�1�D�_���Oŉp9�)�e�N*�[��X�{�����/|Ap�����[+R�g�����O�K_��g��W��=O|ҢZC��3�o����M��ޏȐwcI�V�5��[!j/I._�$��6�������������<�r��{K��"�$-� )�ӰO|��B܊6ƿ�w!nm\7l�I�z��n����ߛ[k��נL7�c��b�,��Nr�.�۝$���R4�A���h.k�\� ���Z}���ֱ��fM��r�tW��ۨ�6*���~��o������JWow.��Q[_YlTr�|>v�8�5�b1�OP#�q]KR]_�z񷆚˫Ɨz���Lo�X�w]@�ţgh�	3ӓND�������wuwOM� �LR�
����+�,֊�n���j�Yo�����ޫ����[���ՑrIZ�N�UY/�sn�;˥|6�0?���e�~�\\XZ)ut՛ə7O됐 � ���aoP�������z����i'.�*�r��R�U��ܻ{�����E�?���	��`o������ݣ
3צ>��O
���*����v�;���t�f�;ʆ2q25�2�֛.��^^Yi4��g�QD�Y/^�9t���#�|����A++.G�:���'�p��g��`�{{��z��v�o�(��������С{�N͸���9G`�H�A�Ei����4:�|�\�kk���v-�,��#��ܽK#�W��,##.\�ܹ��{�0����z��5]��]=$����$IW�x��ٳNR_�X��Z��j��j�Z�W�;�7�y���.�'Qv{N�Ԭ��G�.���!�߆����M�gs���:��FS�I�טE����?��ӏ<��c�v�������'&4�%�u��j���%�z/���<{��ڋ��
+�sg�ܱm��lNu���b)�K�?x�c�F]ޞё�x�]�t������]n._Ҧt�6j��m���22&���ߧ�ӺI�������SOi�]���X�bQ�o�ܹ����3�sχ��9?�-���BQ.+v������ɕ���r��.�\���;�k�k�	�{Uu�{z9>��-��u$5#�d4TA2���C��!;�ŋ�15
4em�7�7|`yvV��[v��޽�%ˬ�-��p������S���^97�X�ɩAS_Y]���]Y]��*=�ʎ];4���.��7�x���^:�o��P�'��M����sq�1JE��jnΙ&&&GGǼ7����x�!~�sii�������7ӌ�kTp�$��ܽ!�v	�����&��-��_��X1rg�v�|�����]����慹��IH�~���7�����SޥiM����n��I��+�g��3���:ߟ�Β8�W_��W^?v�W~�Wz�F��lʜ�>���B�]����c괎�G$�����}��_}��>��Om�Jt:ޠ�"��\~#@��(i���L���7n�q�	��ú���W����k�|h>���Q�&ixz��{;M��pz �`�(��@ƅD��M�Vt�����vwu/-/�Sێ�K:�W.�5�������"�F�S�9m|ӥ���A�(~5;!�Je�b������Js.�T�!�����z�N��w����{.��\[����	�;�7��3
:������638�+�K���;}��������!=���]*���;Ӊ��r�6�u'4�?���Ǒ_qÌ�4I�eWG����Й(\ѧ@ׇ،�e-s�?���x� �/:vA
c3B�s��:�j6�ǚ���U[���6��f��@�e��	��ON_3��AWXI��+����\ń*D^^��g�P�e$fi:����p.۝��V�����y�1����(�1��-#��M���	Ӄ�&�'��0�T�u�.'�����g���hz�?8 E�؆���mDy	�em�� ǉ�qh)�-�hd�ûS�J�M������σ���0@� R� ��~t�P�_�}���,�hw�p��C����ߏ_�'9e�B����"�;�~�g��nJ���կ��T>N$��A����(wX�^r�.}.�`6���.�﬩��ǝ��A11<� �uA�����3�������Y�(!n�J->6l�t�p����_]Ћg�^�D�i��>16�p2>��V;88�\�Qk%&�~�&�ͨ;-�����N�|�&���[��5���7ϩ�C���y'�|�I�/!o�QD���K��O\�wwpF��K0 k0���P����yVm�w
�Y-\��9C���Q����Rt�����ƫvՈ�XXgaܶ���wK���W4?/���NB�@���\�I3���_���s��ۿw�C��3���VV���qg�����?&kІ�����yZCݵkG6�����S�������uזH|?t�Xȿ����������o����Qfǣ����s����۟�J'z�lN�#���AD��Z�X(�+�"�ͻ�a��|��Q�h��M�L)�}�),���p��{�1��Z�#����Z�V_h��y����qfiqQ����jgG���|V�f�F[q�Wzz��|RoT��{��^��o��Ξ�Pt�fǏ���7�v���?��?$�}�8А<�je1M�>?�@�H�/�8K|&�hZM���kw�ǥ�\X�H$���v�a��
I����R��|�#�/J�m�/N�4|�=q�5��.�-��={vjy���t�&�/f]�a�_�������n I��}��J��3��㸖Δ�e+K]Q����4>߼�2<<*񝤭$�jj5�>ש�N��92���I<qm��o���K]ݽj�������V�WJ�Z�:��|���[5-ײ��z�V(wj"�s�^�v���z�XP��JЍ��iǶ= k�����/
�FG�yXǄ+D�׫'N��ղ�g�[�뾅��9�a|ddH�����#^P;;4�]*�<wR\�ʲҋ�l������e��j��|�_454��֡��8@�bQ8�y��ѭ>���.YS.��+�E���ȣc[
�|�@/m�$��-����֯�>K�z9u�e�1���K��[ZD�A*ŗB�"�],Q�$��9 	���< d���[B��G�K��e�,|����j�޽/���E�8�W,�'*�"�K�\JZ��ͻĈ�Np��՟,Dӳ3�m۶�	ȕ���{]��E�5A�Ӈ�[��-䋵j��L��\�[�ӓr��suy��Ĥ����;fP5?��CZd�Ok����s[Ƿ/,.�y�R6S�eK�Smc�b஁���p4���jhݸ�����sW��� W"n\Ƒz������Ւ�$�G^s�R}eř�u��z�E�93=�&鿻W0��91��N�q޲ٜ����-+*0;=�[(&B��r�� ��U�MX%������x ��D
�DR]p�����f._	XW�<���>���7��������n�~ާ͆KP8���g�[et2�Z1n���������_��DG!��\*���Qf}���ژo~�"���(v��]�9�`i�?��믟x�'��#M8��C���m��i~3?@��z��b�}��r���/��裏��$�Q�::�Nf����ݵO�I�y��C������]5X����(�]dY��B>�h�k]z�;3!�|�Q��%�^�'Y��������[y#q�K/��]޷o����T��������w����?�����q6\ �U�r��9%)Y��9�q���������R�Ҷ���_$��u�[R�u��pZ��ލ�}'�3�D������O�>����g?;�u\,���J��q�����e}y9D$�KŊ����\	��S��UeQ�g�y�5�Zq�+�Un�fg��q�0�(���E;q�u=�Y��9�r��M�ؽ;rI�g�g���;�	A^7�	3b��4XO�\H��Ǐ����;/A�����f ����S'9U�^8��� Ҙ"��5��O]��e�!���N�+�:�?��	9�T3
��M�@^{'������%��Lr��R��Nb�=� ~10�,�9��on��_����8lD<Z:&���ǫHLy�<`�9�}$�d_K��[�� �����^D�"�q��dA�Jy]�@�������"�6����$�^#��t�2@p�-��IN�q� �CD���I!�M�ڄTc�UG��"=�q@O���e�E�9�~!�Q�X�i��׎z�!3njP��e���Y��}A�'���4�-բ�@ihh���9�To_��X���&HZJ��0}��%�݇��\��AB�A�G��=z�������p
����9n��u'�$��զ� ^x�C��l�i�z��C6Y�1l9�j�B��K�>�,��#}��wK�!Z.x�\�j.�MM���^r��\�����QY_�:.������o��o~�7�#�>����o�޻h�j�V�1_^[.w9E�k����o|C۰}縆�]q���#g������LwO���]S��y��ˏ<���]��X,G͚���ݓy����<	�뜀����������D�޺r��}w���� �� {��(iHDo��ت�j�T%���<z�������p���7#�b3�I��X�V�8�j�V�V:���K���U,�J�卫ӻ;�*����h&I�7��j�V#���� 7��N\]��)g
�+�ޕl�;��~��-#[4�G?���}��ǟ��O=��o������O8ňO�9�q;���죙���Rm�z����e3Y	�eI	��C#��_�2���+k�[��z�)��Ĺ��d��ZM+���L�����~�6=%y�����:����]��/I������>>g�o���?��?~�S������̓�Jeyhp���W�Zu#�Q[������	����ul��359����v��$Y�0��N��it�����r%cc�W�����GJY�iqi^���L����_�7��������  $T/9F�+[]].	�s���ɒ&�G/�M�e�>vw[��I &��+�{�].��Z��+�iB���f~�a�x?�008|��d���7:��� V�N���*���*��}Ou͹-I������	�Y&�S=�|`A�M,qDdah�}Z�~��
+�C���7Jf�\V�b�3 ����ʪ����#�ȁ=a���k6���G��t���?n�eu�����YBp�7�/��:4�J�$��֑���]T��ka��T��)[ rE��^:�Zs����a'��K˫ݽ}��F�8���%�&=ݝ�CI����V)�U�jjz6�/vyJ,�N|ʤ_�LNBkvu�G��R��WD�5��-�655������{::Z�fB.,��-�;}΃F}f���`�N���kמ5����%�:����gX��:���-�oE^dG Iɬ�t8}���E��y	wQLZĞ8��7O���NN�I������_	/N��XGgN�땲ˣ��̻k��P�tv:ˎ���b�}#.��mݶ1}qe���۩���{�H�8���W*k��1���h��h� �)�H˕U�Q�YS��eT(J1�z�	g��(!���m�0�E�K���d=�t��?���$��Zn�]���5/g`�]&�������_��_�����}�s=�H�^�й̺n]�M����i�{�����9s���}��Z�;vh��f�yᣁ׺Ξ��cǎ=��g$X��Ғ��K���_[_C����wG����.A�B�]r�RG&���`tx����_<?62N����3\h~>�Ƽ�&8�;v,�Ck���Y� ��/���]<[!����U���b^���`�^|�EI"H}Ζ_k�
�B��(��裏>���?��?������_޻g/VV�8�zM�Oޥq���ða��`�G��i�����x����S^����r�$#.(����Z����ν�+_������m�^��qwvv��_������s?�s�}�Rɵ`ɋЎ�:Kf7����Xt��@�NF[�S�$}:����0ک3:���)H�۱c�6Z�D�/����c[ƮMN������|�;o�5��o~����������wG�L�뺩f	+/g�\�.�4<8d�@�46���&&"�o�w<��J.06(�x�0W
�|�>.>��i:y�5��?��Ouw�|��_O�{������ٹ�-�Pԝ�u��\��d'fQpD�ឍe+��LC�INFE��*;>l٩:P��u���UR�:��e�隌Cgw	�ݍ,��9���^Y�%L��z#.�1z)��Ľa=U�"���O� �A�۪w��S�5�ύ8�v��B/��b��梁r)�/M��q;q҅��c�gzo.�i�K��Xr2붭��(i��>K{e^��(��� f�O�o@o��Y�2(��aY2=��`�w�ڔ���>���+4��rr0�7�
	|}@zZn�8{�,�K"t@�Nh�H����iz���Y�����'�?����KCxh
ˬ����Qrђ��z���˄�ƌB^ȍ�P��A��Xk
��]��g�\p�'�CR_��8U�D=j��&��\L�2����ݪ�F�������'^?
������+��r��uj����)^��v@H-���s��7��<�ړO}F��mD�S/�׆��M��{�g��y�#�=*���{�ߺ�)�3���ՙ��ٙ��Y���ۧ%訬�L�ҁ������<r�c����~�y��(۹����I���떴�x�Ux��,�ӓ��}��z�w����ow������ZXT��n$��`WOo�P|��g�9284�ig�$��J�=�x�V&���Jͱ�]�Rօ9�ν���LNN����$!�.���Q532�"���ٽk�_��_�w�}>� rq
I!W���{\�������C������$L��_��]���
��Q��/*��/WH<	�rn��fW��'˝�U���?���D���2�l������zkq���o��D�Kq⪣�߻�����������|gh�o��m�\fi�Z�TM�2����8�ʳ����/~�~Ip�*��z{;�������A�wS�p��>ȰTt�W_~�eb� \��a�[���f���{jfzyue��\o�����F���Ϳ���~ז��C3s����������g��ܽ���cPZ]�ΟC+P)8m������
�CH"�x6�.�S5԰���>�sj[���I���#6~��R�Y����L�������?���޿�8��/|������3����;kk��Ng��Z�:���	���]�=�՝�:�������k=՝$3��.`��n �Ey�B��}/��B�.���m�>���;:`�܍D�b����'����_����g?�ٮ����$y��Ԍ�ť�F���ץj�'˥e��h,ȩlV�N�C��ae�K�r>M�꤮:~��X@�M�#�X�l��������_�N�]{v9�����AՄW���q�s��sq+neK��-Cd��v�޽[#饗p@�N[b��*��1�l�U��l�!\W+u��*ww��RЩ�;��G�:M>��.N����U�e�b!��58::r횋�\Zr�/�=���Y1 ��ܬ�山�\OL�E0�fM>XCt̰_$��K}N~ƭ[��d�Z�kӼ��H��ɓ'�:�;w������$j���jaaQ��K$Z�ڹc�ŷ.���Ud��a��s�u�.]���Q���JfX-���}[�ʶm[��Y��]wݥ����M@ѳS3�\Q�����g1d�G�8F�w���٘n���j8o	�ǚ����LM_�kԖ��4mt���ԭ.{�������
bx��޻[�sE�ڳ������ߌm��'s�?g�'Y]��P�V�gzr�a3�dPQAD2�&��Xװʮ�ŕU�,H�Q`a�3L�9�t�x����Tݮ���[��z�WS]u�?����9�i�:)�u�B#���������XV����/)�^��2��'Gz���hӪ|,�M�3��%�ǵk$���>P�M�!$����]�X��a�V��X�zu�,�����\�h��Ol{C�I����eݦ|��.Xv�1����!�!�3�$�"��6�2)��7$]1���z�"��~���x���b��\�hAKs˪ի�y�7�?�|b�1fF�3��ü$?́б?w�q�C=t��_|�e�T&��H�F�qD��8��g�ɍ[�'����l�fEcS:�ǅ�t/��k�Y]ֶ7�k�{������x��R�qL����BITu�Z�yq�{�;��k�}�ܹu�A���+�m�9 ��̝$�)i3�Ύ6X$��J��̙3qnA`L�i�-�ѭ��W�zbz�V�1'���S&O�s�^w���1X��刪��)���%Z�n�u�]���}]���8&$�l��]���P�Aڠ��Qx�����b�*j�d�!Kp�Yo*�)F>mڔe˖A��k_{k�됦�4vV���?���ɯ���G�tz��G��0OTf�:�Qg��U)VI�3۱c�8#D&�.+� >�@)�� ���!ULz��K��^pƖ/�^|�ū���_���X�sf������A�8��'^O7�R�.Y��a)�]\�ƀ}*,*&pQ>q�9#N�PHL*�\x��u44<����9s$����.2�#�����/>b�Bi:�Sfy���4�6�B�+�� ٳo/h�j_��C��0)�YcD�a�!=�\X�oݺ��6Sy�d�3_F����������*���Gl��'�8ٖ\�_�oH�#�<k54$��D�H;XUv�Q���Av����0wz����.`���A#����<�������7n��/&M�r�J�~���m-8�0V�]Hw��ʌ�S��k���ޱ�V��=��Lk���'�%`G3L?��m��`M�ϟw�e�	>��~��� �X��cn)�\y��`�v^D	4cDv���_#LH-�ۻ���6i�����M��H��[��|�����K��$�G��2�I��tڙ6mҺu~{���>p��i�㘄�	��^�8	¡�N�C.M<$ ����Kv�O�b�<4X,j��ed�?��q�^�c����4ӡa�{dҁm�M��2�rq8o��g����˗?�f͛'�|��'HQ����*##�b�W�"��8��:�l��p���4�C`��Κ	�������[��G-���+��W��/�IR�����%�L=�f7o���c�w�y`a��Ē2"�\t\����V�JKX�r&�#�������1�Z�[K��s�?�wO�l�
�lт#6o��OW_��������؟�i��k_�*�`���Ga�O�ӧw�3㮛W�x���O?���,Y�~��%��ù���w_$HAc�qsS������� 1���p����+D0�6����s��޾e��uGF$*v�A�}����{|�[�M��^�+��q6Թ��7.s�I�#�Z���M��~�b��/Y�xqU;��R锔~���|n�q`	��>^����A�r)ƞ�hq[�	��t���{�k��okmt���.Ö�q��7��� ��(��+�aQ�H��m]�nMw���K/]���~y䑘葚
46�%SS�ȁ/�z��Fu��.d>�?����Ձ}L�����֭�'O��>������źz�̜6k�҅�����?z��'��E�g���ɦL#(��O�95���?�z��o����[��g�z!��`_qt�����9[�޷oO��Qh;	zJ��36d9��q�5V��_��PJI(�IX	���#P퟈�t���ң���<���k���j����P`Y��{W�^��W^1{�l�~*�̜:?�֯[��m,U��PJ�h�!a`ĥ!x>c�Ki`�����u�£cf([ޑ$*ɡ��	-{��--Y������}�j���'��u��׿����z�qǵ�Mٲm��`}]ƈ�M,:rA�\jl����0�@�֩1�03��<G�	��N8�"�X�D���ce �(p������gRN�>��-M��={r���9���>Ό�m��>t�]/�����}���ο����3�724�i���ij��ڹ��Cݐ�Z��E\
�؄`R*��*�!��nb3=@lyE����vJsz'��l?�[ji����J��%K�����������A��_��}𽣣Ro�s���=�w��0Q�9Q2��X-�W� a�G�B�t`�L���#�6}}�����1��LJe�/ց���������"SVY�OxH ������v"�T��\~4[��7�+���ؘ<�啬�d�]K}�a��"�if�H����E�T��^o�p�8ϗ_�9M8wj���O$\�6�?]��t �C��ݮ�������P�����]!�"B����.�o�U%�Hl��K�N��Z�k��]wݵf�fȃ֮J�W ��ccc�/qF�PmNn2-.��������Y�f?���6�n��lL"�R����S���ɋ�_�+��}�Y�ک��z��'�uv:�Y�r�jjn����
h��Gh<��X<#�{kkI�SA��\4�k\_���x��$)�S� �o�T�����`A(�A��Ě

~Cc����_y��s�=wƌ��Ӝ��bp(��N�:%v�V�a�$s��P�k"��b����Bjhȼ���?���XRfo�U�ۈ��z�S��R�0�=��U�V]y��\/��q+)����-
s/p-��b �������P�}0P�����)�:���T������:
t������~_�I��L&��V��C��)R�Z��|�+?�0,���3��� '����2�G��l��HL��
�>}	lD�h����΂~M��U4�	�,;�+��v�͏=����Qcl;�P�єV���g�y��_|�g�$Y�>�.`�z��BN�i����l1�G�@x���ꡑ03����&�������4��q��/~&�|Zn���|������?��al7֓�������;�;b�,sd�;���@_�GL�� 2�af �=]��Ʉ�V�h�����r��{9�3ϼ��I���ݘR�Y���K[7����?����n]}��i�p7��˾l����e�?����ف�y����0��%x $��iS�K|f�"F����}�5e�ąB�����x���[�Zq^0�{���g��򗿼�1���,ذI:P���k����Ͻ��VKωuMX_�F`�w�G]��z{r�$F2���P/�JԄ��n,f��{���'�SQ���T*�cۦ_���=�$�Ӱ��׬Z�d����W�!�bŊ��6i��������=�N���x��ݺy33s��$an?��Yj�?��:n������f<�H�(��yڏ�a�摉ыI}��ZH��J1�ڛGS�'/?L�c��.��\��D}]��Vd�[;��9ӧ�Z�n�4��3l�ƶM�X�nݶ���,���g׮+W�}饗�;bA}�8]ǭū+T��sn�Z�Y��zG;�-[֨^�Z��HBԕ�ۥR%�U.����O���f��y���}p�2t���O�7"���Dbߞ�~w�[K�}/�m���v®��#�Ѧ��!�L�#ã����L�F;Vb3�ǵ�7t�Z��mxf�AH�0>x=�7��K���HC�gv(�K%�U���1�u�K�����5C�7~�#�u��WN>��c�?Ű��Ш[����T��R�pL����dƱ]�ﺎy�gO�Q7Q4��o4�ԟ���1�[o��;��j��,�#^�u�(,�J
W�xRIW�̛��E-�"�5BK%wC��W���_V���Yg�}�9��)�k`B�����p�	�vKȦ��~��>RCC}���&���(Gc���{�=���dҙ}��]�����u��6nn�`}Ӑ�Q$2)
�seDQ�iSߑ�mk�+��'}�嗞;�����Ǡ�;�-�rVuk[�0����0���
�c�9b ���s�� M%����_O<��67n\����ǭ��:n\'��֖�x��U�0J$�J&�w���VG�H)zYtD��n���y�L��v*�'�nX�	^��0s�1f��80Z��Fs�CC���N$L�|�S���}����o�䉓�����_��HJ�m�hL�`�b<>V��n;4��dR��k�|���>���<=�g��H��v���?0R��4�#�L��`F؃$T�[�{��0g�]aHu����˔4	�7�Ϙ>UR�<�أ���7�+.������}�7V���\���nl|ϒ%���k~��o�����NJ��N6~{[k}]��o�X���,��>�4ہ0X�h��=�5n-���S�fA૯�:�|N���\Yy�{ߏѦ2�={{�����k�A��0Ѵا>%��r�����۳����3Ͼ��\���fΜ�{dU�(�߁ޞb~�r\�咏R� =�7m��$ %�ҝقX"pl�'F�#�p2)T
9�]*�~i���uԥ���N�0�0J�ѽ���{ｷ3۸p���ؽ1�N-[<�����o\�d鱟����3NCKrɲy��������GX�N���Ynʊ2:��IV9҇�s�*x�ʆX&�O8z�t���w�,i��߻��?>r߽w�3K��#R�,��r�W_zn���_�җ,:z|�I۷�y��7[�&��G�[��0a�%�?8ЗI'���*�F�)���Ϙq�K��
|���-*&f9��/B)����:����EӋ����gL��3��咤-���Ae�\fPm�+�W�
:V���ߝ�'e�j�N �Ū�%AUB&S.�N�*,D �6��80�	��s����`�wwO]���2����tzXbX��9�uP1���O��g��nnR�@mhb6���I�2lc5����Gř9r�8�n��a(�<˩�T�XH��+!���V���>{��ᡞ[n����_�ǘ�9:,�jC]���ۉ�0}�b�mW�ߏL[�z9�������|��^~���g�9IҊl���{U����bo4q(��ZA/x�W:�O8�����<�Я��wz��J�#6@�r����G��S��C���\H��ṏ=��}����O~:J*+�����9�`\���g�X��hg�𨠠ڂ��Ĵjii��Q*n��0n�s��l" ]hRc~^1T�Y�(�y���`�����n��k>���͝� ����HX�B�	�����, �BL[�����E�{w�ɧ��+W��í7?��3�b��#���Jո e���`b��C�8$c������Ւ�H��o�-�����AK3��;��3؏�%@��'���7�>ꨣ0BZؒƯ�Ӈ^�t�R�N<�����U�V9{�䈄���z��zl���n�L��8����_���'���g?;k�"̧�K��}=}�Z&+O�>�;�=���z�AklP��ca��}��)�5�W_q�+�|�3��Aܧݻ�
p7K�3����=��K.��[����O?��|���f͞��%?�!j1�ӉhI(=&���FK�d��|��Qh��˱�{�Eڭ&>����O�y��g��[a�747	���",��N��믿����O|�S�:��8z��o<�&iK��=}t�`�ؐ���� q+:����H���>:�Ԇ[t;C����G@*S�r����z�G��%,؜�L!d�3�p�w������]r�%نֆ�����u�W����,��G3U��.=�tj۽!4�m<ʳ'���3����O:�	�ܣT�^�쳏�[���J�Ɔ�]F��w��#�}�<u�k���r�WdJ��BYb�S�L�}:�;�-vQ"�uk�Sؾ};�q�q<1/6 HC��ˢ	ɂe/b��nM͌t��6F��iF����GJ�JҊٚ]#1c���V�{"E�Z;M�]H}�u���k��7i󦭖�̙=?����OQt��?�r����;���x�G�L˩��455����Y��P�&O��ž�����Ї>t�q�Վ��Es�+u�Q�Ͳ���i#�1�.��ľ	ai٦a�be��!& �a#�0�Mz���`|�[���m+7nxq��,X�Ȱ�,��ĠA�1�M��46&3Z�iKS�Ȃ���[n���e��Yh�\[Doo�ز�Q��$����VT-�-$tc��PhEd���{a�5ZmZx��o�㕟�Ї �>� ����>�Ң��ٴO��N'7n�$	5��>`���+_��7���[������ork�� R_�8FC,�dZ&A~)��y^Y���YN'I'R���ڤyd�T�� ٛ~��M��:��M�6�T�2���![*�I����_�Y�Rz��Med�����6}⤩3�{����w��bm�MiN$ڣ��y6���v[m��	�SZD�� ��ā�"H��+�1k�*��N�����6aB����0}����'L��w�(�t�2u�;�|JT���9�P�x��,-lF��ŋ��ٱ������?��O�j�Q�`�b�ԥ�%SkR��pr�d�&��ѽ�w���j$��ז���J�g��{��G��غj��O\z9�\=�Y��o&�^O�0~`�OOS8�k����а�F��Gs���߿o���]��v�����x�	�G=��AX`=��cيŒ��SY��L���vqUD�f�Le�:j��]�����}���Xö�� �����3�ԙ�
=��R�'D7��s��Kl2[5C�)�PKSLmh��7��ꪫ����}��O\p!�5#��uv�^���G����Aߚ4e���|�����o~���:�����/|��_m�� �a�3xzI����;��8�y��4l܌�C���� 8��ƘY��D�&-n���{�gx� jij�VOC�� ���(Mɤ���e�vw�7>�؃׭8�c�C���4eႹ;��/�VI�t8��cd�]�>�&6���=�Ab��'ba1~����`Y0Y��ʋccʤIK�-���ys������/
dE{=�ZC�����1�����d��~�~hi�Z���ԓ���K?�+�d��(� �Z��d��av݄j�~�Dn���v�i8M�?�<�M4�a�}��X�SOY���엥����ߍ��6�����'Fy�kkLgRv~��sS&��i�[ڳ�ܿ;��.���8����v���3X_�p:�H9	��n�&A�O50��P�XOL����8`g2�SZlh|��^�?Dݔ���fA=��z�QƖZ�sh�j����w�(hW��w��ԇḀ̄���@ӧ����������e���-��K��^^)�2�2�Z[M�$���Q.\�63A������Q�6�w�ڵg�}�"�����A&�m��k��5�T>�D_M+I�k,}k�duI�/���ʷv��=�y�{?֮0ץbё�{�����x�8c��?�s����-�_��~%�fc3�	�p��Z_��b�a�x���'
#�%���l����� �>�̋�:�,Sn�����g�5��L�PQ�\(��%0�����^x�9saxLO���1�F��4��pAѦaʅ�o�*-	��6��2:��ld�JWW�_��^\~�y���sSu�(Id�h�a�ɹ|��$@e�l����͍�=����=����:U�5��
�\MJ� �� ��T��x�5nYIAv����.&�c�h�����.��bC�����a���/������H��$pO�������k~�aQj'!�4�&�� ����L�a�|mMD;҄1Nr��~���?��_aO�,�2q�H�>	+� �	����	Ƣ���&ݳwH��庺�@��}����<���~P�q���۔��q�e��4?�)z�նP��˒\�pD��Qb=��]w�u�U?���삞�500��奭�K/���]�F`���Y8�vJeU7="����"����o}�[}����}�]�K���9����`�V;�Z�n��t��e�w�~��μ����_a%��g?���ӥ���Ǵ��xck;P��
J9s�2�����)晕�d���>�����?�p��#R�2o�TBc�DBl�������Q[����ٳ0�����8;�����{�$���n�h�g:�1ery�>m�S����	h(�#����"�-t���6o��_z�	o��ْ�^fh.�ԈFb>�����a/�緿����~�W�^oi��a������g����H`�cjķ&V?�,�b���F��[�`��Y���a��M�E��jp�����I)��������arRN��:�z��y䑯|�ʥK�vM��u˖��A|�Q��{�#�)~�bI=a.�m�kA8X�&Ҏ'03�6����ߔ/D�f�(� �tV��0�����&�Q^X���t��Uf������H����c�Ӧ���e�uS�d:oCk�V-]��
x"��agc��~�m��`54HI�h�hTk���3'�|2�����?�!2}k������5�s��$�]�2QC�c��A�T�)�mͤ���,f2iK�}}�	{ܸ�{�b':����{��{�������?�9+��� [ߪ��F���/�kj��sߣ�I�l�ŀi�	�HO�i�GF%3���]c�Kf�e3�\+�j�-�U�����!c�ޒ'�{AnhxhK�N�VsK������_�|��{/���e��:PQC�,��f��=�W2V�uAg�կ~��O���xĂ�?Z(��w���0��za��T\����&�� �V�a��J�6"�4��tx:�B�AB��,���oa'�&Nl߻w��_���Ͻ>�x�I�s��a���J&F�����=�Ʒq&�Lr׶u���c��XÄŐ�`�u����~��0�P�YfV���{c��~��ᑁt2�Ԑ-�r�o�2�m킭vï~��SO|���a�B(�VKs3Lp�y��`^l�v�D0y�7<���C���Y]�p6����ųӮS֥̍���/m�f�V/z�ف���l���>�K�nB�!�n��BR~�{�����+g͚ų�MՒ�S�����V�i��J�w,u����@M���}���w�قw@EC�}�r����f���W�_ΏA��d҅�VXXL���y"-!��Zf�&EөoHC�ɥ���`Ý����̝K����6��	+�(i��d͘B�҄0ٜ��
����/��;�c��_��p�q�/��ҖM�i�J�E����� &1�R6��͡�~����V���e���N8~��y����[o��;W^���?o�Bl�}�h4�0:�� �Ynٲ���f'c�/@��>آ׏~�#�����<u�>)Hez{�[Z�2��Xd�u����tJ��>��N�٘M&��X��M�yם�_ÍةI&ږu�W�X��õ�8��́����XR<���� X�&W�Ο?_zk���v�y���f	���zn���\��=F�Je�C=]`B+-����t�mn���34�o����?���؅�}�G���e��}���hC�g����q��&�Dt#V�1e���l��7����ķ��͙R,��ۻ#�ò.��}FEoh�k,��	3�lk�ݿ���qhXr�'tKF�W����?�_v���S�MۼiӶۋ���	��ش+���MS[�޶m�Apf�{�q""ch�1;�%�tn9ڰ�A.i'tBA�+�${=��D���hV�o"�F=�v�@O���I�S1�A��]���=�-��@��̛7�{
�h�#��i�M����0z�$�u�|��K^P��tM?�z��x�kх��v�z�)��m]K��\�*H@Pb#�PS�
JE�q?�ˢuBIĘم}q���^�Tr��ؾ����׭�bg�y��חW3��S��U��33uA+Rͥ��ȏ/V\�2�� f�3���&YsE�ǎ�B�G���ښ�[�tO�q��W���[����S2)�	�FV�~ �B�����'*�Q�و�6h��:I��2`�z�S6�W��xn�jO�%��&՝�.1�/~�w�%����:Q��$��r^B|H�tw���=��P/Ao�9q�Aw�ׁ9�XX~���3���5�o��tI}Y�Ȋm}&-{��t�"���j%X��%�\x�_������k�<�mƌ�quW�@x����	�$U e��D�����w�}��LH�n3Q�@O �"I��:x�n%G_��/��s�9���E�,�K�$#�ϴ��1BX���z*��j�W_}u� -dX�F����0��G,���F��Y�vS��@�YzNUq�}������D��8kV۫�����`g_p�e��eK�e��o��`���6l {��3s,��L�v�2BZO}p��p�m��Z/@n�a�Ղ�5�p��5k����/S�#�:l�]w������{��c�9��������)����/�����[�;Ɔ�a��yX�q�D�@ �1#X^�}�ʕ�mf%��t(����ڣ�I�x��_ed�TL�#�Ʋ��oRj�\}�џ��'���w!)Ǐ�<�ݹc7���Y�h�1�O���t�0�aC	H7e����
��-����C�� C�+ɳKh��mI࠾��`�G�I�L�#�3�c=�r�W�~��8A�\�&x������yy��71M�$�d���|���#0x"���Pm�����~��/��҄�r����52��/ma���p؝A*-M9M�M�J��,���Ԁ2A�����`��和g|'֧dGl��<D�l�W��Ŷ�==��C��+�n��D��^R� �3X�+�q�p�sM�㆔z�,�ć�J��ͬ������5(��U�h�s�O2��UJ7uVgg�qǽ��� �<�斖�۷(���J��.���C/[��^�Fޓ���}����S�[����l��ڜM9V9u�@N���/t_*B�?x�U�w�M1E!T�����s�� ��\��2��n*����zA(�$2D�&|��J^m-h$M�L�-���6�O�`O{��y�
7U�/��g��z�J�����]�����{��Z��@L�v6N+����In]9��(x`%�x�ꎮ�G߇F �ӕ4� a^���\���k[��l*��^_��3!��>���>=c�Q��+��b��#}`sO>yK6S��H��#�C���d)W	��B݇ґ�.���آx�6>���L��Ǚ!3�9L���cd`s�u�;[����ww������*G�CK��@l�wo�9s�=kO=mI[cZbifq�]�1/���"2���T(��i���D��s8*,����x�Q���L�~� �F��(@�,1�Bި���Z�n�����o��<��L�.y�t658$��Ҡ�J�^��>��];V}����#��͞2�<�fP}rCP~n����+��r���o^Т�n:�� T�\+U�9,��%]r�x�di��Q�D�ï�w��{��/���g�s�tjͺy蚶;mڬD"e%��e�{�o[����Һ}�������k�C�v�@��a��A#*���꣋�S1T�+�9J�D/�B�= T4=�[�HCד��R�����Η������~�#9��Nb��K7n�:���ԥ���ړ�aJ/��;�ADuO����__|�W?�x��g���C���ݏ��۽g��#
�<� ^�<��+M��982�+�д{����7BE�5c6$Ё��##�7o_�d�g�u�Y����!�������w.���F"��)S:�L�a��;�C	�{Ĝ^x���FnY�A
R=���EE����|��_���?y䑗|��$�����{b�Y���W��v��.�ʤ�;e+�64��9�H�1���U��DdDE�6�u$ۚZ��7���8d�e�~�>�:�����޽aw/xrρ�%*c��h N�����	F�vI���\\4o�ԩ����x���T��tkGk� u߰}�*]�0��%s�D���h�9'��I��I�H�OD�˻П�����)-����[��;���.��h���iݖm�C���5�02*&/�τq3@ �LvhD�|�eo��]�����~ʤ�-m"z�y�wO<�̚9!!	Y��^��,#ȍD�Fh������Iߐ&2�|o�\*�Su��c����S7��sw}�c��ߝļ�����N���̤;�o���ֱ�������iS�s{�ZR#C���RN�j�'�r���%>���֫K>)T�R��L��XJ۫z���,pۤ�ӔI�Ki������.H�u���Qf��Us�ƇQb(כ��*;l�u�7
�۱<���ffW�Ȥ�l_�Ю]{�O�Y����Ye��+f��4]����G��Ȩ���&pƚ��*������Pc/��	�(><PaTՖ��ÿuY�7�B�Łs��<�8�?���aX-��7��M�+�1lM�g�]ҫ�z�	
�$�������5^}���ï���i|!���᫋#9�Y���2�̍�I-�Dֲ��2�hl<��X�STB�VSB���_D��dT��S�Έ]a��'Y0�J'2B�rI�6=����5��<�񂥴 T���¨�O\������J��w$�W.E�����\��/`F7���sKu��K/��o�|�g}Ƣ3L�Z�c*�!A��}�����P�ER�j�W�_����ş������f����Z=��3qݿ������������>�'����bʌո��2�����M;�ٸv&���uAL<R�j$)[2��
��2�tXRH�M��a$�gN�9s��5�Y�����̀�~��כ�Z�?^Zx�޳��o���?z�D��C�Ua�X���R���e	��Jی��+ �E�{챟��g`ֳ�2����7�xc˖-������?���������O~�[~�����3��L��I�ڳWz/e�%�fT�>���}�;��;���?_��kN<�į~��<�I7ɞ7􉲨��W�ƚh-nGuǂ��s��x�{��|���ӽ|��<�����:��k� �n���ٙmlRρ`��B���X9ꨣ:����_y���{뭷|?�yj��xLZzHyc���q�Bs�k�c-��t��}�Ż���W_x��N� ��f��w &u�=�ć�(b���ƪ�{�^!�늅�[o�
޹C�흒-dh���'��J���`�n}��7e����	'��sGϭ�޺��7/��ҩ�-�0a�
�X.�,[�ڪI����+�}�^ܡ���YDaN(�.�Ȝ����y/�����Θ��@�N��Y�B�1�X$r��8Z&���<Www;�*f�ƻ��UIL`��'b�#a$�T�̀![Z[[ۊ�Rnh��U�U�V���
��Tr�d�ˏ	���وi*�|��8�~��h��8?_9�X�{ۨ]��B����O�x��\4�	J.��־g��U�zB��-I���$�_��Q�ٴ/.	�CJJ&��:������?R.j2��%8k���uSGH�>VKVƯ��z��:�[��fꁡʓM�jɪǣ��JjcTP\_��T�F�~E��;ǲ>�5D��$'N��!�����g�ǽ��xe�SRuS�9�����i�т�H�x��$�$,�@�SAi�x?|�_�����"��]{vw��;:@�{��<T��{Ȗ�X����!W;� �-ޝT:҈�t���h۽s�h޼y�U��2<�K׮]�ꫯby'M��oPu0�I��-)��E�U@]gљ�0xnKK�А٧h�_�������mμ��VU>�׳o����m۶�}�BH��Ifx��W�����;��U�k�k�P����,ޭ���$�
IG�h��|2����?��O�:z�W��v�w�&�3��5kf̘q�q�ٵk�_y�������O��??�cc�IO�4�K)#����69�����O�7o�L�>�lf�3םYl��0_~��3�:��[���g���7�x�g?��{ߛ8ej2��%�m�]��u뤈�a2�?0t�{O��o���������O���p���b��G(� ��������u�����(�Q饶j׈hH��獌��5�׾~Ú�.>���_��o|�m���	]##ð8!&�*��l�Z��kV���?�K��hߎk��4�}�vcA&Lj�J#	h�=����"SS�!#a1���OME�ƈg0��Yܱ{{]cױ�O߼}���߳�}���'��O費�&��ZO����Y.'/9rp�vm}]R�����9�:���k�+؝�W`�M\g��/q%C|�x�:�!��B��0Ҭk$lõ"R�L�R�#>�j�T-�B8:42q��93�mذ��������v���?�y����om0��=;�L�:u\W}o����>�W����f��P[k�a"'#AQn���1�${H�A;�h%Eo����ο�ޢ�'+�ȝw(g�u/���d�GD-=�	;���%餩�Y���U���D¢8!�;f2펍�Y�ļ�(�ă���E3I�a�yƌ)�kƐ*W��r�U�7��؏Wq-l�3��d��m'�H¢���t� mcRa(��S�JN��e�$��Ջ�?��0������|�U[�p����T9g��$-x�	�}^��|l�a�qZd^:��P��޷ՙ������zJ�CQ�c�<Dߏ����V���j��=|���g����E�
��آ/DR��ţ��3�Ѫt5ռ*�(G�����

y*^����%F�M���qb![���Ch��4T�+\�b>�!�����<��^����wp�D��5^�.�"�aH���\҄}챧���s��]b�G���vh��uG9/���fɤ$ۏ�G���~����ᣭ��!>��`�Ǌ��
��:93�z�qRu9MR~�a��i�'i�ۀ��밃�5E�ԧ>��k�=48x�M7��k���ŋK=tcȻc�lA���,���;E��@{a`q0r��.	�ϦL<z���z꩓N=�g���c�}�'~~��`�WA�J��������+�L�:眏nܸ���ǎ�z�`���,Q� �ɉ��)�~E�'�=Z�m�a��#�m��}���^��X~P�eJ�	T(P����O<��/}�[�~6w��{�����f�Wi1aؽw�v�=�����~���ØQ҉�^�\T)�Ȯ��Q�Ċ�UN���֘(���H ����� hl_��N~�����q��K��\�aŊ��~.VlѢE���}{������=��þ_��Mܭ�E��C_R2���LQ�x'>/�j+Q�6���g?��J�mt�*N�2e׮]�����u�_r'�be��҉ѱ�����zl^����$�!��P����]��֞x�B(JxNN�؍5;��ز��"�D1�Luֵ�1���q��a<�<�n��kZ	�w-��* 0��:��)rA�	���e��L���ƶ��t�.!�^����!%�FY���0*�ʣ�mr���m��:�HYSP)&�'�^9c˴(��qʪ��;sè,�^a�/��A�F0jE����i��+�LY������!��4�h(ٞ�xFB2�C��$Upe�M�#�-�u@Ў"P��֥��Iɢ�L�"��@=���Y��ID��JU�*�9���L9#�Vy/i�j�?��p�� �)����V��ه�eFb��Ac5Ht#���y�i Q��+'��\�"�b����c����ﳩQ�[e��:�qb]��`
%����6�3�P�WK�׉$�X�	���݆`w	t���|�M�D�Vh�X�#���_ǥhV���!+�yZ��R�],���=?(@b��u\��V�Lx��)�3�i�F���#vM[뿥��p�Y����rl�/{�G]�$|����J��NWʅ�-Mnc}�/K���Õ�3����B�m�FR;]Øl|���k����#�q�.vy�_ʜ2uݪ�:��X�;}�d0ʞ��g��ئ?��O>����Sǉ���BZ��i���=p��۷S��V{�Z
��`��^x��t06y�ߋ�.|��s}�!�x��7�X�t���;���O<��n������\�M�0i�n��۲i�CϞ}�=���+WCw9��x����!�$��i���0��M��nB`��G{HB��l0��D,ZH��Pa:��C�*S���_�
F��m	N�ڒ��O������7�,�?{�=��SŚ쑜�%G͛1}�7��馛֭Y�'��Ϊ ��r��JM�F&m�R��]P�/�%��[6|iIV��f�Sv��T��  �S�>Z�r�dI�F�I�wn~�����?x�N?���~��ɝ]���ׯ݀�4ֹӎ[�P<����׼(��n��F�t0p���>
|H�TM�W홂�ϻ�����x_\V`Ts�+_�	a�b�y��
�裻�|㶧���K_��G1h���M�mt,;�v��K�J2?�6X�T�;κu�� "�c������� �5aN7��S �ȬFy�hZ�O|'���U���I����ܗ0*����-Z�_�Z�CVc�F5@b4�C;�n.2,(t�f���S%L�FS�6~�-�5�<e/��$=��eKsZ?�A�ry'��VU��
Ĥ=�_�6��2,���z��6x�Vy:������ahd�J�\�F�J��'k�� a������,#f��f�Q�]����
��q��E�㋛��}�P3�C�X���A�ÏR��
1�2r����k뺪�k	�c
yy~e����0E�ꘇ��ZO@��QM* �<��t��ylE]�p�����F�֗^���`"���T�+zI���aT(AQԚ!���ŘY\�S��c��턔Q���4��@]���*�+��Oh�9`>��
�s���30���j��8�!��U�QV�z�(���c��0��ZX)�t(��/C&1�L�X�Κn"���;i3c�1��5��Y�<	�*���ǳ�:����zB���p��3+�}z�����D�o
G*M�N9�M���&f̝f�:N1�ET8�eb�*��ฏ�k�f��͛7�	���g.��҇~���>҉'a�V��1c��S*>��ի�[@5��S2g3�
�v���=��TV��/q}KϬ��{tcB�a����t/��S�:�N��Y�ئ����g�{.�eX�O|���]-]'v��9{&xո������)���EKs��Ha�	�H(��"�
�Q+�+U3&9�=@��@��Jq���ӳ�u�p�w`v<�l3/��ɔư�X��nڶm[C6����TTI34�MI
aR�A32�~XHNqbVUR�(Ծ2R��֖6v��d3i��X� .Z����?��.��렇�6���'m�+� ���g+A/��hH�@���mx�l˄�AI�"y䑯��
 �a��`�o�p!(�B�%���]��;��V|O�#E�=C�����hT�k�+G�+��ءo�,EQ����<y�)�0�l�qXm}P�$��pf��c��q��*��M"l�r�۞i����m;��F3J�Uu6�W���ͦo�T�e���x ��h�i�O9=SR���.��UL툢ߐ;'m���Y����
�e�)[��]�*a^�Ή���h�O�Ү�1O���K���oX��G����}�%��XV��>h����ٚ����Z�[��� [[[��1%���ȧ/��a��y�s3��U��u.��<�Z�O�W�~u����}����ﶴ���1�!�r�vg�K�b*+\ҍ
���%�ͮ����~�T,�^*��k�O��U�_iB�t�ث�*���Ъ�K��j�Ռ$�I��ơ�;����HH����T�c�u"��b�Ό��f2�b��Ql�򛱛��-T�;ǰh��[,�z�6�M����R_Y�z{�8�.�uu�����%��IKá���+�������?.�UD���)?0{��b��r(er���'�0���zA��`{Cvٹ[��ry��@BO�4�&l>���	�L�m�&�K�,!J� x���E�D�}饗���y��;�����<����3uن�3goڸ�{���.���Ji��{�̲d4����p�>�K{���8�`��m�Ј�A[_S\���D@DI�4�Gj���T�Z�����������h���{o�عmcy���i��̎�}ÃC��A-��^��n۲��mk�����8 rWzv�>�l�a6փ��LM���@{fJڋmz��	�Vż�^,YMs��y~�N ���̼1�����ݖۺx~W}�������>�}�}���--��Ҩf�������m�O��� Ml��3.�q�u�`�Mu��Lc_|�k=�|:?���	�<��ڎk���7��DZB����PUgME]p��>�:����<�"�$R�����:�!�����p֊%��R��ע6�k*��d�ipl
H5������з_Ћ�w������X�1� '.��8��p���L3
Z[��O���������/��*R����4�Y�g&N2�n�a�t P3�p��Mq{W��v�5��U-�J}Ͷ�H}e~�Nk�(	ic��N Ԝ�EG�f�&�W�(�e�h��28m8��h����;����d�hą�xG�Cu��d��&5��/]�d���F�M� 'N|YaŖ���}��li	�co�p��O��Rh�.�"U�QE��QJ�bP�W��QTs���^��I��z�(\U�C��@��ӺPNY,�n5ɹ��{�ޮ�TAN��-��Uv�H�P+����I���cWU��j����ѷ?��ٮ��K�$�;Htv�Ь'!�S��&������t��x���PZ����&2R��]��oe��&�+N�=PIx��U���1p;�X5n��>��-��RK�|��r�tƴS�M��Y�����I�k��$X��ݒI.�px�w�-6��gҤI�o�T\�v-+2������3�ipÔ&K��CK�]��$qjYuͮ�0�Yψ �:E{nں����vۦ�[O;�T*-:�)�DS:�u����`7��I�2,Kf\gۖ-[$d�\�P>)&~���-<��� ��UzP}�����&fȣQd�慥*-^�$��	g�
�dU߆�-f-��ubb��{I��DU	��L�7k��Ư9��6&�	G�]�B�B���P��n.�����[��Z� uq���O&hx�s�ۋv'Qd@�I�_FU��9�Q#�����V�ӿbi{�J^EBm>'�L��!��G�l�k:I:l�J%�"�a�=I��S�A<��f=Q@��rc���w��'LC�3[
.�qC�9Y:BU��~�wA W�����׽�꫹��ӦM�=1>�r,���E��|�I��%^�($is����?�{��5$�Ne��Zz�tZ�)>�ku��{���67->j~6����Lc^~Ų�:&M?JI�4�*.6:ứL2ረ-)ty�ipƢ�`�6�����K��p��&ltЯk�b�¸g�w\�U5�Mʤ(�X*&��핃�#%)7	U��ܨ��ީ{�J�� ���:H����L��tSq<&V8�-�g�egTa�6
T��+�jړ�;��x+E�D�:el�"��,3tb����o#ѹ�x�Q +���V:g-���:�ڊ'��s�s�Ʀ�����Z��1�^�/�ҞQQ�,w r���r��:*m���K�Y�.�~�����=��_m����<f:Ƙ���HDEz|N9�;9b���U��B�2Æ�zL�T.�w�����QF%'-�J�pF�rE�L���|�onmK*��T�?��;ɸ��!�-�U�aݼ��9�����_��"_O��߷g��Y"��RcHE��k���~iE��rӬ��ͣ��Ԩ)��>K�ڴ~ �����~ScK�P6$��h57	����F�3�hGݲ�;Q��c
� �]a�ԩ����Lʖ��8�@�>ƾ/�M��w�͛�ϰ1�)��+�C!��`O/FeB���DiH&7nܸm����_�)�&�1454��d���/9����pgH�y���T�A_��Qq�z�k���h��#ڬV�1��W@��,��~`�h6	�R���Rپ�^���*�ӆ�4Г������������z�%j�فԂD�k��0���aK��k��h4�7��paT�(U_��$�vb�(K�L��1�	� ���������v��\���Ha���=���9��F�{2�!x0�ăr���ԲB�(Xf�x'�_����������~������֤��RyȌ�)7m��,4���� زu;ȩ�>	rʍ�=�B��DHbE�A�4I�7P�����wJ�N�ȖH��JT*+��^&��`�S� v�d�[���v!2|0���v�^��������ɓ'ےu����S���tӪ��g�\CI�7b��%f�Qu��v�81?�W�.�sBҙ5�V5��R�V+�2�m��l}̢2k�f-����
��S��ʩ��.D��X�	S�=�b�EDT��ҝ��>���;�ݛV%V=��n�8�o� yq#U�[�I���E뢝Jgi%�^:$ENeGD��19D���M"��cR��S|�����j+`�T�P�Fs�]�����_�#ҚJb����H)�d��5�/�B�`5#�jTs���ɔ��?L�W�.�De��\��ڒs�g6hDRd�Ve	&����U�7k����4�z���<��}���p��wFscX�4p �KL�_������[�̔�����K䓨�;����W����ԑzɔ��%5�ΰ�q<�u\=S[M:N�v��s������m�FԳѡa��S\o��6m��=~|ww7Q�i�*h���n,&�1D��Zw�s�Λ�:~e6�oP&�N�����������	;�L���v	�ڗ�#Ӵ;��>馡%��l�`�gɃ���$���9�K"Ι9�*اU�E�	�� �.���ş�=�︉�b��r]ș���~�.j����aVk�7�1e��j팡6.�4�R���o}����H�h�9K�C�cމ�ז�T섘��Y�}ĭ؎�L^ZZ�˝�)P#��G}61�r@o?s���ڣˮ�ᱪe,%�ԜR\�Ϛ,b�s6����#�;�`żo��c��w�ï��%h䂢Œ� ��ƴ������1,fW��N��vvb��18h��ql�Q��z��V�P�hC<|��}O�Lp!:�M�"�JSd�I`젩����+�ǲ�Z�Y�l��S����ܒj��+q�H��|Dw6T'1��Qae��%X�nm���V2a����b2P���Q�
�aV3���eVUf����%��(&G�ʏ��3ǻ��Zdz&��y��i̻B@�{9��n�Q�J>N(�1Y,�x��Rl�#��f5�[��m�"��gP�����чv�X,���o9n)�Pk���6M�u��´l֔�����<Z�!E�V����iN<:��w��BƉx�}�~ �z�t�VD�'�w����I$݄��Swhj`Kl���m���ұԯ���dϨ�!�����p��?��#��5�80��/% D�oen2��!���Ե6	~�+�T&���fE�,�����w�ߪ$,x��Q%H����EJ�%&�<�Ȕ�������&�1}��(�\ϨT�Ⱦ���xb��T$���v�bt�^}0\AX��U�z�H>ƺf�o͚50TbL'|�r`hP�r�YP'F%�l!'?����
�*ڕ�JX�憒W�
0�����H�TKdEՀ�1�7��+�ʎ�a��^.7�ђB����u�x7��)�$GCuScL���G 2Tr$v3���\,��4��g�3�8e*+�R�[�d�z�H��8�le�����<_�0��>VE�i�gE���+U�U�����8��t��,�I�C�[�tE��0�G�d���)ؔ7�I7�t5c@Y�%���������|�*Q-�ј�d�<A���[T?@<�����)�+e�%�kuL6(�e�{����2$�.(�0W	/��L%7(��]�r�Y�˰@^S�����4�,��#�0|)��kh; )r�f�K��b���= �_�
,�X{�3%@(������SN�H߁ ͣZ%����Q�Z���*3U$��G1.H0�լ&�/�`�EՎ?�Ǩ�Sg6����x�T�J�Q�0���'��8z�`��bU�<Uq�Pi��<�����1B<�5�hU�\�w���V�w��m�.�+��Qu�d�tx\^Έ5�$Fȍ��G��6I���Dƭ�R���^X��;�/����e�O�Š�AA�q��SYs�pj�/�\l@�҃.��M�C�ե������R)�ؖq(�B�1e�r�>�X¦����S�+ ��eU>*i�zg0\1�m��P�Ī���N�4k�f-�9֡�Z�4S�DJ��U$*�}�)���ū�c�>�(����s�{�R?��աR�d�ԋ��L��t�8��8
�%��0Ggm&��b���J��e��*@�R��k����[��� ��=9p��eO�'�M�6�ߏ�uk�Zo��t6/�q6}�t��\��Ia!��4��y_��L�� -{��(#�%=Mx4T��S&��x���j�H��hPm'FXm͕�j���5�jI��\�^T�L���������ɯpyөt�����rX8S��d�Ud@��M�ZBZ	���f��b����U��:q}b\�G�����pP��
tQ+��� �t�=]�C\�W\��+^H�9W9�j����V�X5HA�R�Ӱ��Q���n��YѪk�>?��*{i&N�[��{6+�1]֑J��/�J�i�=��ឹs�BDBm�oh�,8 ��6����X��Ps��J�z˩a&��.�������q qs,�8�p����]K}�*V��ꇏˮFFr����;0�+�S�@��aS�`����7P*�H7	�R��vUELWwB,�(<���
�PL!3px�|L׋�+�vM��V�i�1�wF�#�dRֲܵF��GQ��ˬ�g��A��	Uw� Z��B>W���>AޤܤQ���`]X��Vr�*z��W�}Y�uS��K�TE���.��̱J*�F�0J�5�r�l;y0ߧ#]K�*tcW�}�X�4�A�]�q�b��Æ�t
���/��j�a|���%,-��|;�"`0�(�D��	�:L�ѱ�_UuY�%��n�T|w�����X̿3e��g�z���
�[�c�*�ـ�Į�Pt�����
��))��(k켉��A�G�>�&5QP�eG��w%o�0�i�pi�X��+|Q�s�¯��"�3)��咩�Md���_*�r%��Re��lJ}H��^��I*�	"����$��AIU"1��N�S���姳6췄 ��i�Ƙ[;QU�&Τ`ay�	�Avv���ζv�4�8����ߏ�N;��`�*~*(aU��F�a�ԩ��1o��)�r�4m��z��ul�V�����l��̖'�d�\�}��Ҁd��*�o��䊅��6��蕻ڤ�P2�dә�����W_D�P3�̈́c:���R��v�8�,�R���32��\�4u:r,=
�)T�+��V�lyA��S���zGPzL����F�^�Η�n�m�+�`*F�b�X6�U��S�����U��L����Dm�i��)�3�NOFa�p [��a�&�&AQ(��aj58�U��R��+>�����6d�-��TU����*ͩf@�!�ػ�r)mY����b}SF2�G�^>i:S.�H�\d���'�1�A�UGӄJ�¼��&��'!�Y�B�l�I@��u�p�MG
k�?��N����u����E��]�mɶ\�M3�65��%��M	����#=!$^ �M$$0lL1[��d˲��ծ�uv�̝[��9��;w�����O����-�}��~��6z4`v�DH���oqnn�T�*O�W��Xc��~n��*�A����I+�B������-'XT{��b�<�G�|�L�����ঁ���M/I���#����m�F�,#��Vr^ui�<�OYj�d�[��fvm�yD{�)�/��/;'>�(aŐb�~E�Öw��y5�
f��}�A�Aa[ݪ�U^|��_��C?��L�șa��+��;���^$�(�	�ҹ̄곽���'�[�R_����D4����>�Ē�%��.^z־�z��M�$�(�CZh�N���B�G�h"1��&~43��w��:�j���J)����Ԫ����Z�"�v�Ƽ>�\�}���̧Dv�#���\ѯj�bF�K5u�:��1�WJ�����dT�n_aBm4��BEP'�� ��u�]799���ܳP(lݺ"�� �V �a B�S��~i���C�BO^��8�1T����Νs6��T.�DKg����]�f�Pe�2T� �*���\���(C>cA)�L^��fa2K��=�^�Y�R3u(G�U&�{�[����0��HQ�ֆ�U:Wө�EqsF)nQ؁���$�}�����[bɢG<�0��C��G�����G,����;:���ή/�k��IJ.�=�-(T�8s�#b������f�K�m��D�EW��_�&&�U�
)���Z�8~n*����M���dHn�������Y�?����O�1�F!�&{�rJ�u��Aޛ7oߡ0��)~��s�+���	��b���El}��Gh¬~�3���۠3���7�ft�ު�k��|�GQ�"&B׋ױ}���an_�%�D��G7��D2�/)�ʽp�a�RN���{�7̳����R���S��>�>�\_�u�-&I�K���'����j��ׂ�㟮Q���:j ���h<!J̿'6u`L����/� ��4����D����(��,5����g���^���@B�Q�+��-TAȈ���mLګ�=y<��܃v��q��8�	�?jFݣ� S�I��!H຀n:Bʘ
S��Vw?��V���EG�H8A��$O��\L�(�l%��`H�N4�B	��I"AC���q��,�OW����!��w�A�O�}R��!:��TMJx6H1���	r�o��ʆ�� ���
Y�UE�G�L+;LZ�V�tHh(���{�	-�6Fq(����v�Q�*nU����^��]B�oڴ	f��Y�ѣGq�@_�@3����'����$�O�4���=������Ck~n1���cǎ�LO���z����ᜪ]Ǩ�GȎ�Ԫ >�}	����_NAya��a�-,����=��g!��&0��TJ�`���Рrڪ���x��w�SȨ(��J���H
�1)����z*D.�'�HT^Փ�f�^��@st�>��\�$�qOI��5XB��h��?f,��K�99A�L@jI�4�U�\����r�^7����m�Em�;K���	������u2T��y_,���}qnF��Y������G�r��&�la4S<�z���a6ӣ�G1�N��j��ܺ%�y�9a�k?�(qD�2� �Y�F������tj� �䣀>q[�)u��,�*1NX��q����T��:.��$�y���Ț��(�������g�O��"bgq��r�L�( ��ղ*��⎈�H������}���E���G���{�c��Z�q��3�1���)~����iN�������p��+P�;n����� W3I�L�c�Gp��f�I�-��+2�%KH#�]Q����_>T!q��G:�V�.�p?��D�+�b*P���DVW	��Ȣ�F�G���>�5-qO0Z-�_B��~D9�G+Q��֗?x�0����p��_���&[�Y��}����bM}��~�	�lJ����P�1����Z�E"���i���8>��UG����y�\ �w��,%�Q�\e8�-��J�)��x��4�\.�v߲eˉ'fff�O��4�={��j����hW�G�µkמ9sR͒N�༸�-$:����/�ד'O�(�}}=[�n��k~�aHtI��8���Je("����A��v�؎s��*����|�,�u���8����_��p�#����Ŷj�����$s�V�}ldwJD�����\�^�0�W~ر,�Q�jڧ�-�GK�'�E�\����g���k,ɢ����.�#k.�i�I���^Y���;�)z�&lZpy�Q��/�Ϻ���n
�!%�3L�Χ�P�C4b54��"��~P��CCC��z{{Ax����5=�Vq��M��P�TH2���>Df�w�
�&���R	Ãf\����y?�ԏ/I"�,�ʙLN��/�zcjjꪫ�H�Rj��?�*�\o��_�47��j�5լ����T:�m-���	=�SԄ�[]��j��:���a�0)����h%���5�c�2�]J��j����
0;V�����d��b�r�����W�l�3u�UL�2�S��6�^j`L3��r:�ɩ�7n(�����Z�&��}�zq�X`�d�� ��NK�U��Gd�3��v�̅��e�	��F5f���r�Bǡ�v��P:f���ir�Q7���i�zI鸖�J���pɋ�9��~��B��$�=J8Og)�S��:5+i��s9l�҆�[́���s�����.��M�HHn�[T�S:��+��L:Tt��z�H�	��ױ���4k��bp����	��ɷ��;*`����De
��S��IeRAN �Te�
)����'\�vF /�?04;_���IZ&��W�D��N3���0��
xD~�Ӷ����q���Ж�U�,��4 �Ԛg{���K����^�	�����I�"r���5�;f�]��â����P/@+[~3
��mT#p�����j9��i?˴�NC-M��Q1�e��~)���&#䫮NI�ήT*���n͜?_+�mB�1Ħ�Z�N�j��ˏ��g>��A�T�{A�gΞ ��������,���O@Z<|�'@��R��ǟ&@���|~�B�qg1߅Bn`��{7��Q2ǳ��������gΞµ=| ��0��gy~w0��F<p��d*�H�j°����c��i�V�-�?�0���ɉ�.��_�?_��M[W~>�X�RYSO�����ǤVŞ��G���K��0Q��d�b��z� ~��X����꘺�w�F�A`�Lv~f�R���ӱS&X��0� ��Jh�I�i�����F���WA�*X�F���(����*�f*��A��t��,�|�b���\ ���[T�Xn:=��K-1m�Mr�ת6�J��hA[Ld[7k���������'*G�b9}>�� 09fc�_��$��-�id=�a�5:�W]�������@2��g)6��@�O'����;�8���^�,�Y32;;�ɤ8����b)A>�V�&�gϞ��B>er��m��y��rwĠ����u�J�8U�D�J;�d4�t*�9��B�8��z
�(L�ą���c��n ���#o١r�f\BG����eM9(_�̎hf������#E�"Ь�j˞�� ���*?���y5��m٬�\'�.C/O!�E��,|]~��.;mه�}�g\�UUu�s��,s'�:NeY�0���R�A�S�i�-}$�1n���\6��a4a�pr���%t#,�f+'$$�u�����^��Du�$�~�C]��@�����l�F�䯶AԨڂ�* 3�ۭ�8a-�g�^4a^�j#��O4'�8բ�;5�2�����+
d�0u�����N~�������	�o�����x�J��՘;
v3~�Y���jI�q4x� �o۽�>&_
x�֬T*QϞK/� #��B��UXT���SO�O�~>��߹s����q)h�sq��O?�7<��qmBR#ȠV�ՠ����Hj���,�t���¾�e�&d7(`��A��7Dvm��n/k0��i��b~�#ܸZ�%l�0�Iz��P�v�G��Y~AQ�R��G���~�Fc��L�г��w��)�~�;�!�I�T��~���2�nm4K2��W�F��Nl��BA��=ͣ �� �7_0A�Ν)J�&ydd�jԹ۞9g➠�JJ�
tq�&�y�_ԣOr��8q۬�[��(:αc�0�}��ᆴ���{�We�2݌��#)Շ�4U�Ƃ P&(�_��7s2Ɣ�bP�}+�����[��Q���U|�������+��J�IҒ�j�����*�|�e1X�����j@A�W(��eLb��m��"EJ�\�|�AK8?䆫`��J�wN\�?��^W�8*f����wu6W)�:caD�n,����{�V@���� �p���SV����I}�L�;Q6g����_�ir%�2U�X���sμ3,I�bJ���@��	]�`{j��X$�ͫ�7�wfx���\J�~�����ŝ 6�pJ#��5Wӽ^*ϥ�j�b�-��t�3k}�� �b]@���I�$��4��܎�i�-.��n�	\m%	��nw"!`�D�#�O�O{�i�D���"z3��d�����t귝LR�CƉ�6�/a\~[���G=`��XF�]]'䤬٨\���|��C�N<�����#�2
8]i���|F)�J�%��߱�Z�m6;�tfn��a�M��N!�O��*�����.A_,�!�k~�ݴGF���984ҭ���\�U+�V�8��[vb�����YV����r�JMO_��-ZIsv��L%Ŗ�XJگԪ��\Q��6�By�v���a��������199U���ǩ��=���ˏ��0ߦI��iu�yO��ҲgyD"3 �P#�O��0LI<k�h�B����p���'��r�#)dP��%q@%T��B^A��]� ��u��ǯ�J��ӏ���5��,X$	2��ď��;�����0��G>J6"_�B��B6i����c㣧O��Fުr��,�G�`�K7蝂�.xD#!���I*ʍd\�B�J��؟/�V�vKl�`�	wu�B0�t��]-ȉ�Zd�	��VK��K)�����	����֜��ۛ���v:��+�6~w��0=P!������b4�ER~�:���_6�_� �r�(</�G��1�08�w����K�q�g���1��֣_�֪迡}�KVn�q��'8q����l�`Ž'�2�CE�>�5A��:uv��1J��hZ&��VF���( +�j���X<;N]a�|)i��[�<c�w5�|��Uq�$>�BA��d�GS��i��Ǩ;r�TB{!*p�
K�R���Ʌ�;T�jEf�� �)_�H�����Po_�Ӵ�ġx��<��r���AF��,y"���O��ʫ/H&Z`Qu�e�_��&E���A΍�F����+W�X��qC�\��*�֣�bym�`��!BP,��"@�ʓ�i�����`܃)Î߶m�vffFr�=B�.|CCCQ���c�!-#�eLPQ#I���Yp��.��`�"@�{���n�t�u7~�{JX-%<ɚ���J9Jw%4����e�f�ׅ�Kpڕ����sq3c����D{*:�_�l���Y�~ ����h�*#YQG ]��~�Aa���o�~H\?"�h_{Ks���u�������=zt˖-��9rd׮]x�b�Z=���J�|�gΜ���A9����}�F��:
��B�B{�5@�&��+B~��b��)����-U[-��Ϩ�>�L���/,����nփ��;����pd*z��œ�T&+U�*�ڪ���`��7��z�Q�`�1����6��l�M�����@F�x��u*�P���4��٠�w��n�[%C��=١
V�f�����NF[��p�s��N��ץ�c�)j��M�\l�P��[W�ދ:�1P ���k�3�KjK�JeJ4�[��6s9r�p� N��$���)�\	�yb4���F�ٲ�v�F��-�i'�I	n2��ɟxb�,gM�J��O���Ɗ�o��C���(\����	�P//=ޏR��^�\N�d��;�@��S�l{�K%q�/<*��X�&}t�VD�4����c;��c���2v��X��[5+	���a9�d2�:t�c��:Ԗ�]&m�ęv£&�>؁]����^��H��&���&5�&�U�j�y�<�e��b�U�J������+8h��m潶B����xm��=p�+.�ĊR�|�� � ���A�8	�]� �ݬ�[�Ӣn�����D�+v��Lq}v�Zŉ�LVO��)x��b�j��v�z��4�JfTE����I h�!xx�������q��׼�u`Ǡ@|�70�	�}��y�!�6mzꩧN�:渁��3��X��"���;6OL��ʭ[Gb�v��[0C��<����l�m�	X�M��-d��DNOo�����b�W��t#QgX!��!�F�]�������V+uΔ�X�i�,�gs�Gz*�)�J6mT*&.k+!�b�\Am�"J�������m45�pu?'ʑ�@�6r��4Qz_&]���a�z�ӏ��X�)����e]3f;^dy��
&D�iQNk�P�DH��݊�����"+`��9{�4j���>�裶��3�$[�*�=o�Ν���T/��.w��i��O�H�.�`N&�r_QYp��(G���F��Fh�:N�B��Z����ًo~��{E����ï�G�K?Xn�����h'T�L�(������l�n�3�[�:�,��K��v5�e����2�-0�~�CҶe#���E)�a��;Wk%9�t13�x�r[�g���}^�uF��]V�6����"�E�>�@B�����Jb����}<8*��C�C�J ��ڥu[��U���%K�������S����WPts5��KPH��hb���H�GԲ��UJ�cf
�}�֊�U�`���\�T�
��{n4��Cl}�W��-$�KDsg_W������*���@�)
���:������M�ǎh�]��ӭ��k��+|��#�Y�b�P�3Cz@����.�T	�J]Vt��aIdW��n�+�P�T��'O���}�v� ����CO�8q饗�O��Oe��-�x��*(�����-��xr�ܞ={�f��+N���F�*��r��*��JJ������� �n��M֐�2����u\8�������Uc�����5��԰~RӖ����]"A"�+9#/�a��]���k{�
����s���Fg�\�0!V��c�P�Y�q�h��X��p��e����f葺�6��V�&6�<~@c��T� +�lP�M���Mjy�ʴ[M|�g�r&&&��x@����`
S���R�2�ʽ�JХ�� �^X��)K"����On�j놽���GW*l
�E�������M��z,GZ~��3ZaGU��Z���	X�*��Y���O�L
G��s_M�J�6��jlh[�K!Q���~'dI�>+F�_��%zP|��׍�"M��1_	���p\Ct	,��	xB?<+�ɀ�7j�P�>s�*��q�B)���e�J��\|*�d�V`�쒭aĬj� �2$���H6���K��e�r�/_����f��H���v:0��X�ٮ7[��b@:1T|��B�p4[q:�����9m��r'1Y٬�xAb1?杖�2A��P6(ڡȴA�u=�۵ğ,���e�f2�uyn��S5���"}O��_|�Q�������l�,Qj�N�)�S�ܭ�0�<Dt)�Rc]x! �Y�w��|`�� �Pa���T����H+�n���'�[	t��IT��!'M�~�+]�	���qܡ��x�x�u��P]1�e]u5v��KYP��!���xC��z:���b� �7��!~v��\z~��M������� {V��+$z�x��ځBOr|� �$��]����>|x˖���{/��Ț^py��+��}��Y��Plg��5����E3���)ιs�Z�����!w�];�B��J�ril�.������v�P���3,��]3Զ�ck/�dׅ�*�wf~�ձM�k�ء��i� ����������?�It�L�n��2:4c$��_�8�Y��*����%�د1����Oݺ=37T)_�0���a�Q�q�y���&����}�[H{
7�R\��}#@56��D��{�����F+�9Q�DBg�S�u�VP�¡C0į��ʧ�z*�&�iX��+���Ǐo޼yjj
�`;�� �%5� �E���OH�_@�%�Ko���pI�1Zh����N��BZ`�\
��� ��W����g�!X-JrQX��C��g�ΈB��J��b�	���E����QN��78T/PZ.K�����Q0�o���-?�8��ѝ�=e��F��F�f*H�� a���6�Ǿ� Ų�t��9���z��S��Ԕ�c�f/v�Ѝ+�5����źvS0�n5p_�X��ߨ�t~���A;�����Z^������x�e#TB����{5��V'Hy�����_�
"og��HE�j����_�1������j��c����`D��+��L�r(�oYQY689��0�Pzp��yҰn�G���`Nq��&Va׮]��۠:�ܱ��m�6�m�ڵ�s�}�s�lqXBccc`�sss8����� ����Y���S�zUb¡��W�'` m�mqX�{{{��G��ЬWGFF00\5bd��ZL7�H&���~wVT1Ϗeڮ���lY#���Ġ�dO��\�g��*V��3��6�~^2���aX�~/!juO��nl^�YPa޴��z�r��Ե��;0���ɠ8J��=���&W>�r����SOQM�N��(z�%�\2;M�O7���u	J�������_�3g�H�ԋ��A�=����L\}��WVa2�3�e��8gf8̏�R��rY|ղ%���3��k��Ap�3�A}�-J��_�1�B��L�G�;)A�ZU�C�q�fS�`�Z���S�|_��8���֎o:��A���^�þ �׌N���	<;�S�;=6��,Ey@ݥ���M��°R�g���H��|�Tk�PT:�贓-ۄqԲ�d:ׁI�&��������K㒓Ǐ��Vj8�p��d��q	 ��$G�T-ڎ���	�@t�$A~"�69Pq�K�$t�DJw�J��OQUI�5=E�d+�G-���ӳ��(���V��h�6����0|5�Ζ(��q}��h�펄�f۩>���fL\���nz�L�{��V#a�+X _թ�^��6D|I�N�4ŷ�s+]�*�ee^�d1�����վ��Z��U�{���n�@�V�`�vw������YJ945��1Ƕ��'�eαr�6(Ɯi�x;��0?���y�[c��L&w�칄��),6#�7�!�l�D������F�����V��.i�� � =2nT�M�ڢlw�w�3�A�i^�ﴝ���)^6Ҿ��ʅ=m�Xa�M�����JXY��5B��L7���\+ڨ�RɎ ���Mr:��*�.g��DM.�˾��3�O-11�uq�ݢl��鬌��nB�>�+�V�1�f-�!ܫ�hCI��d�,XKЂ�y|�ޛn�V�~yt�9�q�HZ����o]7êC}p(�y�l�����k��Si�����[)�����M�mbB�9��5C���n�Yk1��
��c=�к[@�V=9=W,�v87{|��[6�S`�=�����	�S��_�jW�g���(֫)y�l��s�cB	B�(*N���-J�ҳ&qpU["wUq�E"S�N~�@tn�+_B��]hp=E ީ$�s!3� �y���J^��])�P�*'(a4O���F���K-ש�vRGq:^�QO�	�v3�2��HS��l��	+�U8a*
�IdM�6H�@;�h#dͅ��Y��L��N��6�jj��yt�
!�L�?	�"L��񔫮����zAu�Jz�Ț1�md&��BWJ� ũ�G�$: �+�K֬Y�s �E��>A���Z����~�l��:&'A�N�\}��k�������� �Un5�@������R?n�:`���a�#Oq�>�
��\�@�.�HD��Кk����y�ѕW�ۺu�"�k]��V����V�S������g��"���694�f����ɍ�g6b�Ê{�1��n٬c�Bv4�=�]l;��\�n���F��������ϟ9{&���P�!����˶��j"�ϭP[T]ҵlԋ�
�X)� �/�Pum~~������TB-;�-���J(�#���;�����ڊ��"Ư�,������QzN�j�Y��;5��s��%�+ƃ����(�-���!����b]�v��C5���1���ڣj<�a�]�dc��+)!��B)��'ƶ��n��Y���J ��l����c/�<6��2�i� �J����Yz��b[�K�\���M�LzA��{�A���g�ͦ�8T�(̭i�1N�HG�n��vQ �v�|�.!I�tk����"��&�F�Z|ƕ4Xn��NJ�%��R�q�Q�GM]p�00��wxݟ{��a<	7R����QOR,V��V�F>%t����[��̓�С�M%S��Xk�>�Y�O��{��۸q���G�U`rA��` \~���ݰ=��0���'s-� ��L�٫�3r���X�kHôБs�+�cճA�#~Qwy��25n�sW,��u���r��STĄA�0g�=4&B0��H��wB�J.�z<<U�*۾e����Lrģ\��`3�闽��;-D��-��X�0���,�8�ͪd���7o�eHz@O�^K	��� ��
���w�>[�l��\���Z�7��%i@<�8A�@�$6��<���c�a�P���Y#�+�*O_Ʋ|~>��'f"9t��"Y��x&�&ؐ^�H�{����]��w��K/�⦛nڸ~������� YK)+92:v��h6���W���\����Gm�]�6a���^���3�uR�u-a�a�I��^�M-��ڒ��8����Ηk��F� ��P32of����	gΜm���W_}��k�QЈa���޾L��}��;���D��OcKs`���?;7�J�t��`�d�	��M�Ť��ĵ��v��L��{�Ӵ;�v�<B
a�9^�T�7ں�Ģ�m��0jt>�+,�k=�T�X���-?��{�����<��@�%\�p
��s���[�Cal]��sG>�T����L����a��؝z:�M�n���/�G<�m%����X��t6S�/v����'T��G�"&m�	+�p��c�DU���s�.���U�
��_%�v~��a?7�h
Mۏ����E����h��٬Wk��㩉�k�[x��,�؄�d�`� v���6!H�j��I���_:���`�[m�0ֶ]Rm9�EoQ�?�Hǚ/Wa�,��	5�I=�޲km�dɔb�A�G3c4�G�b��Z�waa�J��@;�p�Lɳ�V��Z�`�N��m]1<�� T��~=�yMW�$[>i�-�,qTJ���,1���)��7�i�������'�<r䑨�*JVB�!~r�O�dȿX�|i�X�YH	!7��}ו\0�q�F�^�Ř���PY�:n�47�"��t� �Y�<���p�/���~���]5�$8(����#��e�˥�Nf�����Ir���B�����R��ֲ:b.S�FrL��O%f|�\Iw�0E?H��{J��({_��L�6��x�Wt�	͗��C�Y:z�����y-��1B>M_�8���3\ J�4�Ћ��R�����|�h~��*W���I�,r�SmH��8*��A� 㧉Wk�f�d�j-��*�FԂ\����J�^(�*�q��9P�x��}J[Z���;vu�'C?H�38_�;L\�/#ǃ��D�b�d�c)h�Q��4aQ�j��n۶�O����_��O�C�����02)lU��V*��>$�W�m�E~��}��y�@���%�r*r٠�p۶mx�ɓ'��暹���<�P[-S'e�4M$�RB[p��z��#���0���z_������p=7_�e|�u�۴y+9c��M�ZRmxx����# ��o���_�*ؓ�j0�O%ŝV=��3�z�Yߺ��Q�P�U�B�0����59r�I�/x~�a$ɝv�ܟ����|h�^���[�>[��ӝ�J��*�>�\�aã��T�n�J(���@P�B(����
�5�9�Bi�'����T&6�Oit-��@8�Kr^b�F��e���^A�Z�JdC?~�i*�$���TN��<t���~�/�C��w������d��H~�u����Aa �a��7���p�~C��)��IU��jz�%=%�ح6g�p�l�65rK��~���G�Cmi�G�q	����n����*FE1��|���"��Vu���h[1��t/�A��(�Y_| �� �'�ha��N��QXh	��ۮ����~#��w����ưDOg��IB�#k^}��O��"���N��>�i�7օ�eht�	����r�&-E�0��C �7���ì�6�̕�sN�R49�ϟҢi� }e�\���˾UC�pyI�q�%u��ɲ�a�9��)����������_Rh"];��$���b�Čf��&W��a¨�}樮�Y#�v/,����MbZ�z�e����?�6䨪�i�s�Q�@>�)XY�zpsI:`�y-T�
���s��)���+�8z� �I����K���R� s�c�K��p��SZܶ}�|�����ȑ#O��ϛ�9�>�mR�\Z���gg�-�m.������J�"~�o'Si�!�8n*��u�e[6���Ӿ�,Wˆfe3� k%���?{��ӹ�z=��d&��w�O�zs�Jr	a�[f��Ù�����=�N���!UJ�!oM?�'�"j2d����tZf*�
]��|��㐋/y�+.��2Q�\��հ�_U���h���ȅ꣇Ͻ��{av��;ﬕ���� ���	6H9#����n6����]���9T�Ho��q���\�5U#s��i��n~Ջo~��R
E�<�n6��G�����0PA������g�>~�'OO����6��z�&R��:Pb-��I-�@Η��i�B�p�GiT�}��D�W�5}�N�U�څB�R�5p{������-o׻(o����D�HQ�L#��������?����HX��Kݬ�cfPȠ��"<���ȣ�|b��'��Ƶ���S*/6�R�sͶ���3�׮���?��5�m�����e%�͖w�����=R^ظqc.�9r�i˴(�Q����!�K8_��HZeB(A3s�_
1r7��R�N5۱�a�ZoE�ġ��,d=��  ��IDATT0N���ɉ�'g�͆�Lk�f�i;*'�ԪU�3kՎ��GG:���|%�KdR�F�I�� ������S�b-_#�\���$	�����C�'lGW��7(����n	�U�cǏ�ݷ�M�'G���)��O~zί�OF�&��V��%iPA�1�,��Y�H�Gf�h�F.� �Y�ĩT��m�Ӝ�:�V;�d�+�dj�<�PiV���/��w�;��}��O��v��\�t�����6�l�s1�k�?ͩ���iP�+G�E`��D��e���Qg#���¹DAJ5ӿ6یzC?�ԏ�Hbd�.�b~��R���T�)R_71�dK"kJ���u+]L6?��!�)�$�a�� G#��<꾩J���\1��S�]�e���~��ZDbR���ViP�>�����[��'���+�7���2;;�i�&|�\�������������-,
��/���hj���}�'R_z�Jo<ųW�0��6�ij���ba�bП��g�����RE>,�T~.�/�=~��`��n�j	���F8��ȭ��)�d�]�=:��+DI�`n+�����J����]�:�Y۽{7l�C��Ž�
�2A�L(��7Sr�M�W�|o�=#��嗖1	�HC�,�]�`I^��_��`�T��Wlǲ��M7�F�i�s���=�m������������#�d�������z��_�C�*����'H�m5�ݓ� Ȱ��\�����k_�+��(Dْe�Q���z��%�qC�3x���ǿ��<��àξ�*,Ve3VcpxQ�%k����}v��%�z��	�]|	�QS)��l��y�kn�����I�!�PU쎝0T�j���'w����s�gV-O^r�%J�[Wə��M�=fIZ����Fv�i,_rD�ٱ��[��_9����_z���'B��RMaI`R�v6����{�����>��o�8Nl�+����Gv ��rm'�M�UC�Q
7e@�S�0�
��S���nq���`GTk͙�ʛ�v;4'��'�u��}l[,x���a���<s7�rH�S�<����E�����I�t���c� 3a��MMM��0GXf\&��)O%��X���o|���(��^A�ԏ&F� �ɗB�a�5��2���A#�Gʄ���?��\�~��LL^G$��'�x�rS:�.\�爃�IHezq��'��ꪾ�1�C`�-A�FmX	���*`���E~u���<^�k�Ė�G��ف�b�Q��yBr��D��ԏ-���g%�y/ـ1�O���%��r��5�|A�!�(�Y���K�v��Z�� ~��5�GW��3���=�Ε�:0XB�,��㢨�Z�Iudd�ptU��um<��썫C�b�S|�h��ѣ۶m�}��$Lצ�w�#FGGE����/�=ו�0�W�/�;DSq�coap3S��߱cǱcǰe�%��U�ѕ��������}$��֔����P)��4aJ�TcjZ���Uj8F*������e�ã��X��|�ol���'�O��*�V���X�)]�yֈ�����q�f��p�&�[��kx:�:�1��3�t͵�ݽw���3YP�z�c*s�b1�kJ2V�dM}���oN�U=�$����߲�ҫ��ݰY}�;����z.}�b�S?#Oײ�lѮ��V G�[mPQPO��_����vRK�H�:J�֑d(��>�Je�Z���{7m~��~�Ԟ�_��ϟ;
��r�	ր!�z$�\jB\O�	�i���X%y&��f�m�����3So8��Kv�����Z��6�um�݁�F��M����(��S:�إ�6}������~����~:�RSj��"���D�{u��ז�meEn��2��绢�MZ�"T��'��b~��/x���?<�g-�]`�:�H$���Z���b����7�������o}�ęs�V}��ͅ\n~��s�/ʔԱ�.��N�c4Xv԰H��:nF�Td���þ��q
��f
����|��t)�2u~��Px�+^�ɿ�����)A���=���^��ve~��2��X�٢4?��h��_��WW�{%����u����l��l&�nr:�k^����lB"��jC�?;1�+�O�<���S�$�M4��da�}����:�:��_ D��Rݳ�@1\d�)�ٳ���zȷ����],~�Y��qa����k5�]�����y�)��N�뜟<ד�j�R�2�L�V�����|�=�ڭ
6Q�uAIhB��g���١V��>/���&Fu=G��J�{1�����èOqL�ř�tX�ï\\�����/ͷ�� SD"����&�Ӫ��l�)�C�y��#d�=�d���S���� ���awݘ���\	��H7�6m�Ґ�XS������l�B�u�����[�%��t������iX&O=��@y�3t)+ŗ�!�ؓOş�0aw�ʱ �k�>�����SI�6U}��G�	Ob||�o5}�.��asm߾}�đ`�=/Z�g+�E�\�0e��a��g�Pҳ�6e���sRa�`�ضy܃b(�i�r!'��WK�K���[��X�=y�$v6#9��(4a�ϋ���{2ox�B���x���<�W�g�^���6n�	h@_o��(������Mv"�ՕWR]����׬Y|�̙���eҍT�[��I�ÿ��F{�b�	�v',pPI��»�����W�b��]2�>q�E��Nv:��j�_X�>QV����)}xx�R��=�����}�����_��W�nTb��"'����u*a(����@����L��c�����O^z饿�淌�����������T��!���ݎ��ĺu�` =���7n|�ͷ@���׿�M�}Ӗe��%�a�V���'�a�P\�D@������}�ӟޱ�z|�jRC���*UL4���@�\�r������|������~���M)�7bک|�E��0������,��Fǈ8r����Czl	u�Ej"��a`v�~�׾����/�K�*u��UJ�2�l����w�|�;6�~򓟜<�����H�D�т�Y-�t1y���wvV��
����J�׽�uw�������ν	(��_�B��?��{�v:��?i$�%�D�9*+���×`�T'R,�`��0�6^$)۠AդPt�{H�E��j�)H��XW�pϻ����Ư�땩��'Y�ӟ<vj�̙3��i�١ѝd"�^����A�m�5��s}Đb����#.��Z%/l����V"@y�Z%��Ws�>��Y�~��7����&�q)!�pֺ`�8�FTv��	����H�����چ�*�8���XY,� 穜924Q=[U�#%$
�Ā\橷r"A2{�DMn��!�%AAc��L�w �`<��An*!���'j�����/���|+'��Cg�dJ�O<��e�]����5ө<{�/I�/ ��t��ɞ��c�N�����k�:SMڔV-���'a�Y~�'t$���Q)�OA\W!!�+�z�n:%+��?s�4�b�eB��(:f �L����:��*v���t�6��Fm�#�[�R��u��P�<�{T+T��W �K�M!����9����7�.��v��ے���v,l~L��2jP3h���2����� =��AG7P��H���`g���
�o{�����o���{��CC9����V*��ͦ��P��C�ώ��=E2�dلv��K����V�}���l��Uo��W<'Z&h�\⤒F:�IK��dM�3IJ{ �@KI���>rl^��m��䣻o����������r�J�Hi)�^7]��y	�U���n��6���N����7Qȃ^+mf*1v_�����h���
;9`{9�	�����F��JI���ۀ����j�9�f]�841uaf�۴i߯�i�C�>���v�ھ�ٲ[�g��r�kP�83Ce�
��Iഛ�'�U1��lia����t[(W
J҅�i(=}}���?��(�M����7m"؍��)�\J�m芑pfb���׾�5���oy������ۿ��������ž���J�A�5��΂���\���0,���ZR�}N=�R�v�6f6���d%8TSz��	��?~��W^+��!iz�ϝ�\Z�w��v����[;����Ν��>���c�]w]Ҥ"���b�;��4e��:��m�C*�Zf
�M�8^�r�!l�|i���L*�1\�1l����Xn��>���W]u���GFG[vsfn&���YX�45���%�:3��_��G?�����}��z�O~zpll�vZ��q5�.LBU#�>�6u<_�{<�0����b��S,�Ӎ13�J��*�Gsf;hY�R\�O�,�hpT��v��̡C��S�~���9{&�͂1�͞۸a�����O����n�������G����tO�^�k��U+��LoRM��^۞8�(h���JR,ϥmn���g�Q�A�	0S����9a��n�}�48�K7���˝��mg||�Zk�����'������OO/���r�ȑ-[��:u*�ʞ:qz��uc���{��-���e��T2�nְ��C��=Ŕ���YoZ�p�$�GS
e;�8(�VS��U�ˮKՓ�o�P�m�6����4&���jJ��q�J����|��ŎV۞�Q���j7ff��������������w���1BBHr�X�P�l'Ê��� �8��t�Hn�.�u�X<~�*���Q�ƙ�=_ZX�\c�R�&��
���������;��z���z'&&
�B��w���Zy�7��9s��̒o|����K���l��  ���l2�n6;7nM%i�1��$s��7o��s�J*��zN�.�>�n�L�Ӂ��ԛ5���*��j:�'`k֌oذ	�Z%ѬcjȽ�,������X��@�g)2��av�)P"b:�Zq�Ĳ���cfu��
p�o~�?��m�֝PU�6��b9���Ng�%h���u�,K���Ӣ�J6��4��6�2���H/�0��-�o���ѱ-2��T���nu��ӟ��Dp���g�Ĩ��aK_r�%}��	��}��`dd�X����=|��-��zݵ{��_��ԩÔ�6!?L����D飌���Ing�iEE�[Շ�<8����˯�8��RI ��=�Q'��
�`�8���"��\�&)�=B��iӦw�����{�~Z��p�[c�(���!��Y�#�퇆ae�f�q������b�G��8
j�R�=�����-��
^��[�Х����xY�M�׮Ì����o9)�JT�����ÇG����ٳ������;��\8�C�3�-\G[�:i����S!�����g'���
·2���k׍����[��6ai�$6"^�tg+�3�����+��رc {-~�җ�t�7|��?�����տ�*�yCCԔ��063�jJ���ܿ\�R���*WG�{�{���<��|���?���|�#XgXt����q�vMs'��_Ȱ�U���zx���;��_��=�����ߛڶm�bu�q ��8�%�C4E"SL�܆$h��O��$Ƀ��Eӫ�\�i�].s
�0}l�c����aO-�J�gf��`JŒ���ј�6����ؕ�}��������ا��k�2��Z�z�2���J �Uн��e,;D���p��znKL.��r�l���`�/y�k���|_�����#O�_�Śn߶�駟޴e3����'_���;7���?��+��bp���1FC�<,ϣ�g�6��u٦�����#����k.'xb����)�,�NI#|Ӷ	Ĵ�O�.��Έ�%~���ڵ���S�260�}Zżmذ����G��w���������iB �$�Dܡ�8-l�䢀�����!�'Wcr.��mu��0I����	w|�9�y����Ν=O�(�,Rǹ������/�q����!�Jo>9u�%��4+��/L|<���s��T2��7�6i�s�؏X�6��a��D�a�ȗ<8�|��,.Rv��-��ظq㱧��1ü�/����Hp)�s�xY��믿޶Bv931<<l%��.�*�VKp��;w�l@*Z�q8r�a�C�rH�q��._������
gI*�zVR_"
�7D%�T��Zĉ���ޢ�`��e����{�A�" �ry�X(��s^�16��聟<y�G��/�S��~�����\o�~�����S���M�������!�9>{��'�s�ֹ�	Ȇ��S؟�L\�^s
��t���T.�qݙ)N�T����|����[���L.^�Z�	��at̞���l��L����Yɔ���q�����K_�r��Ҹ��K)���%��L&9���)<|��5#�w��]'�?�����S�sX�f�\
��a���V�ښ�Y3��Ji/�<�Vo�ZΙ������/��,�%.L_P|$���$$�n�ܹ��}�B6�Or3�0�;�b��ׄP*�]��v���������w�}�}�K��y�g������ƭ��B	���GY`5{1]L�����*�g0��;~�)&[Y��Ç'p�m��
:�����y)����r�qٜr��؝�>�a����y�f"a��;N��l�H���i�k���w�~�s��?�c��Y�֫�"��b������6��{��f@ѕt��V�k6׺�I�Lڞ�k��O~������7�����0wln�F �O�H�����$��Tܡ���'�sM5J�(�K022t���s���۷�G�ԧ>���Ǡ405���ӧI��>,����2� �JX�e��eCZc)1�`��mlf�S��~������[�+��a�fKsX��\O0�j��]�10�ƴ��Nfgg���yw�������뮻�lY3�?�87e�l��i�A�)5��zb:	�Oe�v× ���A0YA�n"g��a�}7A�����P��U�}�K_�Rô�h�������}�Q��4�k�W���];6������r�-?t �����#{�\�v|<znzWe�T��j$,o@���(��{ur�ƨ����Ju�N:&�כ͉��������������K0@0����!0bvdx�B���[�����у7�_����o��o���������/n&Ӑ��}��N	eS�}}싢���ԗH#]�s�sg�3��c��JUV2M^p���何R�h���W�#�S.����/~�u�S|��a��ğ�0+�yN����6o����]���ཝ�ѷvP�����Um.t�T���qL#Av���֤7#%"��V�9\�J� +St�t��x�v�����R*}�=���6\����7�|��C�r{����c�{�
��"���ƿ{�}7��Ʊu[���/��_�6;M�K.S&i�0p)@����┌}����]�
�|��r���ھ4�PԎ�4�MP�t��$U��{�1Ga޴�[Wk���5�\{��n�T��{�8uf"_�7��ʋ���N��OR�L���:=�A�L�لe�G��r��氮R�/5>k���ZN�
-��jE����0NOY�n݅�y�#H���)�zVR_p���PL�VƘ������7��Y�W�QJ�!���-��J����$`@�k�@���_w�����j�87��a��S��eOL�_{���:C��耺@���yH��]ۼy��G��M�OBWp�j�L5e��7�O<9��c�>�6^��h��C g(�b"eM��F�wlX�v��4�M����-���䶗��R�S�5:�� ��s�ȡS�N]�w�;��λ��M\�y,/�t�y �w�b�^�l�(�����-�Dj�]��8a����f.W��M��}�O�ç>���A��-oy��_��]�y�TL��n�ف>N�:s!�K@��s�������x�@o^����T�9��{�^v�Q�vЛƅ����b۞��㉅��.�:���k",��|��\�v-�j����Ћ��f���X(􀨰���(���[6��?�����{�'�PA�f�S��Nq��4bM�¾�P"��҄/,4q��gν쥷~�s����ﰰ�֪K���cTm�c�P��CNA�dw�Q���l�2u~���*�+_�ʎm;������o������}�k�P9ґ#��R�+YK���i�Jx�'=�(���x����8~���v�m��{��kď37� K	]/�� ��J�L��P��CA�\��ۨQ��g�6���#G��-�|�7���O|����s��C�>�$)��6A��.�Q���|��m6�e�[�̝}衇����}�s�3�n3X�C��&	�srj
�2�]��!��Oqtt���a>��������_��]�/ٰ{�N��̓[v$��9u?(��7f�A5^��+�h�Qe�>�v2�N�}��Ck���Ͻ�o���N��f	Rņ��ߛ�
�d�q�Epg����о���>���~���{	䪘@��MyE�
�Ce�UЛd#�.U3jT+�I��d�0�^\4�2*��ǟ�	��Їo���V�r���gh>d��19y~�֭gϞ�7PA�?�? ��~�����~���1�����9:�t 
�/�����ځUM��P�/�q�
�whVp��=�j��o݅�ܸa���+Ro$�J\r�G`S��-�?���|�4�C��,}'�,�SW�Љ2N�H�$0;�`א:eYC#�=� 9H�����px"�u�q\�3�
@�X}l������&�����m^�A0T)|c��-V��'���f���o�}�44`.b����cu�^Ͳj�5����)�b�!+��z(�R�w�)U���PY �]F%�
C�ag���,�z���pN���*���4n�e���=��O�.�B�U�|O6YiWX��X�*�<��������e�|��ݻ-+�A�F�M&�<�u�)-�`-��Ώ�y�����ͥ�]qr��).�����];w�������1�p<���
'�l'Te��leqo�~�ئmWMN��������;v4��C�U�g�ju&��LNN�#����-m������b�/ݳ�ġC����e7���~��T��oܸ�7�ӓ��F�Uo����r@C�0�1/{������X�����-������2���!}�I|�5����v��w�D����?��[ny��nx����n%S��H/,�O�IF���'�?���ݻg�����ӧ��z�)rS�P��q=�}�6�d��ff���T�͗�g&N�ܱ�=�cǮ+x�au)���I�3-�=�|�Z9?5�,泐���I���q����5l߱C�S��SI��V�a�(�f�h��cG��n��7��%�����	��VG��	����fW�K�n��)dSI�1�z��-wv���o}��o�ׯ�;�r��f��X�J�q�"�t��Um�j���-���{�w@�7��l:���+.L_X\��e��^�L�34�?:2t��,�*��;�;誫������6R��l��)�N�������g�����F�z������;��׼�|i�r��	3A��w:
���cp�b1/1Ѐ�~�j}�o�X����tf��u������_|�m���W��կ���*jW^q9UƎ���oq�'�3J���uW�9s5c�d_�M[/ת�L1�:sz
O����?��?S(�K9}�\:�+�$�-�R� �)ঠs�=VS��<W��x�~���_��-������ߺ����=_��nLE���VSڐ+����i&�ݩ,і�%��*譺�^��a���������t����ѣG�����o�]!e��Ȧg����ځA������x�nJ4!]��@�a�o��Ex����(4���oy�����}�g>�B�`d�b��k���T����aB7�Vrq�B�\NZ	n���J���+��0%1'�zO&�eۙ���|�o�&�)P���C�H�H�ڶ;;7`���$f�/��T9u�����uw}�{P��[�z�o��S��ۧ�xl�Y(�?}��N��T	 k����N53+��	CO�߹�ʓ|5��E�_pZ�jPV�v^pӫ���E��GOx��ݳw#Ȼ�n�I��駆�uůVt�3S���Ǉ��.���[/�{�ɧ�<�{�l�}��=��9n"�=�>��:�G50�H�1�(ẅ́}ߖ^>������j���4����X.�_�7�;6�q�W�]�Z�����Ng�M^���>�s�N+m��J��z�}�S3�Z'�ѳYXG%��@��KG0zs���V0x���	����o�� ���Z�u����bɖ[�ӈ~�
�A5øN&��Ĝ���್�~��K��K�9��KZA�!N	��b��Hj���-��&���_�җ(f3>;�]��V_;����5��;
�)U)�+��S��߆E���k.�uI��x.���y�	�ɤ!j8X��zՕ{0��~��<|�0�/��W��W�6��f�(����a�9�X2l��vP���W���ۿ�_wn'����kv�P����c���c��~��+���O"?v�����f��������{�u���C~	���?��{�Ť]q�0���Fj���(ԇgB7t:*8{�����������;�������A���[b�%�nĊ�D�!P�`�N)K����;������<gg������g��0{�ާ����=�;tb����bn�f,�{�7f� ����9���'�|��7W_�炼�;�4�"����V]=���|�9s�tu�mظa���'�|�?o������ �p��>�i��":�O$����C�R#�]r�%&��L9��-��H�:VqlOoOsc#�w����׿Bt¸��C�8���iӦ]tɟ�'h����mN���Ņe �{2����?^y%����PK-��V��Ex��p(!�]ڱ��w�=��֛g�y�N��1 ��`��E�i���Q?vĈ���k͚5����w�7̛7�7caD��(�k`�q۝�'��7���K�@���M2�<����!?U��K�������x��C�� (��;;��"D�*Lvʔ)6�eݺu[�l3f̂��
�&��q�#��X�Z9@�o޸��(oљg�8{�3�<������`�(���n*�U����C�
��R���%x��ruԘI����"�b�?�����(������1ŸTTy9w1�p �_����i����;��N�	�?ҩ�"B̢Kr��h_l)�X&&�	�!Q`4oذ!�P/���{��J-v��)��M���/r�X|�`ow�&)���HRG��aÆ�$�_�:������7�x饗�^9����J]9H۟U*�q�k|*J!��X��e�������g��}K�,^�re�bknj�Eb��AC�0D�"#��c�0$,�g�}	É��>�3s�U����׿~��g�(�U��z�~��l�2�H�ұv�u��R�����Ǐ?��Œ�:|���F�J��b�A��^�`�cǏ�8f�h̨��0Mq��E�)�A-u��y9D����i�����ӌ4T=�%u�)<f2S?�J��M�8RWV���m����4ȨQc�aؠR��y	J������*\�eG�LéZx(66X��(���Ʀ�����1h(��3�=F٧��%�9�� �,�OF0�V�cي��D�/^�t�L#$^��f ~Si�+B���o�kGQ7�D���y�֟�x6��r�������*�i��ʉ�":�DV�!�(PRM��������V[[���S�	��%J!��P��x,���"����*4�P64!Y6n>8b���=x�9�,�D`�(:Ѷ(MꍖI�QU�vu�wt���mTqQ���//{�0Ґ!0��V�U��wRn�h|�K0&kJRV���?��h�����b�S�-x2�*(�*(��;|��-��??O<��s�=W�Ŗ�\;4��{�Ν����=�L�p������$��h$�G�~&@j�o:i̘a��Ͽ��+����u>�����H}��N�Bw�;r��a�O��;��rs���E+��=�2�FJ�a�>H�y��b����g_|u��*�aꮧc�@�����С﫫�\v���i�p���%�n�jcq�7��~o�=iܘ1 ��?�dŊ��
��;��j�N������bƴY��T�7�$m(�p����c�G�J+}���?�`���x��!幹y����?�U��~�@#�0{���~�*Y�q��h�G�E�`��IV���Z�`�#��iu���������]^y��իW���+�^op�:0R��E%%Őz�R���;���r���?��s0'�[���Ʋ��29�|�w�}7T�M�C3#%��h"���ظ#G�,^��׬�`���6l����;rh�ҥV�M���
E"�m��tR���Y�۶����8?q�^x!j���rq�˞�N��d<F�+�A���0i �#�&�U1��m������+�N&���	`$}}>/�tw�r�
���tu����1"摇����A���&���J�'FaA��4:_0��;�ƍw�}\}Í7]{�o�1���WmV��I	t�̡�AA��(T�֦D|����ra��a��~��eUUIY��������WQ���@��$�B>��G'7޹/'�ԣ�����%%ef�����?�5j�렫n��vL��8�O��.(қR��Pwg��`4t�xBk�
qJ9�:�M���Œ+�/֏?~�O?IҞ}��Z���W=t���ۿ��{PlIiQ �;��;~4�����WWWp�����5i�7�Y3}��q�G>��?��|L���a~�}��|Y��$�t�;Y��������G��XmE4���	�
)���k�����Ee��`���}^��?K�H�V�(����s��P�߭���fS^�/��݄Ŭ.x���l��>	d2c���U�"�b�άs��Sa��:;z�^2��`��Lf�/��v7~Fk��vtu�=�~���TT+(t�%��m��|��Fuu����10��QMRk0�pKk{UU��j��g�>aM&��6�"\�H��PN4��c�p�->R�q�'��n2i���Hg̾l�ǥ}��q�q�:�!:.��+���ß1�3�1F�}�&![����V�����I�In
(�Z��ȧ\�}m-1&"ВE!<v��%�%�q�Տ쭊�&h�p8��޴i�Y��xٽ��%��t���YH����瞉��k��?�`����$�'b00̱y7�t�?�F�s0Nr�a��b��W�6�H;�xsXz��w�_�ᇗ�p�����G6A��K4(u�ট6aMn���%K��[p�!>>��Cx0e�t"EN���PQJ:��Ӆі�U`$ &a#GǕ��]�gӦ�I^~n]]�Vcj�3� �F#�e���駟�x���^{�Ö�O7���9na��]M��;o�����;w��7]�r�':a����44�Kʬ����t�5���Vt\*�-*����>xj�j�Z�o��ݽ�v�ȑة��N�'��F�
��Q3��Z�`ߕWPR=Y�ℕ�R*e���<�W��ܵӤM.X�x��S�yꩵ� I1``�*$(������AO����g��9�x�	v�
I"Fr��Ċa�-�x��{�1c$V���0D; ��k?��Ӑ�C����=O�>�!
��]�?U�[�����y�f�����Xl�b0+1������y�����]��� �aw�+�=�\�ߐ!f���O?��sx���c�\��G}t�]��=��H���)�GN,��-V�����[��ݳprM~V���W_}����b:[J�EP����-�[NQ�Db��]g�u�Y����?!v�P����>�ɀ!a�f͞�+k�o��q1����?��%Kr]�H8=��p)?aGj4�V^����M3f�x���o���Y3j��^Ǒ�N�����?����݋�_���g��3�-[�p�?ò�)���ׁ��������s޴�ӹ�uٕWZ���%�n�N�®UUWs26V�������A�_}��f�9D��R�#ԟ�zψ_ExMZ��q�7ud��`���V�x�s/��z������
K!y`�^llj�C��v3l&��aذ� ���çH�o[k6�Z2��"7mڈ�t�I'ϟ��c���#��ˢ�2�����R������G������>� �ᄦ�����Gًz������t>N>	�͠�֤L�lÎ��c�mMTl�Ny�#'L��n�n�>.��i���3���*��vG.�@'$����a��� L�scLf�0gΜM�6U+f�>�{s;Wճ�k׮)S���V�H]#f�?�&M�iչ\zs��!�����O��/cEȓ�6ry�IC9�ޑ��	���\�B�:Q�(S�װa����~f���ʋ���J�s�(�"�T���^�lg�	d�����-��`��h��I����H<�F��i5h����D�J-�d��B$��O�ɄL��d[���8l�]��`q�N��5R�
 p�?���&S�H�I_D�2�B��Ga�܍ǂ?8'
c�6�e�{�1HI���jd](�T%%OR]�3����� )^gH�rW�V��j��K7o�r�'^v�e�����R��!ɉo�����rHQ)db����l���U�_��㉤NT;�tt�,�f'~��6A=�?����ܹ�@��\9�*���V��tګ��J�" M������U)�Ox�pJ�~�e����_�r�~LD@��hP�"���cɘ�椒m��\W�2lؤ����?�yt�C��쯪(}ᅿ�a��q�&1�ay)I�V;�Q5W������GO�����gw��c7
�ׯ�谛E�84Q��ܿ/�X)t�~�m�����۝��?�7��aJ��4����Js"%��\y�?_w�S��?~��5� $8�#G�[�쿦L9^�-V%�R(UV\��$T�i��)�L;!'����|�_o�ևYZ�b��%2�	ˠ����_�b�ܤ���G���Ұ1Av�(�Ħ`�v��=��U�V�\��k�7B"P�@���z\����s�[̚��|��s!��[�'��q�Mć�����_N�X6�*��ʣ3�3.��/���kG��,.*��>����Mơ�0Hhe�ߛ��:�'�t�˯��˯~<��pCÞp� ���k,�4l=�=��㎻�?�nAa�x�"z�I^�=���[�(9��;�qcGb��m͏>�� ��$�r�~��o�����C�@u�(e��^��nq`Y�
<�B)�ܰiK^��tx|��z�?_yp1t,��0�h���bdx$̢�3�"�׵��_���uw&ljj�ֻ��<��j1��A�/���6�Ps܄|��H�x�U���#���'����'��H�N'�Ԓ��>����WP��ex($̑�F���U^�M'/��_[[�1�-��B��"+QU�1�̽}�}Nχ��Z[�[��o���o��llj����U�R�6������8�9[�n�0~쳜\���;�y������ſ�$	5Էj�����D�h�mji��Ѷ��;w�U�={�57�}��e�ܻ������(ͬ��t�,1�Mʁ5�����Z`9�HL��V���	ݒ�Ο:}FB��54t�wӉ��E%�Vc��@�S~�I�s�Ǝ����?��CXH����$*�UT �N����~�)���
l��`���O<����a�a�S�N�g�:BQo8���ḚR�d�'t�`J���`�ϫ��"����52r@� ̺r��l�:��s��&g"��'���XԿu���\Snni �bx7�岦���v�*�?~8�,�ܐc��=#Fknj��މ'���C{r�;�̦�K�ټc��LUZ��q�"e?�#=��q��_�->�}�`�RDv>��+�"�_i}�>8�V����lh]J���{Ί���/B�C���)*"�7!c#,4�4N�3���6*��̩gJT�b,�z��������KX�%�%�v��"�����Kͦ�NY��xZgW�85�L�2�ްaò���D⹹�9W����<���.d�I�J�2�
��QP)�2���^X����^z����q�$�ӈe�4��dd�>�#E@>�c'Z�Lss��-ml�a�[������~�Ic��*����ف�L>&�����9M��N�:�]�v-T<���>[��'H�����B��tu577�#�SO=u�<���]y�&+	l�t� Mf�(Y����2q��Y�������s�`�*�J鬤����	(_�N�UQ�b�Q2WqH���.����;�E��Rڶ7����'@�5��N�Pb6D!\�^~����6e�X��Y'�˦�χ%�<yΈaz�f��\�Kx�Gy����'��鷑YO&����2.\�&�7� �o�C�L�6����8���o���?�|��m�ݶ|�r�2�Ͷm��mL�6D8w�ܔ���W0*����b�g��Ő���'�4�Y����_��"��?���H��;��>�y�6��Yg���q��q8�� �#�C�b}>nroT��p��w_Ok���<
/���Jx�I
b2����SN9塿?.)P�j[{[  �(柄aG8ݜT���1M�������-?�Vcƌ�2z�8�r���;�w���7�g: ���d��qAsc���:TU��#�<������|�鏤�[��Tol�L��Ϗ1�}��u���,n.���G��] �O}VZ�|�葧�~������W?X�$~ue�Pw� ��/��w���㧖���p��4`l��"�.��[ZZ&7����Z���o����={g͚�c�@۩����ͱx���X�m{�z�u��v��2����&O�gA����}����{<��a�y%����BV������?��>|D,���b^%���0���?��d�vh����|��}���sA��ļ|i��`�bl6��2��U*mj�����Λ?_�m�M�[E���j
,����C�u��M�8{]Z�Yx�n'V������o_�dɘ	��z&L�)��`͵
����^�Jw3U��>�l����������$`�	�r�v�9�c`X�33�ÇA-�1��E�-3�8x�;�m�{$fEh*�{N�� �A�IIIN4ݹk+d H3��E�T�UĢ��	Wb��n����W̪�'@����f��A��`g�Q�vd������4���Q�tg R�_������]�T��kp�֟��P�񨁛��?_�΁Ue���)�g�/T��<|���������㏯4��ä'<�d,�������^'k�j�I*��Lmr���-(H.Q0K�?[P����P��n��qxֆ�?��4p�cҒ*ur'h:��5�� '�*'����j%���}6b��]�w<����~w��n7sDb<��ժV��*R�j,N��~�D�n/�O���D��>oQI)�bf�7�}��ҋ5TNIŭ�ÝT4r$���+��(����ZZ;X"�T^s��͋�1�<�ӏ>�����4AJmo��`и�z��h��h}�M��u��ʁE��\��wk?����YM1(����S�E�X��j����c�Z�&�^؀�h�'�RR8g�H$�mt�^VV:s��mݭ˟���Ƥ�]JWI%"0e��7��\9Nj� �R��kS�^:����xɏ>�0|߫��3��i���lԕ�P)���d����������?_y����_X��'ȝD<������ @'�����`Ρ�V�W��=�4�7)+-�?|�<l��_L�P�L"I�ܑlz����� ��}���7A�_t�E��6�GF��Nf����A��O������Z�>}���^#��h���]�9��r�3b���r�(�)XҟS(�]��i)��\�{���V���K��[H� �N��c#XN+k�;�6B	Z;���?��5~��3O�;�=t�������M�����eU�I)����)-��`���g��"�EG�y&�v����?W�����Ai��Z����<N-����'���[߬����o�:}�Q�q��-�ޡUUuuu`��C�����`�ij��z�M�y��U?�����/���uӦM�e�bp��)5ij��x���O�=ɴ���
=�b�d1k��T��)�su�5JJ�vm�p�m7�w9�O��uw���%z��/���g���-�[�:�h���Pd��+	���*�����vˢ��8�y/<�,��^N�+��66����ܵk��b�9s��U�"�ܱ�����O����F2���;f䠒�B:�J�x��>��Jc���x(M�8���i�)s/���+����,��������w͘:���	l��B��$��������q�����?�[����bT�Ue�d�`Ҵt�:s�A|a�htt{�����c�&N�[�b�w��vt����(��D�3Z_cccoo7,�I�FP�Iy�Z?��㺃� �&�L�l7���;��u�Y�ܲD2^첹l����G|�`h��Z�F�0�F#%�l�6tPe��I��3��O?�j�'����yT��ģq��Y�$�\}~X��N�=�����\W]u��'�U�Cu�$�4f���j�bi�T0�����M�1�#ؿ���6N?n���3`=��<p���ϗ�;kw����z�h�_P�v��ᄵ���gdq�É&!��Rj������^
lb.��<�L�>��Bif���|6��h�@�	�k�~(�3��������3>��@�s9�1�a�`�)S��������X�� dxEk�X�/vD�L�G)]� p>�!���Z�v���&�FU���E�ǇB����V	��[�ޏ�']y������
�!�]�(��O?m�%TUUF��!N�If*%m�h9#�j�;��b��3!wT��شi,D�wpXO�{"++���{f�F#M���b6���`�Mq�A�eeEYo���|:	?�����E)�#�Ҋ��(��o���d�j�� �A�Nh\��<��3�;�wH�W]z�n�s�W��T��f��b2�2W�i���ttv`�F�~�����5,���^�ڱ&�}����@�v��[IR��A�C�_�1��N�y0#c����zx��.0��L;0�ͦ��).��Ꞟ�(S��V���d�YQ��R�fNI��#������p��l��r�:r�H$U��GV�~�	��@�c�)g��m��/�_l��-ð���^P�����Q������׿�����eI�Ќ����{3���k˶���#�m�	���{>4�3�|~��%앢\�x4�O���q����x`���g�}�ĉ�i/d��h$@"�61�G���b�[�m<�Dכּ���7߀���oP��냹	��O1�>�W��|n�+x�@L*����z�I�m0���¼ˈO8P����}�2��0T�Ơ��@Z�P5�Z9�F8R����)ӧ�س矯�|�WUW�A������Uw�gbGr
I�twtP�e0��4�I�V�FHZ�ЊҲf� �a�Ν+^|��wߝ0v�G1�Dz�G�����Z�lٺ�[�t�Ě�#%%9ssag@`���Õ�`n���S�m����=��Sv�\�pZw�����;�i7�v���'`U�[Z�[��EM�zz���j�wQ29���l���ͷ��s�MTy$p;8p����Y�V�\�f͚�n��SN)()�\��۰쐁�C�(�*�Vv��a�菟9��9_>v�}�V�7m�4�#��O7�E�[�X�z��q5ؠܼ
���H]���"$��S&1>�
�`O^N^n^4X�~�O�a%���f�WII)hx�:��s�b�{��x!�����\��7!^��XXø�es�v�I3V�X�	Ξ=��Ql��
�Ԝ<��7�����=��Z�Y�B1Q�3.���bv96����z��n:��Sՠ��p|��S���>�xݽ��;f��ѣGnhھ}{�3��+�B� N<|�o�"O�Z�P�SEFCm��!��eќ��隔߀�j�s�n����*E�9�ʁ3���>��������E�x1�
�������2�Ʒ�)�g�d��(Ym��� w��\*nTRO����T�B&�,��,,Q!3d�(����v�UUQ0�5�z��1���t��ܶ�f(K�˔IS��������R�kY)!�����:	��h��a�ΠS(�OS��*Y$iE��Gd��r�n�q/iDEK�|}Ԡ�l$��o����.Y�^݄	sr����5C��P<:��2��q��B�QM� ���>�ꩧ�ػ��A�$��</����S�t���w��ȯ��@�J�69�\�I$#n÷��<���>��o.����C^�ծ3�E�׸��`^�.��{���V�Q�nwO'6�vРA��7l���C�|��'��!��$�<�"^B²�P8A�ꉤ�ˁH"�Ft!���'�ޤ7P�^���j�DmV�����n�i=l�I5�@nqh�ޒ�=��3�l2VV����H8�G��s�\���(��י̶�*�9�$2ž���x�Yg�A4�rC��Q�X_�jdN^�;�3��7)ɪ&��8�KQ��?~�G�_W^y%נCN��`C�XF�C����U��'NO:��b�c� ���!�0n�2n�|߽���[�fL�y	�_1�>�J�2��6��]�dv����[�����-8}	�k~I1nX��\̮��K��䑖G~�̪S�[Z�����<�Ȳ�$�M���^.���8z����:>�9���6��%EŐ�Z��H����~��ATTVҐ��&�8�A���M�#�]�����#���}���s�.��8�U\������S��!_��C�Jo^��{���/��.���^��ŋ�|���)㵹��`?J��Ap�X���e��Qcaq{���=�$�A�E��$�[�/�V���RRҨ�T��c7X�r��w��uڢ%�S�*�(G�D�%%���������=UuÆM.�cjM��_�����w������҈��x�s�9;W�ԐQN�=v������p�QNqa~.��M?x`9���׽��k׮�ˣ:C�*�t�0:2�����i�u���M�_1{�l��������ø`���8�w�R�A ��_u���u�o9���7����W���������6+���:V�0���_z���+s�P�(cK��a��t�j4�:���nwo������p�s���g�~�2�{Z����8Hz��fJ�tY�U�~i��k�qޤI��J᪹��S��inm)�:5ڴ��$[:wS�P�㼋��4yγ�>��#�X��g�<x���:7��������6o�qNe�S]]�Ѭh��p�������MV�E��A�AP����
�T�3�*9VPB��+�_P�ǋ�?���Sw[,9��u���U�.۞�4J���ݶm��`�����E�
���i�Xґc��������ƍ�p��c	s4��K��"�ѴI����g�1v�$�D���nv���o��٦�`fe3/0^mm-�s�=7��8`Ȑ��XM�p���تʸ��:I�Jq?��f�|7/�|��m"��%�W��-d4��8���5�eݢ����\�ުGyd��ZD��M����	�����v��RBJ�dP��F?��kF4V!$E�x����BL�W^�ꫯ.���?��6����i�aJ�L%1�]�waA����``��-��y?���׼y�pOHy6��l�#l�e
������_�6M����%"PH&P��c�=���kaN����Tx)s��&�V�]�.��2S��
N��ϠA�1��n���WW��0}�)�%L��w�`2i"X�p4��tAs�F:�,-)��v�G�L-���|��9�v�g��XВ$J`�?X���\X'��{z�-ad¸?`��O(��X\T���z�]w��	����J��s8����K`��0��'>��2r�(,�|P,$��`�X��.\(�s5��� �:���m�{�?DM<%	�1�?6�������pk`awwV4�?q��p����~�2�&|qQ��cw�L=\V^��� n���%g����3�>�Z�ͦ�&c���Y�1괝]�E�ԏ���F��^0�A�',6���T)7wԨQl�s���~���d��&����DR>���̗��c��s�=���jBM�3/ϙ����q��l&���ܪ��\��SO��
V���v�R59�P>�$|���^������^��C{��VՃQ=}[��h!(�T���z�i�y��V�Z�����܋˫�v�A:�2R�BG;y��t��{G�V�T]5i��n�a�òQ���u��[�B�7�*s�2(�\TX$K���x�E<���7@$�i�~���5������k�nݺ�?��*���e��!�Xr߾})U�h��m�a�	�?y�֭�ZUy�V���ǯ}�э7R6��q���?�Ϡ��?�;hn�����@f�� \YZZ<d�X�]=]+V<���{�r*	�F���LhR"��Z���+�x��/��t��l���{O�e�<7��U�gaA@ؘ5Vl��	/��ښ���	tˍ׃A�/_>z�DU��ٷ��`w��>^o3����J��9��#G�� wkk����3�N ZQ���_��Łz&���ȟ����K/>���O�w��3w�ٵO�^:��R5� )^�/?		�����G=٣.��j? G�]�l�c�}JK��� �{�Q�G��������v����_T��[��9
�i˖-'N�J�����y��x:��*9=>oCsSR����H%u��D��IQ�"�>�If��0�xB�0�
+A��G�T�F���t��n�Zmnh�򪫲���b�9EMz�ڏ��zݷ�|We��ɹ���Z���V)ũ8�%�
'S	���D�ؙ�#AY��pwR�3M@�DD��I`'��&��WՀJP���~��ꛯ�a�ԩX.^J^UE�=��'~���O=WSs�����W8��Լ,z,r��%�C.�%��ǚ��՟eOqf#<�P8�Hr��F����c2G���T���.>c�W\�V�A�F5q�����D�d6i�	�	7�z�B���3��jn��6�Ͷ��|X��<Bq7�	�B@4���r<* ���DRG �c�'�&�Y��%# J�����&B����;��y����b���߭[x��g�s��X��a�F����t�&`6��z]w����L�")�:f�x�������曐�cƎ�*r2�?���A��<J��Z%
F�.N��u��g���������u�RA����{�g@�C�G�
����aX`M�Lp�
��F���B�	����i��W`���I�lbQJ��>i�,�L�L�,3��G�ؒA�[IIĕF��ra^��a��~��v���� M�^��I��p �F-6kWO����7P_+�n_Wg��Ӏ�[�^?tpUeV�aw��o�6���1l��HUv�IJ��<�%���JMaS�Z��#A"B��j���&�8��P8��,)-Z��7������r�䕗J
����aSR�d�q��Ba�NW%Ȅ��ҭ[)}���8����	�0�,&�p%n���Y���7_n(*��L��vw�B��9�pPk�'�є��A_�0Pe¨�S��U��P�ڵ�]�`��sοpҤ�r�v�ЋI�kF.�\OX�}�m۶���i�ŒjsK�b�;����zE$5)����%Ų������'JOOkue�eH1�0��:$J%���KH���=�B���E���O/{���|���g�=jXCS7����(�������f1�b��J��h�ݸՌ�_~��5} ��{�IX�={�:t����b�Ut��ή��p���-����c)VgԆ��w�~�?��O4�;��1N����a@V=�)�H����B�C&������R߯[�����\r�i���S�{i��֮N����"�W���e�>�n��ӗ����^~u�ڵ��8��?����{w7�@
�VU��y��Q�8xh��a��zK�)�<��;��㐌�p<������"�0��
T�e���p"��K���&L����9r��	;v�p��D-e�� 6CT�p8��P0)ЖK|�Ȅ��n�#���c���8�d�;��wX&�-��sk�G�QXZ*����/�>�^�>7�}ʁ��1�;vp{Aili�t�d��g�=�8�tCY��$��M��%F(d,3���A~Vi�$�[���B��k�����χ��D�E�a*:k�԰@k֬�p͇��<�/�����X�ʫ���0?��R�.}~ϱ���2��cQ�R�%m'�
"ѯHGb:h��v2`�ß����	;�R��Syy9H��;�u�e���C��E@ٱ �/�r����%���?ge�i@��of(>O��A�!.:���x�-��<g���F]�D�*<�B��D��*r����O>��>����UTVb���Y�5Ɯ��:e$�U�,�����H��\NJz���l0R��(��e��Cd������o�|��K@>�N�����]�T��ki���q��JHS�^u���޵���8E&,��^тz�ÁU�����L��`�R�f�>�y�七g������
Y����)S %!/����O?��of�a�̙��5�Qlkww'd+\���PWW��C�u%Q`��<���9Λڀ)�=yŒJ��� ��j%\m5�tww;�(+6V@K]�����?��`�je��D}�}\#$�M��Ô�%�D���-���5E���H���?��O$�0k|���EF+#8���ŖÁ4>Qf�I���ܗ�̩u�He��q���v'��[��Y�_������9Ҁ������X(*�3�9#�萍$xo���A�6w��z��w���в55cp16�2l�::W2|I	��8�������M��Z�T�`�;�k��SO=�K/�_Y��y!���T���{��JH옦*b���	+`a'LgРAe�Kv؋/�!�X���奎�j��2A�![˸j�i�OpZ�XXPH��s����x��e���wߘ�5�4�v566��
9�O���9r�~����3��7o�U�B��>���%괚�Q�������;шj�b@�=�3f�V��	 /փUM���X�D9����v�ZìY�z<*�އk����3炝񠚚�};�0���z��G���a�4hh�3�SN9eѢER*�����Vy��0Cb��Ņ��Q�_�DP�0p7WU��0ws��h��t��j0R��k�u�=�D��▿�5v�X�/��TS��B:t(�C�~�'�!��St1�&%���I������3�cT3W�����L��`er���b�nͼ����i�i��"p	J/��A��������ϗ����;���6G���L�� ��˱��I�� �*��xWg2�BP�/0�&�	U2hd%.���kD":���.�s�BVJ��O�5cHɄ������c�8p����M�6UR�������	ءaY�<�x��O��t&S S�
D!�I)8��f4N��(ʞZFj�F�PI$���֥J�'i�j�*���~$�&�EStʡ*:U�$�ɐ����Eg;�y������KJJ��u��A���t�g�N�ޟr���`���]�ׁ��T�$լ���Ԓ"�'�Yz�>�0fی�XRt\%4u�֤�t��6k*J�	A{3VB"J��&{u��{��s/?��Ӕ�$�rL#%����$3k����ږ-[ �Xg�C��;$�:�S{���ҒT�h�1уG�
)�X��[�pFC^q�J�։�&�j�^"������3;�������b�]w�u�g�]�Ū�(���V��]���ܱ��yK��?m�}��G?��C���añ��?S�Y��!eI��x���meuw>x��@�Q��rV��a+�Q^����	E�c��:R�<u�ࡓ�λ�⋗.]
����޸aCUUU���+0�Q�3@�r9�	�&o¼�僓���q�;!���hXP�.�0&�I���x���i�+	���f�uĤ� ��TܭM�z�Q+�0��X��$���o?|�0���Ao�P/�X��0z��{�vL[OM�<H���-����)�\���;�}�������%k�>�a5�t�T���=�`?A>fTj*���1a�kRD�v	(o1賙š�ӭQ#r*��v�}�	c�c�Xz�;s��|˭�M+γϪ��S���;v$IL���̉F<�-��m��v�*$����v,���I�����?������a��┼l2���W�x̐㌉��uT_�jt�xJCF�A"@P�?ѫ�}��UYVOD��d���_-Y�dѢ���\���0ޗɢ��x;;Aڔ����:�}��e�d�[M_���JA��X��pQ���0���ڄ|��KO=��դ�5�'�y��dĦK)��R<	�����UX�q�	z"b7�%l�A�&5�/uG�6�����̜�4VY��o)l�p�����AU�ruKa�ϧ�^j��q��/-�ApB�X�_Q68
�uuB�:�8�B��n{��/���2qp�јJ(-L�$���\~���Ɯ�Da)��&�v䐁�5?}o��o�}�I'���9��ۿgϼ����J$�&�����M�D2���ǌ�R�rZ�U)���)����M)�v��,.��o�����ʩ,0´��>�&�H�Rc4>��+Ce�R8�5�}I�%��9J�����f����`�?����64v%��7�h�j_��e�l2�-��r8����O?�J��ۜ�a@�Q��}�$��^��z-�\��|�����7�ᩧ-Ԧ��I�K��f�9Kg�6>M�"��6e�B�%e	2�<�_'e�d��X�%Q�G�"�#�?�9��0��O�]��-�J�<��������g��CU	S��W�ejV��� �/g F7h�����IQ�g���U�)���G����;d���U>��CS�P�NeG\2�`I>Z��}:��+W����m�˻�d!����=a��C�[n��_<f�~�b�a�H2��|���% ���V_���\����zΓ8����w�������g�]���C�9�&>3�l���r�	&+��;��í8I�7(;w��u��~Y�D�����\�z��U��/_�fڴ-?��!6hڴi�6m�69�����{�b�q%U:�W?f���q4�#���*1Q�i��a@p�L��"�%�nK��(\��/�=z֬S�f��Q��.�~aF��v��f�w҉���n����k�2N%���sx����I=ab�	�`�l �$S�=��a��N,&�F�ak^z�3g�������.���ˏ�5�t8d��A�LN$�8�����NX~���k�?&B�����Ͽb i"<�դ2ؿxA���R������S%^��y���ỳ�>�f��F�%��(��&k,��-�X__/�(��T-�w�n��̠���\<��o>z�'Z�O�81����!��jFv?�F�Q�ͤF1=dK�gAx��0.A�?o�7{���[z�7#4n��`xS���TQ<����k/(2r�$�Q���g�fFjI)����#U�cp�e�N�Z�H�J������n.;9r$
���v�i���a#G�����0�a�Q��A���B��5 H)z���1�Ǹq�}\J&�^����F&y�hR�Og��l���2o0Gl%���ɳ�~�훯���o.**�8p�O[��ܐ�Sը�p��$�xzzz��p�����a8����E�a�$6!�8LJ�w�a�?��#�~�&q� [��/�~f�>m �����mx�Q!o�1HV���-+�~!�g���t�*I���dr	In�T�K��p�)n�D�F�����چ���)g�nL�^&��;s� I�1�\Mc�����W�M����QJ�Ih�����1��>0�q��g��!���(�뗕��������ߌ�AnQӰR��0�ͯ+��j�0Dkkk������% 5�^4�r�����d�G��\�E~"[�� X�eV������ݻwo����~��2**�����������^��C�E��T���e�&�6��D:q�������Ϯ����3����\Q/�]��+p4�\���׿���p,�Zx�u���_}ݺu�|�n��(�t�-����+H&{V����,$r�"�X��r�VY����S�0���"��b_,^�PkKǔ)S�'L�;E�m�;��MRO<�Į��1_�~�f��b+)�U��ދ�B���E����j$J����%
K�*�P0QMe�z�xC^��h�ҩ���q)���}���N�:�w�4ǙKj��PX ���K�����46ٱc�9g�UH�M�W_|��+����ۨ1��D��tg^��~�.���_�}�J�$P7�����в%E5
v���/U��a�5,mm]<��)ϝ;wܤIz�n� aE!��--����6��P	͚�G���@�[�|�=q�L��d�S܎s�Hf��?cA+�&�9�<��Ex�,��>_�V3u"�t����[~�mw]x�ƌ��X��'�ް�`�nm4)�v[����'-f}ey�NIi���NŨÆW�ޮ�w�y���A���.s��\���_�R��|M�̴����8���T�Å���˖�}ܔ.��,�GTw���F�h��b�b)���u���9�ݻ{o��Rn��
˫ǂ#�=͛7{������TJ6�Ai�h4�IU��f�ϯ�4#KKR#��+�������ut��{n�3���k��:�*t6lܼ{�6��Z��+�:��a�	{
�����K�UK7�Jeoۓ	V�|F@���>R�W^��{�f�������7�Z��J�2x{{���?��̼�|3�=U3�%��S����hGV�!M:I�@@E�#^��  �<:�#�9�ե8;T �R�g�үrs��I9��Yg<3n��fʯ�ƹ�w|a?E3Z��}�P��Q"�ҽ�ak`��1����ZU��;��և��V��WָB�pf�����|�����e��W\����ŏ>&�s̋��3>z:{Q�Е/�-�X�P:0S���,;T>| ���xay �H/��������3v�p�I��_�/�z���;�l�>���5֍JL&��T8���w܁ń��\w*/�[|C�%��2<�o 2rS@	���^"�� �~�]�&Ì�!������wߥ���������0��n�
ɖ-[����|tك�}���q#����z�-zJ	}Æ�&3��8�"� ��g?2	�\��;��:#%���V�)Wö�l\�z��o���%@�<DY�6;iPj�.Z�_~���[o�����(�ڮ�>}����z����IIG����}6�R�f��XmA6��u�D@?Xa,V��O?��Z3}ڂ
�J-k��&d".�\�8�	ӌ�l6���=���~�f����&��NJ|r/^�_�F� �r�f�����J��̺�<q���;��W_����k����	أ����#�iZnW�gU͍1�D2���Gm�П�j�T����(/�ʒ�S����z()K̲��'r�ދ޵6o�6q��L����x:�<�ng^!��+����rS������mI|I,��0ǃI�E)_G�k��Ǩ�c��|�X�RC4:ۢE��{C�ӟ�yu������w��GL���4�)H.>g�r�GG8�$	@OQ.�&K����!͕Ҫ��"r-�h1m����yn"Ѻ߽�4{Q��]>A�"M�bI*PR*�Lx�}��f�DZ�o���$aO'ɾ��4��nÉ7�+Y��&��A�i郀P8����v9})SP���M��g�]B��󃠹c�-{G��1������ȑ�_���P?����K��L*ef���"ي6y�~e�a��Z�_�ʉ�qfnΡZV�	��Q�rr\!ǀ�� �o�������:���D#�_�X1�"��I ���Ҙ���'��`����� ��b�C:Xm:~:+�~e��q��Y�Rl\�h�#1��鍊VOm�0�_�a��N��[:�N�!�aϾ��jnm!Q�Í)3�L~�uu5c�T�����t��A��*mL��M��q�`�׫)k$���h�A
{����@�j����;Ml������z�n��[55��r�4�r��׷��8(:�������"�y=��,����\ԤFp8���yh���JRWvV_�6��h����H'�:��Ы1�u �ը���f�W�ۋ
�W��ݛC��<W�9s����t`�l��B9wUU9qݟ/���-�Tu�KQ��:��bI&R��W����3��iP����LP�L	�񔨥&�+�๋C%�DMVl��K]^���x�_�����N�>((ty�z*e�S�~"�5j��j\����?;a�����L�zE�/�ǡD}�^��+�͌�#%�ʰ�?U4z��К�԰$��y`^|�BP�E��?�S�r�]�R��
V,����).%��Z�Fy��! ���|��w��h�Kɟ�Gz�=QYK���C44
 �!�S��>�a�	n��l����F��
S	����1��������ӗ�-<��z�͢U����:�����ʵ[R�N��0�0a���ej,���K�^���鴘��y{0@(&�"��8(8�8H��|4��F�q�wwt�avp�s��q*HQ�`=Q��/�蓯�}�z�%W�?a���?m���@�C1�z�M�KJ����`Y���l��=۟�J�_�Y/į�
�d*ڄ�����N�����;�g����@"Z��K�!LA�q|߂�P\X�F01�/����/�wT>�d�B>F�g�HZ�z���ys��p}*�����üu)�Z�&����0�� ���ؗ��|��?�ѱ�>ۘ��I9�bJ��(�1���g�c����g�ɂ=���~# T,x&#� ��yF��/�7��%��UĶ$���6
�3p������/md�6�21ꌓ��>3���HXg�"�*1� ��g^�����MP43�������o󇙓)`��fX�3L$KՌ��h}#��5��.�a��2jDD7,,��7e�>D"�4.�"f��.f��Q��&�'�r�Ce�5Bqjl��`�����,h��_/�������j$�FA�h���ᦦ�ʪR��S��ʶ~��V<�1?%��)U������b.fR��'��r�μ@یGD�0݄��RL��m۶��`��A.8�#�8�C>�/{�J32d�A�A&"���BVT".�oRr����<�,���u��iY$��IώOR8D�V��V�À߳~����A"O����mh�`z��a�˙��y≇���f=���T"E�p���ԔzT����,9���a\�=��C�b�x1�����!��Χ�v���g�}�9���A0l}����@sO�����w�5��H%(��ũnB�b�g7]J�93����1�� L{܊�8U�;Wa�y�ѣG�~��55�~X���`�8�
-H�<JJ�#�7o>th?�[P@�� 	\���*�0%���t�%��8�o��zs����*�I��d�̝;�������n�m
���1��{Ϟ=�`ϛ��Lr�����VJZO jIB�1JF�I)Zd�ꇬ?j�o(=�d�����ÿ�?�%z%�ك{;��`��}�������b�'SP��E&�j*���OVe�%#	W?&�!TUƟ����b��2�e̹����������,����}Α(<���w�r��>F{�O�?�,2��/A�)NO��TU�m[d��h�!o�=9�u�,�Q��럹C�R�+�HL�C��, Q�N�|�[\-�,����gް3M&d���Z��כ>zg������oH���Gf����/��3	x�����,B�F)�M�o1H��
�`o昀+�y%3�'|0ĔsTڊ�r�1�RKY�TƗbS����;q�h�C[L�#����x�C�$a1���|�������jEu���@�fl�� >��@$J����HB����F��[:R�&٠3*�^֛��E�P >��b08���;���>�hq���]��5�-}^�$C����,i2[����n����r��z�����/�`�$X�;�T�CwrJ0)t��%ˁ,fC0@�f�#@Г�Q]�/(��iRe�Ũ�?| ��:+(rm��RoW� {6��:*�]
�s�7�i�8ĺ&%��T��kC��D�A_��I�_>V?iu"4%�$�ɱ|�xa��Q�P�#M�CQBp�����UV'�����L�9�a�@VWwG,1|X�o�5b�Q���&
�G#qYIB��C~��r��\��
�J���\:�~:�%�`��#C����WaAѨ�b���ʋ����ү׾��K.�2qt{ ��)loi��W�ђ�|��X�Ƚ*\�]١ӠM��)���o�N2�e\�lG���!��f#�����P h�h�S�o���2蔑�+j���u�֧�/�6u�ڵkUI����-M��E�o��V2�n��S�>Z=MBJ�4j��LheIg&�M�ZlDU�/T������(�3X,�@��8u=����k���}�is`�Θ>c�Gkv��	[�=�fR�A�\S���R���;>nww4�߯�n��݌�[�	;�LѲ���W�A��V�����6ؚO�8��C�%T"	� ^נ꼌�ɑ���K�ݐ9�R�l5ۢ�;�n	ܞeR�</G��U����/���<[�g=�7ռ�?���_:�\���3�"{Wr�|!�%�𵔦#D������&��]U��\���>��S}����H�&mPi��%AC/���@�{�S����\D@y��pC�>�TU*դ�S��N��ս����s�}*(���d�]��k�1G?�Qb���4�/%V�=N���l&J��l���9�V9��4��îf�֥>�t�y��X��تG�t����̞��"G�Ɉ?A�O"8�`	G�HҩO0	��S�e� �qF�P:t%	5Fe����1z����2�Ab�58�_b0�(�R� PU� �� �V\�X@���g�)6{H����{g��#:��V�z��u���*I���'v���s��1�%�rO9v%R^O�!E��ZZo'j]J�S�Ѵ���a{P@7$�`�,G��hf~��7��ɺK�	�e˖-rc�l�+�c�ĖtCY,��R����]��3�'YV<�	F��+螁K~��ƹ���90=͆����}�K`XZ"�' H�|���]�nux��!.�֤̩VO�Q��0�2��MG�Rh�&�^m`��{ga�����k�i�����{����N+ھ}�b0���M�e\s��k�5�9�x>�j�'-�oF�4R�|�j�N�8���b�+��L���;w�qף�v;_��/����y�E��q�F�U��Z-�6�"�γ���%����'K�k=,�W=0*��m�M16�}�lW��8�I����=�|�;������?���n/`f�qX8M�'��1l�7=����U]�D���  {('�ti#Iގ0�E��+�G��ag�'��@S�<�{~�q������׭���:���=�����N#
[8��F,0>u�e:���n!︎���_���zܦJ(�<̒�O�-�֙WZ\l--Q ��UӶ�r<^d��jʙ}����i�.5�_Z+v�H%�@�K�!��2x	��T�&�m{�Ѡ��1�&k?����y�a��A��)NK8�z�d;�?��%�-���MÅj2$��r��7�J,�C�1����P�G��X�X��M�cr���"��#w��	�0+b���}1q����Ԕv��#��|�X>K���⁔1k�p��Q�-��K \����1�d4��a��x�e�e��D�$m�'x"fOJw��Ru#�+�dVAOB��aa�ź��2ݙ��r>������I>�����
r.�}�C7,�^~7�M�ךd�������i�����;��Ն~4�efl��-��a.�\����[ȹP[m�jKb�E'���1��8>WK�	N����O���vq�@YD1�]��'QL��Ё�:ԩ��i#�S7�犅�8K�@3��}0"�:�*&^B�8q��]�$�,Kqa�$'u�Z+�d��N8��Y�8OȘĄ;�:��ϔ�nm�D��ŜG��%RSS�.E\"0Q�.h#G�e��r�©P@9����n������޵R��Vgo"�
�r���x��~H�~��(�z����a� #$,WF��Ջ^��'N.�9~饗,����i�'5J��\�n-�re����@:�{{k�1�#:�RF�%�aLN>HҸ�х�٨U�+K�������w�.x|�.�e�ZZX��h����罀6�u� !�]�NN�n�m:p�^��=� �uY�z�e���][��J�F�R^���J��ӳ�wl^�M��]�}!�	b�;Y�D��A���2u����d!�m!X[м���⊫���߼���3�R&��m}s8N/J$NV��������x
�-,Â��W�E����+D��st{AE=I;t9ۗӪ�Y޷oiCő-�sB�c�l�]NFi
���糩�6�)Z�K�wčME��g2Q�~������g�]�o�|�vAO1Ø��o?μ�Y���91@��m�ڑn2*��c�i/XS0S�&^�4��с��Ǐ�")"��@˥[��KYaC�R��V3�����ka���=[G��0npO�'��lc�0�dff�|7�]+�c�M̟Ƌ`�[͗2���d���ZQ�y'V2� (� |^A�ǁ�#yr[?lѦ��R��R3Z�l,�\i�'�R��ZC�}F�'v%K*����;��&us�|���6�U�t�����Qv�Y�/��jHj9�z�=4��U{�X�L�/2�7�����3�$�"��d�
�C����k�M��$�?�4��K��U��(�Gl6r�#�7���V�#>�!'S�?�C�%2=�pU�4/=�sW����<�q��[R�J�TbH��������C�΁/�ס�<$�Ͽ%�/��$[b'���(�r\1u�J(��� pV�n�����{����+���C�<��~����!A`��{L@B�[ik֬�ԯ7�������3�a�I��ǔ�G,S%�o�D�)e6C�)�WT�8�܌��'�;�O�M5�aeάټnݺ�B�Z{�o����H�=�6L�2��B�(�~�=��i�P�A�#�a�PVe���-ƽ�0�T2�e8�C�@����>!�ɢ����s��F���U|�"��'a�c�!��R���L��&3ڒ}7s��T�p1�@���L�.�������<s+����r�R�JIf<��f���Ӯ��I�H*��"��)_F��r3#��y��T�L��D\%W(�u�#i y5�Gss��}��T��z8g/���l8��n���fq��~frbb��/�Og*��	Z�KR/�zԖ�#�)����?�!�@۰�
�IF"o��a��:��'iu�eiwx�P̛�؇��\��B�V�ԅB�%��$L�N�9	��nBj7�	�ʸ�&�`�@v�R5D�:1�O�?s��a�*�1RVlz��+�cx�n�u8nA.XԺ�8W(�YXbd�B��)͍�U��nr�ވi'����X]����:��UN�f���	���.!����&���0d��G�T�I/_7=�栫��#��JKr���������<�(��#��
n�n��8��#�	�&���b�󻡃��e/�J�r�Z�t����t(��GR�X���H���L��Z͢`�6+�YO=���P�������	 �t;�\���!`�/خ��=U.�C8Y��������C�޶��bu���}�W���0���g���lV�<[� �$|nwV�^��.�kZb]Pq���e��.1n�T�1�ᩤ.�@.EG�V�Y!<�IO�/2�+fM��c.�kކ&0�UG+M��/�8g���'zY��hH����}V=��1 �M<���̒+�!0��uL�ll�c���aآBi% ���(�o�k� �l��΢)�oaIue9�ʠ.�,�������PQ�I����7 J�}Zo[R�XV��յ'�X�7����l�GY��p�Ĝc�S�38��L�A��"����O��?�jhM��7R����I�U϶��3W�JCR_��2���%��$b��$kG�	�6*�˳���*�MR������%�ĉ�*22&���_Jx��퐍�Ϸ�>G�x�˙� ]�E{���Kk㈫�ċ ��k:��W��k���4ߤxR� X�"�4[�f�?��;d�����*�MEi�S����,��ik�9e[��X���D��=H��S�#"�	�/K��\ϒҢ��2�۞�aA�ZXY6�a_�o����'&&��YA�0ʾ<��c\���t�ܟ�U�;��	/q���z6 1�M�a@�dψ�S<��v�9D(�.���|	�J:��O�K��V��g�g����`�6V-KI���B���EXc pvA������5pY���'t$*G%aS-�*��%�щx
�v_ٲe�������'��+b�WzLJVȸMt7��$�)|>�u.`�sss6l���kz�!܄��u�bYΑ�U�'pB��n�]�U�>�)�F�=B�Z�
��s����0*�T�= #�������/�L逺�ͅ��,ee]j�!���⸶y�/�m梬���H{1�Hpk`f�7I�O&�̀k�m��r,�E��$�n�]��1��e�y�3EPK�w!�/Q1UB�����J��c"�C"[����)��^�&�a��Dg>�ԧ]��Fs�(q��� $}lإJ~r$�=r�����O��?�O�� �\"�h;�n��{4̤������� j7t�4$�QLJCCb����z� �HJt]8(%�$mQ������qɬ�z`y_�����ɏ���X�l�F�ӂ���z~7^�=��)����n��N�S��d�	 ߁6��i�@�H�AOq���T"�"'��MF���.�����+1�I�"/��(��lV*du�,�~z�y��T"� ���UK��Fk��k�٬���#��r$�]�a$n̳�SN*������b���dVf����xp�Ӄ`&Ow��ސQ���O2X�hm�c]8W)�c�h6����z�4	�x]�6UU��K�Q�r>�}&�閱�����5�<�l?9om�p2e�O1��P���^G���f��hu(K3���"�ž�fC��b���N�����0� @��&��Q��W����?p����c6%��sI}��  $7#�tDI����0<% C�Ҵ�����g�fb��wi.Za�I�v�Tţ+剽{�R�C�<K�����F�I�ф�����"q`(K���z6g��x/�yw0�,�R7��s��d_������7Ұ�j��>g�*s�њ�_S�����*	�p6M�6rt��Sd&d`����F��N��VC-4�,K)O�4h�y����FTVP?��贌)G�aͨ�OH� �=(;���y�,��x`��o�ʬ��$m3�H�ƿb
"V;V����m�6�;�p�LF�Ȼ�S�|O�ZZZ�d�C���ׯ'��n7�G��X�eS
�H
K��$�ՄN|���O�'-줰($�Gvk(�1Z�.﯄q�ދɘC�\v��̰��B'4���gb`��pހ�bJf˝����&���l��a�ֿ�f���Y�B'?칅���ߌ��Y�}��&`�I��,�<�"���6���|C�>wp�\+���+w)S]09$-?�j�!��b?��M����j��6����rkba�2T��+8I7��P0�x�م��w��P���h^D�Ji�5A���3%9ʱ�����1�ɽ�iKҘ 
��b������ܱ	`��)!��D�.�!&��s�=u� ��?�O��kpamo~���@�j5��ߢ�(�B���-�3�#;P	P�*~]�w��8(�?���W�v�:6�Y��wI�b�3F�o�%�i$V�TX���m�����A��җ���
yI���L��14$����U=�i�C��(.5-3��^���l����&q5��϶�`���F*��r�ַu�Uw��?�υ�
�!]�A?R!��3i��m�ꩴ<�w�a����^�{G�������"�S�oo��lN#G�[)V��ɷ���* ��j����崯vh����?^f�<䮓�O칉O�3��P��?a�s�9Yy0��f�~��y��))�1RX-#5����R'S����kX�c�����ǃ(I���s�L'i��f�n;A��f`�V�q��{���]#�U�=�1��=w8%RAMT��s��.^��xy_d�Qg<��|�ܨ��d=3)@�`U�#���唗���tߣf����z�r�i���w�k��ɣ�c���'����!�Gҗ�I4��N����1Cb��L�e�H��|f&ɡi�?�\Zkw,|k���H�o&��9�/�J}��j��\����)���;2&9y�${��<����Rڹnڋa�b�\���>��AY�+�?.��J7 �G�ġ�m����������X���r}�� e2q&��jF»$�`9^漍t�|m�i�����.R�ZJb�����Y�S\lt��]=IAFϥ���(}x�;��Oɔo�{����QW�G��:�?W��`j5�'TR�+!�H���\�}�LY�gMS%�	Z�Jv�'�����D�9v ;G���4l�;�����h��E(���Ҋ[j�D�I8{��jWS<����j����ɑ��U�42'b� eޒD��I3f��B���B�?�!.�{�J!6��ѰP�)����^s�}�U������^u�U�v��c�8�N�Ji��u�D�=�,��neL[�%��PY#�����F&�i���ڳe`�f����:�����d}�u���#����5ǲ��}���ʺ��ŕC^��jr����c�n�u�ˌu��n�"eyㇽ�Mr�U*��t'���+;�
�CV�TE	�oX�J}�c���������q��Ht%����z� Ӣ,k�o���'I�AЙ�3��R�s����,�oɄaf=Dt���$�4�s����~Y�g�0�w��Y��R����aS�g���&''Ӵ��j`������/�?(�}�d�ff���e�������~[_Y�t�����0��g��>~��$��1V�C�*�k�
�m�^L�o�ڔ�1�[��DܘP�-%�Ih���W�=#_�޽{f����Q���l4P�����U���A��{�r7�(�(�;�iӖ�/Bz�U�O/B����X�����@e.�
�
b؎�n�^�F������X{����%�^�]/�@�+�Ɯ�t��SP�H.>T_<}��ܙ%���hn�\��BF�#����K�R�݉���ةP�a�+ 6Y0��E�WVԔ$�ҥ�=0��"i5;�aB�pBL�r�x��L:,���,BG���'�;�[���J�@�It�9�u����G�}��b��G�^�HK��cR�?��n'�Ǎ;�.sp�+I��&�q9M�7ҖF�U;U��פ8Md�`���;�z\�'I&'�w=��R.���J�s)��iļ��uA1D�
�CM�bG��Ҋ����� I'�e�����������(xwF䎎T%@:@����t�M#8��t�,���꒼���٭�ޢ��tld���C�S�o��:��8>��ʱ�aƲ`��c�}
,`/@���h�BEm��\��+ˉ�t���]�P[P`��h*'1~���S�O��r�J1����,��T��B������7�����©ё�ҙ�Z �N��oa��Y���ԍAT^�w��b\���*�n͏+.���4�F��Z��b�
��ꐳ���H��'�}������9Ÿ[�߿��k�D֗�#U��$hL��n�CI/p��e�sG�/0�n����(�;� <��dGz97��kՐ�&�y�Q�$p�;���j1i4�"'.��|n1��,�O����v{��OU;�<�I]=.� ��E�ҁ�5Z��2�eW�9ΉtN�����]R1~@Y�I���	�3~�&�)s�n�/�:M�����KT>�+B��F�m�4V���;"���~���({����9Op�v�����#�W���F)̿"2�Bw��n�� �Ns���Ry��l�rc#���뷐1]I׎�t�O��'��~��IPJ��Re��d�s�ɡɧ�(�\��G	N7t��`��9�hu<��P0�NSzc��1�e5_��UJ�$N����l�a�T*�#G�H�����9����4������ӓcc��N��	��ڱ����ȡ�U;I��s��#�NU��њ/����\~�O��<�� O4�%�V�J2���B�rF�������J�	�׫�����do���[��8�s/�9�cP�F9�{��3��H��8��|�64c~��1m+�v6��h��Ɛ}��k�i���Z�}�L�����P��6�|��ñc��kb6�.�l���4>	���^}�|�e0ToQ�c}#zb0�q�"�᠌�ö�^0�.����vA�Z�)$�8���|f���m��#����r�sv��~�О���sb/�����X,$�[pؓ'c�6ڒ\*r��ij|N�b�������\QW�&f��V�;Kk�$�����m�/ٸ��-t[���8�&&������B��o,>�I��'Տٟ�a��T�t���	�J��3g�xQ]���1�e��x�!#u}�p;�d^�%y���T��9�B�M�<�c}�C�����焛lذa�\z���k���ZS�Bw�z*
�4Y��Y���~�t$�%�w��U�y_��&*GsT�&��BW*����z�>x��s6iF�h?1�ʥ�%�W<9�"%���B�W��5k�`�W+��/�N�q���b��b�
 gb�0�_��NL�H�2�@8^p�u*�O/=��]333���}g�ag�4��J{���4�"�2��Д�Ϙb\J�Q�Y���GW��Ap�N'\Ynp<L��Ǭ���"vFv�ҡD���� ��������y�4�F=r������f��g��R�8����(�f�';V2����p0B��8��6f��[d(*��5�@>Hn��߳Eqz���0�jأr���ʒ�J�5�>��m�5�A�hJ��i6����=sI�}����C�.1�9lz���󩹆������aH���<�o���"���B�P.�T�M��L0��B�|׸(\�gV�C�f.���~vcv���@i�����]f́p�����c�3M�|�\.�$O9�x�P�d��%8'J����nU)��`^�b�b�L�L�Zپw��eݨ���ԀR11���J�`l}��Ѵga~�Y܁-�Xb'���F�~�4r������f��7��D�d	�R_|Qq*�R��"�H%�� ��z$�����
�e�]�=C��QY�� ����(a�\�7�FB�"��qyz֟.`=5��~IYd������P��Di�R.��!��F��5��C�o쐄۳A��*Yњ���t��e`J���K����*ο��%�N��p���Q�|�8R�@�OOո@�4��G<��q>bvH�+A�\XX��,�r2�XM��W�����RŬ����W��ȃO`i*�P����۝�~�c�n��Q:�FNb��bN�>̞4vՀ�˗3`\�I}���0�(;��E�0�{	+ֆ�o�Z��MĤ�&��ы�}bOY�@[T��,���[�V�R�!�gU����¶jǫ?׌�-�ܛ�m�>t��A /~ٴ�rU̧��!	S#g�~���\��1��`�Z���σ��*��i�iD��|Z�IHB�������=D�iT�����f��
bN�Q��'�o͹�iE�j}ǶdK}�l4a7;z�1���}o"��R���nrV�~g��d�Jw0������hR&��Ğ��Zy�v�p&M,R��4.%ĘD��tc>e�2W7U�.�^&�HD0U��,����H���f��&�.�R�a�,�R$��1��5R��R��'@ω|#��I!�\�ǖI}�ʰ�lSZ#��]�t�-t�SL%�ϳ���|���FH�K�T���x������l޴i��q��N�Ҙ�5�2kzn1��A�����55�6�o�3.�>\�#D�$�c�
�G��s��{�ޅ>�c�̞,H�N��R(,�#��Zm'�V��nv�H��n�M=�>I���,{X�b��G���P�>���3�IK�z�v��� �?��R)ڶm�-���)�͞t٣k/	>�Bڄ.���Ν�y{��]�qp��I�'�z:�h��.GW�]���p�U��^���7j�=�� IR�5̴?���;6Ř�䟔I��R�	|�֐��쌳�{�Ր�MR{c��m��8�L�g����DԜ�}e�Fpj!J;JR�M*���Qmy3#:kd!�ũr��W4V��(Zm>�U�k2��9(�.ly��aDY������fE�*C8�d�'10��i���L�Of�Ɖǖ��Y���U�칕ZVQ��fD���.S#8]*=���@�+�����ŔZ��܇:�x	�~���O�G��<�?V�X���Qz�p���;��lN��đ�f��廐���Q]3g��};�7o��b޹����R��c��� Tl?� H%Jb��B��]�s��|���8=���`�y>�_�Tgn�8�_7������O9G~<J�p�ԗ�o�k�t/o�e����������3i�:���t��7�,Q�EO�K2�T�Lb����e�R�����m`�%@	M��(�W�AZ-sN�����o�c�c2K��tQނ?�`!bjd/�L]�!�v�dUi�-Q�$Q7�H��	��z{yO1*�pf�,-ET����sZ K�(qL��pBO��` +��w�T� B[u�)S���`��WS�(�#j�۞~Z��j�X(S�LhE�Z��'W�/S��I~�Ty(�/��5���?v��Ν;�L�Z0�r��tݔ�(���uS;B�\�#��x}�)��޽��K�'���R��_�1҉DiovAA)b����|����L�����O�.�8W(��OJ��o,�/%�d�V7Y6��dIVrͤ������/�C?$_�~59�S_����G���c����;���,�z-$�y�����!Ҏ�'J�4��,�/�� �%�[�h�P��\��ͬe�*sC���&-��;K{��E(]�?��l�;�%�E���W�O�E�!D3�������O[u���d��z��ЭX�9���2ˏ9i���	Lˆ�N��Y���Ď��o�>�a3~�*�HuH�L�=Krڰԗe�{	p'�:sorq��c��5IPɑ�!������t~~^w�U�������:�G�E�g����	�?���I�I��XK�X��9X#�&<�Ό4�^�jf���T!\�m�L,6ӕrA������ ��d!|��j��D�^�g��+��@ډ�N"��c_�n�+'&&��/�J�ޛ0�8CF��]��bQ%�!��
�;Id,��������`��5EL��0�"�(�ʺ���h�����A@���,�/J ����pS[�i`�Cl�7u��"�[TYU�'����v*劰S������A������Jz���09��S)
�|��]h���C��o�����k[i�D �ji�r����x�R���6k������L���3��lX��t~d�ȓ]$M�c�A�x����!0#i%n����յ��Ȕ�[Jw�$��~ٜ�u���o��`le���#�R���\�'��'���v�v3�[f��_0|�{uv[�ܳ����-�4�w�c6�ɔ�WJ�Q��Ab�Oȟ�x�4 ���? >�^�zzv}žs�Z��-�͙�V�h'A��x��n����4e�id��C*i!~>�rd+�M�9Y|�wS��f�=��z=����}-����MaM;�\�J׉D >'a%;1lmq�V�<�a�v�z������K�=v,�Z{~��*SW��J�b�Q��n��D�z\�a{��I���|��I�KTKҍ��E�s��#0�!�%#uƝn{q�e�E��(
|`Լ�H�γԏc�kR�/(dd_���qH&��+���cLVx�!�)'�$���[m��{��	�p/_,�k��0�O,��ANhk�#��L� \9W��	��!��B�L��ё
��$=_f���F�$v�'n)����4�RD?�߁G
���"�Z���++6�0���-֢�T{(U�3ty/N����ʕ��\>��zT�V*M��C�i�f��x�L:6��P��I!b��
yG�`�We������Բ�%�"�Ə1[��L�����gzlb�����X�Z)1��4`������B`�Y����� ���?~��`��R�TI�ݥ�%X��i���M�V��aw���=��o�4���U����هJs7Q�\]R�Mz���ٟbeV����c�/�u�;�=#̈(�fȬ��̍���tYQ<��Sv6߀���K}��v����ڬ:c�i+��o�W�jH����Y��8�d��J\|�����`���l���VK���L��ԝ<�F��'�7�N��e+�ZR����M-\6�Q%%C����0c3�hO������JfrDC3m�w�R]��j���XW	��:�1��!կC؛%�l�&[�PgQ�����>[__�� T�w�,X]'3,u�n.���DS��]�0�"�&l�5�d������ruB�8�;/,,h�DƉ`ye�5o�[��`F��"�� &x�X�F���WR��3������F����Y�u���E<"JS���e�ک6��o.KGAE7��P�U��O���n�f��<ⱋ<���cɁ[�{O����#��>!��,/���v��#�ԟY7&����K��e�Madt�� �z��fw��	��0���R� ǳ���:s�̚���îe��r���We�����2Ə���֮����!�2�{^֚9��I���{�W�TO�:�{�n�̌MMM�P�?�|��Pc��r�vG�7�'�� ��ز}��؆Ç9��׽"�M��b��� ���U���(�)4dp%uB�UAU�U~�Z��q�~�K�5MZuO�ԼB�<�P�0)�b�_�P5���3���]&t�6��H5���hm� HA���P�1��,�v���FyL-�Z�6���J�"�e^/�x����9:3�>fff���������񎸼Ѩ�,0fL'��x��BːJ4iYn�4�TeR��:���x�핕(�###sss2<<ۿ����$��>۷o�a\�RM�$�_.�*�b���Y��a3G#�� )J�$�����N̅83�V�/Q^o����3$l0R@��lقarC,����כ���A����1;;��@ �0�0`�ƥŕX�&MO�8�w��YYY��N�KwB�$�  �݂ps�dh�0��=��cJ�չR��t���`A��|Q~��Gʇ��Iv�2��5��"�\�;Y�N�&�fw�����J"�KI=�+jc�[-�eg@�d�mn��K��%���4J��B�p����R-qH�!$G�x��AZ�$&��Zi|t$�}��lQ�uP��:m2���g�$y�aӴDw$ҡz�ci����N�F\D>KKN��|�"�34ڱ�9����heu0Z�R����)�jcT��f3l5C�,���8PO���BG��b��K�xy�/�ʋ�ġ3a�q؉:�:$>�SnEw��E�!o���fjj�d����x�%����\�iw��ڙ���s�ic�45�.Em�eЉ�-�ۭ��&Һ7���Ɋ]Y��	��4깅V���x#��aG"��i��U�
@afu0����`{F�ڨ�'���[9�n,lu�"�����*�4sͦ��+M-����wTVԩl;2�b����;ǎ�8�Աf�C�bx�zD� Hx���|�!q�Jibd���o��.��;o�a���5k�`��p�y�a~�[v��a�I����U\�-{PHgb�����͕�o�{�������,�L����]�;�� M	��U�|��}��2��&7��՜���u2c�YŮ�w�>zgݐ>Hs����b?7!�w�֭Kˍ�z�Ӱ��D��D~�ƠC��Oj�Ȣm:�����@ڎ�����7�S�O=�{#��&�ܰi�v�/o�S�� #	��d�&��g;91�
ړ��=Hs�<�'މ1"i@�v�Zhu�51fV��q�FH}!�
߈��	`�� �2.�f�V���|J�f^:f@�P�/���� �Vq7**�%�%�(�r��\���U:t�7o���׿������~3���|��H�S�qOG�ԯVA1W�o}�; �2��i����ŢT�7��C0�!�':�-�,N�h+�>@��U֖Zv��a2υBN Β�&��b��o� �Щ���q�\���f/�4SM�(��d�H2R����b�*�ԭ�b�rƦ����D,%�8�ɥ=�W�k���-�K�ٕƲ�I�6.$�=-��ꉧ�ތm�zm0�g�I���i6�M/͟�el��%��P�aJͺ�����ex��{���4Z����.�9�'��Je����ĉ�0^O�L*�]�Y��Hҏ�KK=^н�O�m`��6Ԣ,Ƕ�sEYF�fQ��M������a�Xà�=|KcX�ܳ:ӳe!��d���9���ؤ��N��߭��q�T�w�	��;��;w�u���T
I���ݻW���>��.�U��36�#��(���T�>���x���)��x:�/��r��!�M#���!�apx��Ƕ����(�-:ɺ�0��p�x�\Ppu��-�0	0���v�<8��7�`�-�R����7aB�{�G��@HŒCDI`�A*�	��H�cĘbK��(�v=fS�|Ʋ��Yx��$��݅5��pvE�.B��YrY`�z�e�Ϧ�)V�����0jJj����Y�ḾԌ��>�m	��`��N�<�AJ��F���il]�30�q����}f��.Oc�YNp��wjz�:�v�Z�aT����20L)]�V��:Wq��W
�!��I|��E
l��;K	 ƃW���x;�?6벛J�p���.�XgXCr;���AKƅ� ����)|�(�y�r���1e��q8�B7�E�#'S��5�1��l%�3�-}!���0=`'xB���}�]�+J|�#iHA�va6A1�`�`]�J��4?��m�8�f�����A�7��y����m��xG��N�.
]-031�ݳR�˃.�nH�G�b��/]�T�N���	�'��.�Yc�̎����!�ѴS�>¿:�rA�~��)�iT�&'��1�O{勲�,���Y&%hL��wFf�G�tU�~�q��T�.~�v��W&<�k����sub�fm���bW�Nڅ1���\񢁴:-�j_�?���e�S2�NFQ\��90a��b�Sw/~�0m�Z�:�u_��8������h���Q���RPb��U�L]�����"
��*���d�nS(�<ħ���4*��x�;�+[�����TnЩ�
M�]��.�m�'�f!�_1��K������x�0NVV��墣]��aY0��ߍ(N1GS��f��-WjIJ����!���U�2��/�/�u���Ł����k6��q��:Ǉ_�餾a|�����a͆j��a�>���r8y�iʀy�<�a�	�D"�$̈́j!
U�n�H�|���w���O^����_x�K�WE2ɳ1��L躵k��o�vϞ=�b7o��E�JB���qL7�Rm� 5�c�);6�йʊ.����$B��8[×���>7"�*�HA�TAH����9ۃ�`�+�62ղ4������s�Ht�7�y/i���� ��谩�/AƋW_��#
�trt�����w>C�:ۼ)K5q�<pR1V����[Ǳ<���캢�J��O�>��#��&�Pى:(�Y��WҶI.����af)͜���w�����ӒXQ�6=ۿ]7�I�3��h���c�R�HV���	L8�PǱ$]Pf�F(�:�EB�ƚ���U/���W��_�h��S�����RF��Ms�^�s�U�����rO��H��
��*+��a|)���%e�޲�e����V�r�w�����I�yk�h���nGҳ���W^��8"�8C<f���D�&{��$���6�Z�͜�bc�Θ��v)���J��?��,ˏ+f]+�CL�,~_'o�T&�����I�6-�E���:��%��,�Z����i���X�N"�#�ͻd���{�NϑîP���b��0�#G44���e��RGO0��l���֗?e2+�d8I���W�i����w�;��G�;���f)G�R<�BQJ6g�V�4��7��������;w*�>o
������+������³��|,qߊ�*��R�|��r���ck�.��RC��
S�!�-�jο�������ߏsF�a��	p�Ԙ�4����ӭ	��Y��B1L�\��$�(����J�Ʃ䊀�k�R��㎻N/�?��Ͻ��7r���a6B�.�� �%ٶu+��<���~���c�\r�4��3Ϣ��Ѥ���i4�ԲPiޙSQڰ���T�5����8v3���_�����Zq�9�+�1�ʒ�������痾�%L�瞇���p�1��z���K#x�f�M	����A�OLN�����{���?�y�S�L�9B?}�ᇯ�ꪏ|�#��Go���s�9�T���2wڋ�����,��1<��	D����Oq鋛3��}�����v�ر#G�l޴y�΋�R�'���̤���hvJKtF:�/Nt�J��>\#�n��Sz���s�=���;���+�AB��&
�\��	�|��/�m듇?�Fj�Y+���2��^�F����������cj�;����Z=�s�i���v��./O��5x��O��;��e�O��τ8�O���o���Y*(l��"���l�,�/$�/�8rB�]OWa�c�N�J8�S'����y�4�08��P�A�����s
żĉ��򯆝n��J�Le��éxR��z�#u:��L%\X$=�I�_Y�T@DT�8I��ͨ�x��S�z�t!��� ��^�Rr��ﵚ:ax�AO����3j p�cL���@N2�8�� ��uV� -�l�"��/�8L���BMp�\^9!�/N����P�YЖ��taI{NP�:q����|i$_*�8۬�4�����ۅ-�҉�a�F	N�Dmp��Z���l���B}O�����l��gc�*p0��5S#�~&�����#M�z���J�0tJk��\q�F����Nml����P�����)/(r4��/�\y���k�X*N�t�uR����k��y���-�%ψna?=�_P���Cq�gb�`���!�
�B�w���R?��8"�߃�ǘ)Q��{���z/{�����۱c#HU
�r=?�T;T+E�:tw~��o{ы^���7�0�p�Z�*1o�5��9���aX���e�t�{�E�]_ۣ�}��mٲ_BՀ����t�M����P��<?
�$*-�o���W����Ї���o@;�F%0�{>�L�����I�����1V�(4v�Di�!m��^����'�{��Mo���?�)�F����d������PJ~�7~7���?�gϞ>2f�y� ��)�|�\z�^�ΰ�rs`$6��=z�c�k�y���_t�E7�p��Ԕ�Y�x���{�1�[۷m�`��JcÆ�K�쑘Ǚ�����7R���7���J���`@9Nx�X��[�8p L��/�`�K��%���=r��-���F�H}���34{�~O7�+_LXB�P-�Ѫ��Ԏ}� �+,nv�I`Ӓx������qk9�gWr,?M�-Cߜc�|x��w+<uİ��|B̯l���i�Lo��9��唪��wy��c��e7�K�z_A�s2�,.�����D��$�8�"�{��3t���ׯ�h�%8�r����Q(Ǝ1p�C	���.�C�D2��d��7�pa��j��т�;u���q�+G�?��O'�+��c�.�-H��-E�w��1��P��K��7�K8giyB��ȒN��6T���yn?kgj���N�N;��v�sW�2��?8<T�׼&�����z��������֗}-�u���)Q�HMq�����ԧl�EyH�ÉYs��rq��ɓ'Λ��F��e(�3襫�-�>�dևP&���1�;�c���:I��9~�ԗѤ�Wc��ex�Z���`�߭T�"�Vu��� z��c\�-���|��؄���D�1��z���}���<'V�T�G2Rs�X\�W���[6b~��>��-��������?T����~�z,��g�7R?���L-��s}�CR��G@A|��}�V�)m�KY~��TxT����H��A�5�����{����_�r��|`n%=[|���M�$��)k����u�T{�\�%I��}O��+���/Ca�V�XSP��%ONz�W�w�}�a�{�k���9L��]pu��leU�Ij�E�yK,`Z�QhD-�i����C�k�y�+_��7�`�װ�wqwމ~���v���R���=#>5�N���[	y`$P}�_E䋋O�T!��r�������׼�5���'���v��U'���+���}O�������ƺ�#9�u�r��:�G�k���E��9ؠA>���!_�Ѯ�5������>+9�Z"�:c���ǻX �b�4ꭙ�u����'8�Nhoa���۟%+>տ{���>%E]HF.SC0!Y`�.c?�I�҄��.�f}qq�43��\@�	�:�����f�F�NC9r��}b9�
�Ea���\���e��F�#���t�}W�����8�����!2�5J�p����NL��P�1�v��C�� _.��r.l��@��v84��:Fz���x�<��&A�¸�y�ȱ�|�Ҹ�Uf&����U��4L!��\ o|���iG�f��&[ܿB��n���\Z>1;G���N�]�7I_	�)ET}�eײ��]^����z���͓0?�j�����םy����H>�>��J! .��%W�����m}�º
���`����e^Ѯs$�D�|V	���z�u��m$jtl��/u�lL,��*S�X�4̏Nǡ�*�IY`�*ce�V�<V� �n4�;�q�W^Ĵ}�t�/��ƚ1��G����?�|�޿���y�@k۔�L֞ne%���r-��]J2hv$(�y��{�_��f`Ðl�j�M-X���T��4:����������W\q��?���������I�X�4�eFe�P����Cmtļ���P�@�����wOO��a�DY`�&��@�D>�j.�ׯ_�W��O�� �����O�ӏ>��{�e�5,ǪRߠ9V��"�Z�ۮx�s�Z�{߽�֮���}��oy������xuX��3t�ƍ�U((SS�y�/>|���o��p�e��i������`{fʌ%�y��8V�#�H�g�}���?��R�|�|�_711����9��J
}kii����g�K�����hÁc�UB�c�Ɍ&!QX)+0y'u�	���w�q�o�����͛�t���pC?~|n۶m���g~���C�h,C#�w9"��&]�lْ2�&~�G�B&作\O!{hE�IAzW����\�l�x��,��c���9c+���ԇWVYJ�� ,�mկ@�ꂹ��f406\���z��ȳo�pv*�|�t�̘Ù��&6�cT12�Z�xDb�a���=�ə�-��������fC��"_�LB��axK�2)���"���\v�(�da�i0Y'��xFeq�y!�?BX�Vg`-��b2ggg��I.0����d�./5�Q!���b�@����u�{$�t	)�דďs҄҇�U�!r��魛f �׮!�=�n7�4�3̘%��I9��X���jV7`c�M$�����i,}m\9��P�1=����j/�Lg��xƼ�G�B\�5ٝC�;�s YgI�ǟT�ݩ��0"�)X�~�nڴi�֭?�0��]�,�O����r�5��t��ZZX�b92:j�u{8	c�:+=�h�<��3'x���C�Pcck���Hmd4�;���x�Tr����QHAE/�P&��ow��z8>���خ�X�����7W7�؂g�ڭb��(u#߳U&mf&++�p!U�b��Z39V��V�����o~X���P	�y��k$���T��+�'�C�).�%��Q�z �>��#W^y9���G[*��O����n����`S��gR����0���v������]����o��m�{n�q]N������74�}K����!�R��j�+�E��L��̱X(�Ϝyꡇ���O|

;���I�� �T�[cS�?>��mڴ?'N���ǣ<�����w���G�eW`�p��Q!�dؙ 
>����=�.v����O������s�Z�L�V��zlrb����Mo{���x�A�G��[aMJ;�h�5�rw���'����
���/\Z>����/~�Pb�+6{A�q�7�J �,�+�ʥRO�5K�ڜz>��h���fƈ�+��S(�T��{�Ϻ����oo߾UqW(O0�λ���{�V-N��n�tp������w��>����vC���q򞽏����s���ԍ�j�v����STS�@Q���GYSR0��uGơ�-��m+K�������6�/)�s�<�&��ݳ^x�7�>�{t�c���������#~R�������w|�?�����T:�Ȼ�t)��!����$�����p��䜷�:2��E)�\C2���[��q�J,�r�\��*T�����-��./>|r͚Ϳ��/j�ӕ�R{��n:k�n]31�:uj�ſ��O��થ\�)�s��m%�3`��|k�ͯ�>�f7��U�j�q\��`=�5�}�fN�XE��q�4��;iC|�
��
�9�8-���r��+Ku|s�Ё�^
u�� (����@1�W]^�֎?�m���q�
�]jKgN��vg�`���9��%����R�X�Q
p'd'R��'��A8��f�u��H.zN;�N��т�u���/�:]�sL���|*W�;NM�?��}7��l>v��]����N��tcwa���x���Hu��!__�Ļ�<xx	ꍟ�*V�Km�����v�����Xhn�\u�����=׿�W�w�a�y���Tj\tN���/Ϲ0��$\(�jG��H��JG�f:{|���m�ϟ��^��:yr9G1Sw~ai�y�(��
@]>��!U��|M	'�S_+
�<F�	w���DC�@�v[�V��T��n��;8���"o��^�%�?QR�´��h��#c�0*�'���7�@�#��B����q�*ac`{B��������2=������'ǫ�F������&���ZQg��nS��R���Fv��SO=�ࣟ��g�&����7)N��K_bt(c_C���b�x�ŗ�?r/���ߞ��g}���^�|�:�~q� IY+�%�(o~�X6������0�~�6z�����%�s�^�%�VwrrJ���ÍB�ĵ�Qpή]{0�?����%/y������w���yآlx�).#HA]%:e`��Dᨵk�;��C�i��?��_x-c|��I�+@�@ ��Uk�|��@'�����MO���`�r�o}��k����`�~�s�ûc60L��@ a9v��!������L��,�X�%n1VL����?�������|'���'�u���(~� 0Q20���`�(׮]���O��ko���O����/�$$�l��*�]>H=��-M��eWA�c��Z?8�4����j��{����o�y��͠����Tu�!m߾'�\�
 ��gN�)�O�h13T�{�o�|��o~���������1u���N��)���`���ۺ��n�y�fR��/ps���#3����ꫯ��[7�DA�%���*lZ���-[:���]8�wo�yϮ�����⟰�]vU��S�����S���� ��Ss�dJ�a�x����Ъ7p���Z|�g�ϪD�(S�F(�����߻c�Wy�ΐ+�8p@��cT�ϓO>������ܹ����d��]+R}MJn�f��P�"N%�8J8B���lU�;$�/bN�:J����Ն$��6��!9��<�8�|�W���PN�����r��,M�D~�'�x��x��>���|�+�>����^�n�nT
�!�@'�:���仾�	H!s��˪z������~L�'�S�m� ��p����G����ڴiG��|뭷b��u<���=�ԡg]��n��J0	�u��q,�#e]�������iCIe�+�$�밽M$�B�)Hf"^Y|��V���cx�r�<��*��[�W��U���cGf���T�L�4�ؿ��������KHd�����G�DA�vڷo߁��0��Ɩ:Q�g)�Ǚd^t���N���0�j��%2�{���ڵ�?܅�?�Lԙ�&�T	�q��hj����#���ධz����\t�E�?�-��j��Y�AHSU*23�L�c�� ��.&��@
spf1�\��v�j,�E��s�`�4cq��/
�a�xq��5�iÃ�dz���~#J����s�g�$~�Ѐ��K}GG+�%����c�蒋�n�v�w}�[����g>�W]u���4-,.I���~�m7���=��7��u׿�E�X���rÆͮ_�)416N��̬��\�R�14/7Ud���U��f;�Z���
�m�ϩ����{�*B�"�I񵩬;���O�G��;�㎻�$�~��a�MMOB�5�N�4�.�MKXeϞ'/�����ɗ��/��Ǳ��9<�.0��+��@U� �xa(rV9h}tt�3��̋_��j�L�Dq�$�����T���
F^$U�N�"�ݙ��LOO�g��?� ����o�/�z׻~�����ׯOu��iӦ�,V0t���,����vRJ��c���a{_~ť����Ԓ��&'�%�#%ڇe�@��ag ��*�]����~|��驙O}��7�x�����~��ߛ���K��c��e2%A	�= -X�b���(4[�㟶nی}A �{寿����<�d$x.�:UF/��R>�m�����S��� 4��mqa���
�>��ϸ�����׾����̵��ة@�EXb,��/d�`�A!�(Ai�BGp�(���a�����O����sՓ��*�_8�G9ozͤ@ ��v�<c��z�̫~�5�<�����R�cM�g�]������{��8ܴu�����?u[�4�E�9���;ȓ�k4ۅ$�l��:a^�`��wdr#���'��k^��K/�<V�<9w
�jl�V��5���f{e�|�fz}�z{��;�t��憛��G�?��g&F?�K�>#�k)��f�VF q���G�� ��5Z��|0�~̡���[|�V�ϱH�lq��"��Ʒ>�y�
��맄��9v���[G��+˹�����m�o߲�����\�W�W���iӚ�'磴�l-��v%_v?l��iy9jE�j/NL���	\��i��}˺���F���c��T�
뚼����ôw��f��_��7^s�uPn�<�DP�nٺ�qsK`��;�������������ğ|�S�*W����`;�H��=&��2V	�rjff��0�)��&���3��x��^�#y���q��̆�ӣ�p]�s��>��>���[�9|bi�m �g����(L{|�����#���!vL�����W��/��S���C�-���#F��n�b�DY*�^u�������R�l�:v����1O�O��;v������x��?�v�����f�q������ȯ��K?�я�ٵ�����ӝ.�c�J����?������K-�G�^���n�U*p��ɶ��D��'�Ͷ=�K��S.A ��M��K�\t�7 )�hS̋�&z��8��J�P�ZjƋ��V'h�V�ֹW=����'wS�{���ASD4	)ۓi�F�j�#�pc+�0s���<��-��'�?d,�����)�/8w�f������RB�[c��u�]d����(u?�
_���S���O��_L��'>�w��zX�{��L������kǤT4S�M-Re*�������;.��xm�"@9tY�mQ05G�6��c��>ɑ��G?z�w�r�7}�����_��?�ԧ_���f���26+68~|�獵)Ob�_���k�����o|�8*�d^du�|`���N����
�~�[���׿O����	�PwY�g�؟dŏ�������_�p�3��w� '���@�P�a||�\���G�*�����}����o<z�(�I��_�#����"�\.W�{��ǀ/��,
���Q��HM�������
���6�dS?��c�Pر��'�y���mۿ��o�˿|�mo{�����ŪÃ�A�q1E���%����W��@��|��;����Z�yl�D� ^,�V'��\.��0�a�<o$���wߋ���_�?��_x�{ߋ�1�M�6�L��Hy��`Ga/��X�E��:,��y|�#��������wo6S*�R(e	�@�=qɚ�IS��9A�F���_�e�[��:�������;� _�r�>o�߷�޽[�M�:�%�s�"�A�Q��ǧ�����T1��]w�/^s�r�n�y%<�Iqcp��|E�U�y��aX`��ێ��v�mx��^��y�%���`�&Fi�㈘W��d��d�M�1��2A��o����I����u�p��D��NS3�˯z��}�KI���c��V+a��6fRʠ}���������Z�O����׾��}���l��z���O�a0�\S@r0���C)N����l�M3��px��s��`�K��K�֧�,b$׽�u��nvs�����{��Z/,�1Kkg�c��2�N��}X�?����u���?|߭��z�;D���&D<��.�c�A�euJB��TW�g�+~��h�u91 �|��+�/�B�cN~�~�Y�~v�r�ڿ�P�$�v�D��#���޺s���|��_��W��ͯa�q��.�c�{�1�A���qے]�2��˘�B����B<0*���ŗ\r�e���Ì�M�����c�Q�1~�������|��#G�̝!��9眃��a)�_}�5���?��w�sם��Y[6N�9�Mq�Ҿ(�}�?KCi��Հ��q%)�9�*�+U�8�J��]T�9�s�<��@�����%.�1�i�zJކ Kf��^�N�6�EdxS{��T&p9p�O����lqsI��?�Ͽ��曧f֝:={��q�.����_����rY�4dp�R-	��9��w
�q�,/-oݾ��7����o��W�j�Z[n�N��Ԫ�"��<���H�'֮[7q�3.�Qͥ�쩘F�d�7��J��
P/�N�vYQ|�3������~��+�<v�؍7����������?��[��֋.�9>V����uӊ����(~v�޻w��`m��~�W~�[n���?�[�]���WA|,_G�������+�����O�$�X�1�[�r�蹹�{i��&Qz���/�#|��}����^��nz�^���㮀�b#0��{��͝����;gO���|���ׯ�ٟ��Lp�r������0 ���t(۱��o߾��|����W��PȢ���V<�
����A	7�t���׾��Y��P��x���ɩ��H���ø�u/z��cO}�C�]\\��Ғ�CN�����EY{.�>|[��c���x�k���wq��0��tJ%P����{�U��ZUIyRb(��ؙ�A�>��k�i�k��o���l�{��������R�X3�\�t�4�s�E�^.S��ʉ��b��������=�#�29g��`�P���p�����/�ȧ͛76W���֮%k�=+����>�}l7X�[n�����}�UU��9Ǿ��t���H
���fq�f�0�1gǑ1�"fL�* JNM��t����W����?o���]�^��{��g��U_ծ��ǭi��H�K"�;=-+=-����M����n��5YB%%x(&�
�����5,Fc�?�+4J����$C���)�g]p!��㹽�}�jƎ���j*%��N�?Rk�]m[n� ��HQ�j��(�N��i������t���g=YC5�Z�R#������
� �6��������D�����>�B�Qc��>/̹�{���e�U����r���cw��Qzi8�l���u�����Ne���y�=�b���XТb"�ؽ�h^wh�W�}ޥ+�ys��ͩi6GN��@���G+�N�cV�.!R�2Fi��\�����������)L*���)WÒ��ԍy5z��ٳ3�)����-�������& �/0��p!o�'�P���#&���h�G��g�=�����-#�Wt���RS(�>���<23�L-�� ��$����+)%�J�Y���CS�yB)w���~HN��j��h��Ǖ�\v˄	�Z��^����j�>����u&s/�ט�3Zb������'k/���\��/<�N�B;pdoT2MV*��"J�t��lHl��
_Q$QR����C�P":���v�����c���w��	��zw ��؎4�%%��B���2c��o�V7����5[��Ee��,�}���������Eǎ9|�hEY���_=j�Y@�ǎ�.�Ͳ��������4�ə�Otťr�O��
���SPsI��O� �	Y,��(�R����HM���+�t��	ѹIm}�ͷ-)..q����D��ח챋�P�\���(�^,���������&���a��O6A��dB��Z�[����j�5��Q:��$�+�;�H�Ҫ!�C�>/7�W�*$2~A�7I���7�6�}d�'N��}x��.�Ro�y�Ə�S�Ł7���M))���y�Ud��Р'ߴ������x≶�`ұc��j+W�f����W�X�f͚�K��r�-L���,jw79���555-�m���ׯ����l߱}��x�� Ҕ��y��s�g���k�.6�N��2P2����0c'N���a�_y��T�:�6����;�|�68�� /^��ή�,�i�i�f���e��y�&Mz�ɿ�a�����㑹[3��/+pe���Ǿ�7ol��I��FaK�\`2Q1��,�0F��3� ����}��k�~���s�9I��Of��� ����=�+#F�x�ٿ]~���?���={x��C�@�/m��E���V���W_}5VM�&<��f�p�Z���}�!��]x	�s��s":>���(�׏��s���P1��%K��<�aFd�n��~�)8=�_!�L���X���>��-Ř��R,
&k��CN["@��`n)e25U��
��g�9x��{U��2%̦z��|@6ջ	q�̔vI�` ������	Zee�w�% ������*m���C��Bahy���KP����r�2tF:8�bᓰ^���XJ��Hg�����/^�����͛7���@6�(Q����L� r
p4���b��/���� 7�/_��b����n�N��s��Ϗ����Kq)h)�a;�:|l�ԩx��۷cT��,�3g΋/=-����I1��TJ9���H�Sf��O5��-��D_x��+V�<�u�p��b�n�m[k+6.XTTt��	l�֐�|�6�'SW�*Qm�LNN�������{��BT�
��p�R���d��0�W�2Ⱏb�����#����(�l�����ٙ���^�h���{�@�d
��M$hV�g�D�Cb��i����l`�x4���_���}�}��.h`8]�GE���#�gy���U��2Y���Y�&_%��pY�p��������-=�N-��"n���Ç�N7y�}��Ro�������r�^�#�-lm:��SKGFf��W_}�`�?� 	Ǌ��%tP+?��T�~��/���@6�@�R�C{GqEb"�F�-��*���F���<f�x�AKK3��='w0'�%kİ��H� ��z�r��#�����j�
�Ox���G5)�����V?1�M�����ܽջ�i6�#����:��POoW�=U$��6�"n�����ޟ��Q�$���;dTY+�Yɽ�=��b��yط�w�:p���p��i*R1�NJP�T#}ɤP4���@��J�p��������/}��c�N`�@wŧ�f�p���t�F���>�������lٲɓ'G��6��
%�SZJ^fkk��={'M������SO��V�fƸ��l��8�Z�oܸ3"aLӍIVp�'b7�|:5����TU5��b�[�>�]�֮�>bޖ��!?�c�=s�}�]q���+������A���e�}��^{�E@�s�=w�O?͚uޮ]���&���Eu�^H�]w��VRR�\�@�O��Z2���a��2�>f��|e���/����/����+..=u�ĕW^�>��C����OY"q/ 7�S>|W�����w�}�����ox��#G�X���<�h�ԉN-�`�6����sޜ믿��C�0wR�_�Ovw�>ǰ�G�"���o?��#Pj�P��~'��K.)//��̆$c�P=��+�W����V�1cƁ{챿���".R8��e��a���������D��ӯ���Ӊr1�C���@l]KK��x�A���.�&�׿�u�=���Tj�Z���܎�K���`4(U6l"�َqz����<C��O?�t��-�zӉ'���I��pG��JozLDG�ф֨3��q��"WvTWgf>���z�G�����2�1=�	���sv'�:.H�jv�r%DO���]�>�����:z���M��B�pMWZ���xT��+�|%�+�AȶA��h����i�J�9D�p���qQ@Si�f�NO(tF�@�Ɍ�vw�=�쁧�:�lV_@��]AGF1�����1 )�2,Js{�[(-�F�j�2�N�r���f���8����X�7�8�o=���.�<�Ϙ��F����)B�1�U�ɇ��Ź.+2���1���
o�$�	�UGj�*�y^=㜹�B�m]ԩvΚ��o=|��ǖ��te�fQX;r�����`�L1I©�Á����b���y�= R��w�~/''=##���=]�'S��8��oL�HPu�\	�M~�w��WK�L�5��8Qפlj����@�{*�RsKf���i�XuzCsk+D���=�a	G��E�����!T}N��h�Ԑ��:^Ӏ-����:>�����T��<z��'7+�_6xP�/
}	E�d��*%�W:��P2�l��gmimw�]�I������L�4����:u\Â��#������oWo����� �[��K�'�O�4�(���[����<�X#E�2@Q��AԍT�!2���?,�PyY"�KQb���
�F���{L��#��P4*:�o���{��צM�����gX�`$!Q�/6(֚�Ű.�,��s~�1~��YE�F"J|N�p<�j��b�2$���p���������V�w�'g�2�!L��xV_bu����5'��fxH	A-��R���j���z�X}�ܹ��[�VY9LIO��,c7��8.��r𫹵�n����67��3��/ y�"���;��'�z�{��9����M��� �0�xj�'R.���ꂂ����R���إ���'L� O}����E��S� ���/�3��t���G�bf**ʷn����oܸ1'�ҹ9���L&�F������/���?�kd�LD0�� �NA��Ҕ)�z{)u��_ +�����o�u��㮨��sM�o߾���g��)6l(//>�y��p�(���&B��'9�D���}��'a1~|������?_z����r�� �ד���1�Y�-(.( `��EW�Ø|��� 97�A*��3g@�a�y�I�]Ώ��ĺx9�=~<����?b0�ѣGc2�mq�g�y�z��q_H`�a�c�"ǎ�P�' �%%%���n���n[�z5d@�S��d��D����9�쳡��Qj���+��k�����Æ�����G8~��(}>GS0�_}��oT��u��X"��H��"b/L�#-��<��}�Ν�0�o�\"�Nyd��ON!.x��F��C%4�K��4F<ݨ	Ա��i0�1�֎VLfN^.�C�� N���NIIٲy n�q>��Gm��Cm��$���N��q�:�DN|��?�oߞ���E�}JW I��x$y���@A�m�|,�U�������n��z�V��FN � P)�~�]۠O�pY�%U� 'L4��alF�n�޽۶o���>����yk��?BE��P*k$�����-��wE�� ���<��.�w9V��	�߿��	pC/�Ke�R[[+���k�ƍS+��P�{\a����z3�(�df&P�?�z�;n�ӟ��{����<���OB�u*�p�9�߹�TE5��3Gؼ}^\Μ�����Z���j�ǌ�^�ꃎ�v�Y�V�.(=8���X�DVv&S�M`���,��x�g �~��������1�wW�]YY
�7.}+Q����3 bQĐ�բ|ɰc�n���wC����{�޹
��z_5�]FF&>o����9�FKi����מ<Y��N�A�ܳ��z���&L��W�&�-�'�Id�e���i��"D�,Wi���A��x����p�\y�5t6�H�<q�����̦*6���u�\����X�bg�KT+��c'[VG����� !�m̕H�����^����L.p�>d�j�0,-�Q�k��my���y<U]]�YgN�hu�������%+;����V�O'�"��؄�A!k�55]*.*�]|(!t���%�SJ�+�Rk �"++嗍����[9>�e���6���R���M���I%��Ŵj�*���
����K�o�B!��3��A�V(���R� ��k�VTT̙3K|>!Th�lQĂ{	��:t�;i҄���k���G�ї�U@��O\��ӹ�Nk�'���Xlj���/��ᇟn��!f�5�:#<~�ϋ���w�f#���~����fϞ�|���zK#��á�c�x��O�:k�$Nd8M���f��jD����x�oq�o����G=r�TfL>���sO�Q�TP0�u�eW ��2]|�]��<��FƏ���;r�ܲ+��]q�wb~�/�l�e�^K��k��}����
L�u%jΙ�8sVǃ���:��,�-ȝ(�6	B{��~��ǘ\�y�ص�!�0:�ŝ@�E0� ��h�"LKjj:����t�~��q�:`�k����#_S���XኾH$�;̝��;��W_{^>�<==�4��������{�����;`�~�� !�v�Y��FSwf�)�R7���9f��Z�ڰ��&$�B�^��+�Ѱ�b6�����I3f̼��k�HUm��Z�ipa��^�v�d6@�ܮ^��|���L<uu��U�mL�C.:�l�=�c�.��rc�9�u����,hZؒ�Su��V_@�k����+6�|��m?���Ƶn���a��#����}�@(�0Y��	OSG�9@ܥ'���P.X�`����A�$McK�N������n�b�����6==]:�RJDJJ�y��+W���__�	��W\�19J�
q�n��j�ɕ�M-Z�~��3�[��]�>�n��;f�Z��{��?PM��V�2%�BX`9��J�l�c�p��:$��[ty����|�#��hDY_S��D�%1Fs��p$HM������  ��IDATIKu����ݷ{ǎÇ�O`Ł�P�*��0>v��uocC#B�K�T=^��[+���\�������I�`�Z�(�+B��S��?@���=��d$E���s�x�Ʀ]�~�(q���TVcN��_|���i<t���?�{Ĉa�5�k�Y9������YZR��Ɛp_������N�� ݂�/�x�o�}��/��Tk�J�j1�飚��8b���¯U*��2m\�wB� C&W��,'�_�bL��+W]y��(z��9�0t��n]%�Q+=�@Wg�٤��Ɛ���Nb��^[ggd�9ӷlٕ�c��^0�b��l��r_w�ʷ���v���(����EZ�����L��їŔ�J��4V�Ue���xL�9)2r��ۭdݎ�Ca*7 �1S-C$B6��/(�������u,:G��Ą��ƈF�?}T0���<�!+;C����ٳ��o8�4m.h6��-��n�����a�4��saW��>���O!SXqhm=�Ԕm���dd?QG<zi�B��f.�)��gH+�UH�;A�F�25u�ș���w���量Q ֤K��dk�	��	���eu:%�\�z%��b��\>˧h�s���_뭷r�c)������7� fd����˨���$��&hel�@C?�"br�x�G��ֻ����>�sڴi�@X$������&�t`bĴ��6�����@������Jۄ3�N7����3�< ���`zz�s�=�
����?���3�p26g$J�|�b�~���fQ�&&I���4��������H3~Z�v����t<LDs�����/��=���D��way�{a�gΜ���ܺu+>_��k�9rdZ����إf�x����ƒ��m���{a��&��@%������1�@l��~��O>�le�Cxt.p"��?y����j��.�dNb���_z饿��V~R/B�T_k�g�j����څ.��'M$T�������MxR��p"��%�� P�/.��Z�%Ce���*"3��@^v�8g�#�s�=��O>��UQF'�z}?s�cN~�����Z|���rɔT���¿4�)�q�;e���f��ݽo��VC�q�ͩ��MG�^V/��;���'O?��`L:��2� �1{�p �!�s������Ӧ��:�U���W\\�=1i'�7��2y���;wan����J��T[��+�ꀈ�1r���D�X����K�K�i?_��k>����1���)�Ι:u�Zo�"�/����Z̛�h�k��kƌ���DYY���k��-�(����C	�� e���\~�9=ܾ+r��!`�K.�,��X��O�:|���̢3��.�`����{�cTU���O������V�
���������C��666S,DbNR?�C�d8�}��x�%�]�O<�8$��������G�*�P$3#�`�	���>��Nn������[U5�ꫯ�a��EĢ��6~��z��'��`⬗�'��[-����e˖��_�d�M7�"QUg7�5ő�� ,���p�� ���`�7��g�����¶-�r�ƕ��p^0h�#����!�lb���5P�[���
.Z���BU��__�;o�T̉�bga$X <�
v��C��_*P5#�ٸ �u�N������t�>q�0�����W�c�Ɵ��w3�� �V����1A1��⯸7"' .�z��>o1;�͛7���p1�p��o� ��$8���#����[����5-���*�cn?d��3bѓS��*՘q�Ry�Ş@{?����է��@�a���T�#��3dFFP���͜ݝ]�����BC%�^����m�6��<e�$6�R,DG`�'I7��jJ���U2�i��C�==������o��۶o�O�����|l`<2�Dz$I��I
97�T�^��f����*?���˯�U���`��~x��p%9��#++C��[j��6��#G��Z	;������_\�zu4�=�<I�x`�ũ�*���eD�' 9�
�F�&ÿcǞ��b�-]�433�1�H��_$*3��#FV1�hn��3�I�Ƌ����Q�,K��Mt��Bs��-���}���W�Z��+`��J�U�'�*29Ɔ<���֜lD 3�駟_w�u��r�`����H��I��C]1$�\4\|���F��RVV�r��aڙ��ɡ:�P�������Çc�^�����v�uk�5f�"�����@���X�7�x��w�{�٧g̘,;x�`�I=&�i#�����E�H03�	�.�Г�)��>����`���tR���
}=xޜ����E� Dh���5V^HK)V[�W�^��;�$����4�p�?�f���� X�j�������SҮ����ϝ��_��C>LsZZJ,�kn�g	U�隷��e�-C�B�uzc���t����T���%|�Ռ>Z
w}����`��#���Ԓb�����M�'�-�D��h����Z�̪�Y����A��^o��b�RV��pa{��x햢�����������:�y��a�m�}:�#3�غ{�
�^qu�С�����X4��=�剺z�0����:l��T
}V�}��
�A�w���>r?n�9��@����+�����?=ub�ys/�=�α���p�N?�����ZJ���z�lp��rs*���l��?��Sii.0��z��Ս�3�O�*�������]wGըQ��j���J�pD�%b���ٛ��%�NY�;������]�ׯ^��VU��x���p�qÆG}����ϡ#��.�	+�rza?��d6A�45�t�w>��Z�x�,���ɋ��5T����1�,M-�d�����U�u{jj�m��~Ӎ�,�{�����f�ݖ�y����OIK�hkƊ�<�{�H�$<�؊<�c��#FT��~���{����9��$����G��2�������g�f����x���|���_�^���2�r��A^6�7H��Z��+
a�1b����59q������ה��T�q��"�M�+� ���A%j�i� �v�a޼9�ݵ�e�����s� YgMp���?�;///+���9�:Qɕ�ꃧȩK�5�j��o������4�"(��p�lI�E}�}N��Q�^g�y}�P<ő�Pj��H��=�l��5a��;�uz��z��^����A�?Mħ)%"�W�%^5P>Lu�tp\���𳍐����nNdQ�;Є�J9�o�)�i���>�8����LGCJ%|8:W
��|&���ꐄ���]���_~���kS������d\٧�YS[STX�P�^z�/֬� &c盆��^t�I�Q���s�%������/1��4\��{�����{�g����yǰ=P͂�;(�"��/��*Ud:�XH���u_}�|Y�~\��bĊ�R�QQ9П[��*z��I��<����|�����g�ٰap��_n�Y '}}.^r����f%?[�yS������	6jUi���0�X;��S:f�YB���Ͽ��˘���|a5}�ׁ�������LIĆ�+O���hp�~��\�hѢK/��%��P�(/��XC�1K���g�W���l}�m�.S
�ػO!:�A���>�𩧞�ύ�5jF�yy`�ov����pD-�=_�����@�VJ/�~XS> �<xW�����UUU+W�.�?q�E%�D��3��qC�;�T\R)��;묳�
����4���+�h�� �4������Ձ���4�}���;��p����'�@/\-7'���b-�&ĸ'P&��ˮY������v��m��2��Y�L��aA#T��7ZDĎ���>3!E)A#�<y
DfǶ��}��Ɛ���\*Q���� ���M�0���]|啳�.�3gNfNMKGd��t�8d��Q�#��҂�*�u���o�e��͛��P����������a$li��dZ�ck�ps5
���ge��$[imjz���D�L*'O�q-1o�R�\v�B�Cح�.�p@������D`9�81�FC)�x��}��.������E�2.�&%0�߃�Ν;w����h���W�,����b}�I��x�Q�K���d��������C��J
E��\���"|��Ͽ��|��G���Z�&'"�}�'
j�eб�23(l߶--�1����W_��,��b�%�gf�۶qN	�qmڴ	�����z��g��޵Kn�Z><��bO�����ɝ�������~��f����/-v(���d��KN�7�q�Æ�^�|9ѱ�ͽ}nQ��Ofටe��Hd�Ν�j��{֔�_}�{+q���TN��,��Hs�� ������>��)�Fy}�+���T�Ź��Qow'F���3v�8HBg[ۓO<�nݺ��t �/���믿����M�4n\.6��@�XIlL�]ܷ����g�Cq�Tۼ�t�6~���55�G���R*��]���pB�j��4{���9s^4Fa�ں���v�XAAlzZ+|�m�r�������v`,�$az9��˚�������p�9�X�)
���Ǆ�{���ig�[��\ę�1G²D\
�J��@�BF�N☄�a������)���L�|���wn��zƈ*�i��"T��Q��m���#���N �.*�\���/�����a�)m}�!h����\Ȉ�c#Lk�z����dU))}�/2���A�en\H'	8�$��������c�z.���?]��O���g���C���)�$(�`+���ywW�@Z칃��^xᅖ����Ϡ�K�\�Uö{�]Ԫ�� ש����b�*H���K$��>btMM͞��޼y��ŋg�<���t�b2���2�f�����)332-��D�^>Y�E.!����C���'�����X"q$�-���գ�B]P��%`�].��K����v���:td��}pm+*ʁ���V"L��&Sh
j ��U��n��G�d�
��Ŗ�#���/<�ҿ��[��6�j�O������)�<iW1��(+���裏֭�7 �4HJ�8	2��"v��͆��Nz[�nŷQi�ă��6*.�G��QJQM����:�N9Ю����g��� �%�e�����uZ6|gG7>I3?���$Y ��qkժ��ޚϾ8zh��\y啥Ut���n�c�{z�wn���@ex�S�]iY�g͚?f�g��
 $�B
G���Mf�L&�tv[(� �➾.l?)�2�BR���a떟��,�Q�Щ��?'!�+d�H�@�����R�nO	�j)r�E�m��SñW\��t(���0�e���̬<��IdJeK����IVd�,���/���;�K�Ĝ.�d�%Xp<WGW����E�0N�����SP�3�H����X"�����]�6�g�X�JY������|�	��ې��ά��ʦ��ew��`��!�gh�D.QQ^PT0�رcr���uC*�����M-����@���kkz��2#!Yc�)l�sν���s%�����K�B$7�ҩ��'w$D�a{�nQ����e:��x�e�ռ܌3����]:�@�[[T�Ȩa�����s�������>Z^^������pcJ������8�D@F8 �������c/����/<����� #�M��ڏ=:��e˖�R_4���Z��'S��f$������S�Z�歷]c�����_������U��>����N�ݞΚ�Z��>i\UCC��)��upsf��������x������$E�
�=x� o��e�7ot��{Ǎ�b�'i5*�-5�%�&9%�;n�>cF09t�z�G��Eޞ�V���Z�)���(��2)�ww}����E[���
{:�O	l��7����UO����qI4\��g,5=O����`>C1׉�f̹-���;ٷg# �Q'OOϖ��-�qD	��ƃ��.��>}Ƅs�;�1�<p4��%e�˧�%l)��.j��H1��:�Rr<P��))�
�K� d�:��ЇĹ���A���#�d�!�nN���#q�H�8\T��ʽ�t�����m��s�I�`���j�X����H�
pge܉����:�
�
����}w�;���B+�@�R%;�|�ç�[4mm���`�;\�U3mڴ��vX>�R���DR��c��EE� *�4�~.������>��	<>�����	{	���7.��
�#N7��\��}�����_��ʨ��ܽs��7�1�T�a��=@�*�j��ԓCp�kT��9�Ϛ�AN��b�P��$3�< 0�z��a��~�8�]�6U�,e+�\&��w{��)!�Lgc^Z�фm�m'O�
��4�ټe3<f�sfZ.l3nĔ����	��H620O+3�.^�7Щ�&�DoȂl<��s_}��M7ݴd��$��O�5�����G\��I��2�����̎[����۷;�ܣG�r���M�m�>���ظ;5'o����s4t�����gϞY�f]z�DYT�L[��[�T��{��!�I�s?!]��aZp�&������KP=��E�=�}�e�`���fѱ�͆�B��«����%�9���=�V�����/��S%�^�&�9�E����҂Z[��fjZ
q�8lJ����b.�+��X9.^-�]gU2��d��io�l�;�
�0$G��'Jd5��I���)�0������������2��7�q��h4I�𺺝�(~F|[�U{p������R���}��;�:���6E�ק���q�7�<$:K;���+߂�:�&
�ROg7�sIb�2�̘�&��>�E�˯�9sfaQ�J�Ž��[�I~ ��� 3�ةU$K��W`@���7�g�<s��?I�����E���0p�7�P#� ��L":���2���ѻ��رC�\��#��".&L���۠?$4�����6mέ�.��[K���ܫ��v��k�I)
+�A���cF����;�]���G]���7o����4�	'�F;z�ԩz�3f ʤ���:8�:1lnH�լ/T ������c��&��!4<�Z�O�G�C��bʔ)o �i�fO������*c�k�;�s`�v��9c���ǚO>��?�)E��V�݊�h�h�'�?���/��@sss}c#Q���YRk(wC����'��ʷ������vR6�ZAQ+f��#`�1�~�̙Ж�̚;q��~j!�Q@���'�����+���=^)^۷l������"��^~_��TS׌3.�r�n��V�Y(�-yy��^߀'�LϠ�I�&AK�|�D`#&r�n�S�1�_a�Tɖ��R�����o{+K��)�8ۻO�bi!���>Gx4R4�י�n_yy��lko����Ɗr4��W��YHF�UR(�[���Ŋ]����������^*������X&�\��
$�G��u,��ENi����D���	�"�n��x	�/�Z&�'a�J�#檔�C��$ٰ\dt��>8QB���r�\iI.�
R\T�-ۯ��z�Xl�L&�"�%�Oq)|������o޷o����d<JK�9V/�_��.S3��O�*�s�(�x��H8�qiqT������䒑��9���������3g��fU)� �q��*�1�@��pP�ڸ��6�0(���pݒ���k�L��z��ӾDnD ֔�r
��MBɻ��q~%� �E��BJ���Dª��)J8���߰�W�|kĈ�ͳ̈V�fqH ��8=�� 
5��z�`;��{���~衇#�R3�d�Yy��v8���<���������;�0����I�`�	ӏEd���a��n����z�K�ऌ����Jh ,��kk���6�3�G�JN( ��І��{��j�*�
�wȐJLHww�@G���HOό�HH��׸Io��}�FJ�L�0\�A�HxXUe8�@�~���_����s,��(F=]�ʆB���>��Ok���A��h�Y�>Gw}BWjSN�4j(E|����8��Ἔ��3���w^߰a��\[Yaz�G�u��ő����`�1Y4D'�+�*�N�'`�HQ&�JɯQ��MI����򗿌�8Ӑ�p��55��b����P����F+$����/�n��6j�������O�f�c>���`1��:I�p<tS��̐�8~\f6q���}̭��9q���8;pvw82�v+!U"�(����a�x\�P,,l�ڬ&E������?a�eW\!)��q�tz�}}�U0�H���%e�6�`~�R�>��K`S������.:H̸q�����{��q���hԍ;
K���/�|���6���b��}a_��� F�^�<���k�U�U99�G#3ӹ�w>\����w/��Ά�Z>�͡�����p��ފ=��kSSSǌ��/�=��>1r�_�+P��Pw�۪��{���2�z�S�3����Yˊ��TG��<p���a����5Ǡ�FeG[]J���^T�;��\���O;��у���;4c�E.OK�L�8��]m�r�G�I|ᠿ�棤j�m;1o�^�/y��������Re��)�-Z�������St���A?�7�}Vv�h3�T���S�
���嗍��jlc��@�6�(����R(ti��ؕ��ݹ���5�r��ˊ����m0��h�Q�Rg2;��T)�++��|N:�O&����O��.���Ԝl��)[x��UU�L���Q�����)(��Le��ȣ��Ѻ�}���v�I5��ə�4LlNP2�8h�Q�u�/�*�)b�ʝ�����'�	܅�
cQ���R+�C�gr~����`���00/>gX���0{�p�O�P8�E4
���dTE�n4���xhX:dM�Nu����E<G��^���۶�:x�����թP���<w\E�֑9�1A=�+'�$�V���tm��=��*�۪r)������j<�u�]�r��'�xb�ԩx�c��i��dl��h��n�	l�����
T(S�FǑp4ٯIE�}QN��bi��+�r�6���'���p��8�dt��	c���k�;��9{��Z�V���~o8L�{a30��}�--D�?i���裏���:x.>Q�s9 ���87ɺ����I��"�45B;��x�6�E����  %��X�;~)��ҥ̝��.��FM6Ģ��>�����S��#�J�3���2�oX����a5�}���Eo1|����\ѿ|x��L��~&^P
���*5�/|�+by�a��Iܑx�[[�#%�h����hq��7>��3-���y�T�%Z��q ��D{1�Y�O�0��&�
�J�#W+U�L�j��C=�f͚��X�Ք�֊�?D%������d 8�`\����`���1ڊ!�z�a����x{�נG���^b�Q�8��)�<y?Q(pƢ�(��s�
����&����X�|����o��ք�j�d��b��of�3jԨM�l���Fz"q�gg��c4�L�.���y�Z ���Fl�{G�3q�3��y�l�'NՔ?����4 �Y���,��\5j�x�T|�"���oL�9M'� ��ԓ"���#���S-�1������"M`�������1��ډ{@N���9߅a�M�����j�
�)���oߡn����e���t��H��=��sUL����˯�0�ּy�����������(s>��	O�"�\MK��1��P4��گ�x�!%�Ç�z�������Z�tQ�>��W�#X���V�l���޲eˡ�5�sΜ�sMVk��r��q���@��I~�\�9��ܘ�M��`�z��;�lٳ}+����3p/��HiLmm@Ղ�C���z	��T�k�u4͟?��]�۪�*�"E N	[�$s�`�3�0`A�1����_|�%�Ɍ:�ش�8���ڨ�U&z$�:�ֺ�Ęk�v��͟�G]�Ï���_\V^.�RN�<|�����v3y�Z�"������!����j��/8z'�#�J k�-��'n.�D=��"�y�$�$���j�\7���JAΆ]�T�r�>�_Y}n��t7>��r��-[�#Q��������d�#�=~ٶ��10����R[]}���N�E�=���z���2S��"]�':[S6e�7
DH�ig��a]k�	�ו���DP��k���,�'"j��r箦"�DMk�N����CJ�>�F���Pʃ��`�J�/)��A�pD������S;;�
�MF ��M�6������z ZkjnIMM?p����.�-�ˇ��ھ>� h�|S΃��[8���̐f�1P=��W4��pS;�O`����r8�
%�٤6t��<Oȥ�����M�4�G?~�,���EDC�hX�I!�:p|�����}�.���v�je����`&�>��P0���x
�$�<�}q:�VG0E�w��p�,/��D(ĳF1�"��Y5J��W�~��o��{��l�V�>�m�*�u:���R�<i2�y����|�I�PzZ�Z��y������/��Y�0�p$*�Z�
S@*&AF�����3��MJ��h�]����}��'˖�{�=�`�l����`���Ä���h��k�5`B�(����W�^�7'L���?��v�Z)Ku�)K������R.��dP�%��`�g��TjJq ��>��+������Y��`WO�F��R�G���YP����//��r(�x�/����Ty���>oCC���R�����������&h�9�������3�T���X>��p�d�F�m>�U:I��U���G�(�x�D}iT���K	n*u�#
T������KI_�����Ċ�>;yrn�>ۀQ95:�##B����������(u]}]eťD-��>0[�M��XU��?w�>u6�f�^ʓ2�E\�#��:�Ы�o�Э>����)Q���f�<�!$k"���D)����{[�_y�<�����G���Y��v�fYdW3f#{p�����ܼA�A�Kȩ�� �]��)��0Sf�"�t���9sD���u��9J@�J�SO�EW���I����cqIe����@XM襄O.S)RzZJ<�X��@ E��}��?��C���3ƊE�bT*����8��X�D�fWg�[��c����̖.�s���̴T��#��:�,|+��sStݡ���_�}��7�8�mg�-�@L��T`$���c
=&3��r$�'�puR�%�W�t{䂣IRĢ	���?�|tw����m����ʳ�
�ˊ
[�꺽T�y�:!]�Q��ꩯ��V�~�\ ��}G������J����#F'���L�N[[G���'Lȵ����o�?2|�0�u:����>�7	�Yt:xfq�D�Ԣ�]��ģ}J�oڤ�֖�/�3|��k�P����x����,�_	U��vwz�
��ih��Na/�[���������^_WW=�.f/--��1{z�Ξ݌G��A0��F�A(9.��v��#��M=V���,�tЙ���ׁa����>|QRF��ON�h�@�Č�Rӟ����ի��ꏟ<����'O��Ke��o�֠�_�Q}}�.��~��c���7 ?9���mE
�"���d�@��=y.+�ȹר������t
��#GN�0؟��=�`r�=�	,'�����?C�H�"?�<��A�)��9q�{'����1�,|<Ϲ-�����ܞ����MC"XM��i��C~R���L�B�����C���ec!^z���g�eq��0��ߩGֆw�y'�R܆G%���P"B�P�*���i�w���2%�f���{H�l(*�8��3񳣣��7�ܶ}�%�\��?/�%q�r�@��xaa�=��-[�i�&��TF!��sƃ4М�AqB�/�LVB&Y���l����8���L ��/@9.X�`֬YX���:lH�}�dN>�}�Ձ�����ǄCl��������!8jŮ'3]2�]�Ÿ$�S,�<��B�$��H� ����u7�|��g�S�W�l�MM&{zyy9�5��X��NCc�`nCA�������ouvz�R�.�+qDy�Qԑ��"�O�0&�,��Ơ�����������r���<2�5k��ŋn�����t��Ot��u0i��%�	x)u�Љ���5��Ē�_{��S��,Y@d>�
'�-�P�nX���)������#�b�88G��0 Z�yAѩ�W�={���~�ԩj���p�L5�-	�?���ii������Y!#��!T�[��w�L\_{�5k����,����SJ��p�u�4��5�K��(Y�+�>nSS�M7ݴp�B�ӕCG���<pxǎ)������'(��{CC�b��~��4��tEb�~ʤ��Ӂݿ|���'�����R���@�B��/@u��n�����
�n�Ņ�������q ��.:{�ر���삂Dk;���N{�I������["o�X]]��QDC�9���N���PDm˖-��Y�%�?�r�ʿ������ʙ"rε��#�NϏ&I��0A\����Vč�;5��˯�qΜ9c�O�]p���C�9߈:0��I
�lPn�H�V��c�R'��>f��;ZU<iS�a� r@�ǎK/�@����P]7� ���*GF��g�и��9����ؗr��8����=��I�8q"`����\��l��J(�&�LRp'Jx��͛���N��������f�Nof��lt�#�Z��(g��I��"�~�O���#�$I��fx`��@k�$��G�F8%�Ƿ��h�V$'(����O��;\)�$Ȟ��I�Y���x�A�r���R�Kp�B�ov"�3
����w�<�~�_a�8����'n���9{�v��ĄaR���������n�>�/����駟_{�`�#P�R)8�
R��
��Ɵ�;��L�`T���RRS4�0���Xo&��`��'��ڐ#��Pn�� �G�F�i!�pS���j�����d�����˗=�B�g�%J��J��L������aV���V.r�%N��q)����RU��=MM}��?� ���c�a���C��q��-,|����z���ǀ��g�}�ȧk�V�C�ib��˜,_SS�ʅņ��9�?&3�Ъ� �j�"�G�~"�����}%�iG�6}���G�6u꥗^:l�8�Aǳ��B^E8�p���eu ��1c:����_{�o���t��R^� �J^�Ƙ��p����פ��~*tшJ��wvQ>G�/z1��FcL��JF��(�JY4F+N]���MZ�wwm�u�x��TRGK�LaLIM���$�XL&���~���v�z�!�E��Q�E����?����H�k�9�)V�R�\aJb^���#�ͥUOhوFh�G9L%#=t!g(�;���}��j�m�Us�w�w�VVAAm���{a�tF��u��&�'�fUiԒFi��w�ڼk���3��#�}�W}��.,ha!�BgD�	�^x�~������8�$&�P(��&|~Lv\0�P����+2�dx��{v���[p���W�***lll:U{rPn��b�����}7����0'z�
����9���d��6�#Ɩ/[�ɪ�؏U*�g@���c"���`oE����@���wu�h������!���$?��j�g�`G��T��/�.�3k��I�p_�s{�{���{}�>�Z��b��	O���Q���Z����J�m�0a�#�7l����/�v�^�@fUH�-
�";�D�j�v���II�+vi����N����UVٶy�W_||��µHO1�
2��=������{�^~>[�u��p�����Ab/�S�gG&�:'1�yp}h? �"��N��{�3w�ƥpMn8�?�d�ۺ�7�L���d�'��8b���O���\?�<A�� /z�6I�����~ff�ʩS������X\@Ϟ}����tr��MZ�~�/���f�=֚(��p~c��]l����>7����n�	�Sy���
1Zd��}�9��c�X;%	Yc��I2n�kv���K��*��`	���R���+x�7-~�^���)>ɵ:aV_ (^�JX���(͢���ђ�6��Ң)��gd���)��C4��{�����@�6^�<i�Y�X�����-�7��P&$=o>k�� vu�c��Ma��(��V����fy���&0>D�d�v~���I��p*@|$���#�B$���E,{��e�����B�a�9���7ހ�����~3ncW ����>}:����ѣ9���Y9\����3Ce��,
�79�첰p2��I�l�r�EJ����������N�}�v��	��/�|+7//!���}V�L/	����cǮ���yz���))f�N���-X�$��T(�?h��nx-R8��-��L=���y�,N�T(��ƙ���0H�%1byya]]���5�w��06e|zvvk'�y{���&�ҩ�}}�'�=o�y�H`Æ��w,��|���S�(J���𧟪���`")��J�
±~.zZk�@uB�q�-�h�.��`A�"G������'\y��B�;q�ē5'����ˣ���>��{�w�a�:l��̉G�
t� �P�B�D�M"(Ğ�I��G{ϯ�Y�sK�p��bHt�-'��ీ�P:B������[��7��������%�T]+7H	d��S�� 9���C*����駞���M:t(�7an��«!�%�xZiC������ �B*���9�0�y5�"�>!QLF�m���X�1�'`w�MfQ�AeGý�J�{-.Zn�.�/Ď��q��I|����ܵ�O>���o�N5�d,4��(%}*f�`���f���`��33�UTTL�<yŊPA�.{���$gPщ'�ȱ�E7yNNn��� �EOss3+@�"S�ko���*.�P=z:w����J���A`���	&0�r�=��T���|����=��?'῵��e��`�IIe0ŭ01/iDG@�c�(��s�R�n��G$yB�}��J�\��C;�	���@�	���K�Jg<)�{�kr�VC���Sur�R��)�
�V�ߣRTG�"�;c�8����&�4`���a���.a��
qu#("`r*M� b�HI��qAo�>(�0�u������G\:6[G{{@��Q�pd���A.� #�b��~B\���'�5�`�h���'�*�$V
.�`r����-�@�&�w9�,���<Cŀ��$�I�%�}R�����/��:7���d�M�6Y�7��)&?&�������D�)�.�90��
�&-�iL��?��B:-*p��m{Vk�A4��3	�I��uu�ׯ���kE��fIP���P(�a��%%%EE%�dT���grM��v��������y:g~�g�(�G&�5
�
IR�5��	�>�HB�R�Y|{}nn�F�����ˊͻ�ڶ��8q�ZZ�"��ȑ#z`T[Ow��f4�5C�'���!H�w��1�1=yH�N�RDUA_<J&����j�Z� ���4Z���5'�Ыh/ <h�~�,��Z��(ߚ���{�����=v��.s�h�lShT�������[g�B�._������[0xT�`�ۭ�ǃC�Z�N�x�Jn0�ԅ1�E��Uj` �J��'DD=�\qy�LX(�jE8��*D�pT�	huZ:,�(�Dhft�վ����,��
����p��=�Fb�TiS��zCc��)�GY���}�󆯨�C��lD���F�ҋ��0�Fd	Q9-;��'�S(���O�"N�t-��C��H���A��GTİyV����~��;v,\��..��cG�df8 �R\��H���y ����SE���vÆ���딥����&�V���p�b�{���<"R\�`,��lsY8���-s5�%a�Up�,/���3�SmkzJV}s+X�����7�=cz�Q6K>�m��$�4*�^�ҀR!�<���VX������Z�t����t����%$��b�
����hq�+":�;k����z�
o�FO'���S<���fL����K�(_�Ҫ�\��v��)%�����eJ�n7,�.:eT �z��Z@��3[�?����{�n�i͚5�g��ٸq#�}2���XE�IT�f�ƭ�9я۟�A�%��b���ix�[�nť*���Ok�_Y}����?)~�d����
(nC(W���P6���^,rs����o���:�hҫ?	_)���y4���R>�mH:|lzEj�;\QƩ�;`+ŧe\q�N?{fI�!��e�̂d�7�[!�?�K�mOʎ/?]2��aa�Qg5�������A��W}�w�wߒ/�̪�ں����j-��e�I	L`d36�=a(b�!��A0K��㰬 �
�	؎{��gF���F�^�n�z��5�*�̷�u~������̒�Y/_�w﷜���w� sa#�T�t���LhB��2U���A���'Ap�� �[L�̙�4-�kZ���S�,*݂R\�&�T���f��!l� t��U�w�"��{�	I_U^S�'36$_dg�aF�lbڄ�佩i!\y���h���C5���։�t����D���\�&I�	�dkKz�`������v+�y���*4��F��#��R��̸�n����"x�Ռd�@"2���tCIօ�{pp�R��x����{�7�3/��7�71���9���w�R�0�KM��rL;���MR�:uD�ů�]e�c9�Z���~����*-����?,4��|�3?������(hmcM��q�'�|r�7�������D�&k�Ȯ+�̕m�g��5��*��s%����T��*�:jJ-b�Tq e��P����83������k?�7���w�:.`�]y�qRv�]�~����3��Xm�� xm�j�I�a_�n���Q��VZ�����J�o�c֑6q��00�p;;{� {�4v���n������|�������?��{�?���$��Fu�K ?eP�ǯ\�~���_��?��S'��p�#b����tō���%.�˲	K��p��"��Շݙ� 6I�U�	�T�{�9��ʒ��1�W^y�������O���Z��76�����+X=��� e����?���	��x�3͐�){��&7ϘD�s�����o��6��R�d�g�#}w>��Bj��_��?�C?���;k'׆�/c��N)�p��/,�O|��g�z����?��_�Ņ�k��<!|c�?��?�]x���{��<��#ؠ��~���؃ K�7q��F����
L��(3aX�'�ꧬ3���-I}�l%^~X=��8��E<I��C��LF��F=�Qnnn���AW͋�ޗ�H��#r��"[͏<�n����w�թ��z�w)�K��L+Mr����n1�N�^��>4_��cHss]	I\M:�����6��U�#Z�o0�B��D����b��G/����a��1o>I٠P*'�Q����S�n҅�y����P��;��,O&���ivD]$��������{H衮tJ|�ڕ��#s�بZ��a~n�ytx����o1�8f:G/�F�5ߤ����T}��TU$�`���`/"ڲ��h�� ���e���=���7�R�qM�~*=���ׯ��Kb�|�FX⤣�A}S��2�����������/���%��B*4�T��z����x�w�����uB��R@�u��u�V��V�������=g��.��V�=ٺ�N݅�` �����^j��-��@w�e�׼��~5RE��RQ�ێ�oH|�?�^�H�^d���ȳS�&^1Qj�hK���#!��n@r++����`�ĉQ76��hqy�`sg8�4	$I'?|酗�Z�c��6Bg4��>؝;��I_�t��L$9�;)�	hL>Ѱ]/�B_�y5*'��/W�7j��yC}�FA3ϝn.ߊ�|<پ�x���I)���n���G����ʯ��,M���ݭ�Vo^{���wy�������/���?<���v�0	d5�<��_Z�����3N7������M���H<�M\���Y�����I� 犥Sѥ�.*�Kz�����ěo����^�m� Z<����3{[��c�1�y������7~��������'�ŋ��y����ܽub�y���4���T.�}��)vE��I�e¹=�`�g|�GP�C�I҈����nK����z���;�z�ƓO<����q�͗������������y���D��斮ݺ��;����A-����w~�~��G?�����bl�� �$M�Hz��|�{40�K�3
q�y��H�2�'7�D�nůy��/���H��L{&��yE��������<���7�����/��3O
"�7A���F�����Ɔ�>�w�R,2�����L��d� {s����ƌ|�ApBr�4����[hO����[ke�#�g�$:�L ɤ��0O���w?p�ؾU�O�����HJ�j7_���1LU:-*��r8�;Y�e�4n�6u\˦�<�țe��)1�-5���%�=L�
�J���_��@/���]LQj���d�,y�(��iu�
iEc,�d��L{r���%.H?���Q��DF�	ԐK���	��*�i2Ԭ�s��&4*Sy{�'� -��3��z�\���}��ڵk7Ο?{��9fMc���)�0��[7%+S��Z�͍/\cs/*{���CܙݲI�tx���+v|Nht:3�Mp~#��;���%�;��o�=j%=+t)�*��`�}i��/
�J}'z}��!+2�i�>��Be�� �Y,��������J�-M�-*l`�DQ%ic��\�"�6��;s�>x{
�?�L��ٞ���DR�����.�-�A�%&rjEp���!6>��vv|��47�/"~(f��P��[���F�PhcuՕ
P��3Mn)�/�a���6��c0��?DA�a� ܸ������,8��ʊX����7v��fƥf,v��b.�t�J��s舞�JcSyn�(��r_HB&�d���}����wã1߃8����K�	قe+�J6�u��mg�S�!���!8`N9�6��(��8a��'����7'�lWO�vQ�0'p���1����goݺ�^�xq�H�jQ�گ��Π҉(�RnCGU[A(	���a�������W�� �C�:��'�-�q_:P����^��&;��ݘ~�~��G���'�0�=�8��׿����3���?����?�~gV�?`���ظŅE5�J�+�,uSSJ��ӠbVe��4����n���� ���D�D�(��lw��g�y8���'?�������|�w�X��b�xF�cuc�����������{�޽K(�h,�$�;_�v4��idp��J��U.&(�1hc�ب��J���2t�T�e^�4��>#-PR<�D/����\KG�	���f*W�<&IY|�K��^xAN�9 ��o�q��=�������LƱr��۝k�:҉�rb����L�E�	�>�H�^X�Y�׏���B����B�cЁ���*��Ξ=�C��	v�	&~���ͅ:qC.��^�̖��!
lml�g�i,F��r��S�0�ס	./.�MIC�P�,� �q�^1 �ub��)D�h���F�[Q6�ⱤzHۗ��pԇ����
�ҕ��3q��I#�$]
uBQR���V3���ZK)f���uj+
-~��p;I�5�v�4(��a����=O�l'c�<�w&I�
zb���In+�#,MZ�
mw�v�So5f+�L��zZ9�>�ZN�j@��D�;�J_Z���J۠���}wX�j-{>�#s�ymmM�x+�b��+����q��|�Ņ2���jt|�by���a��I rh2ɓv���`x���g�(D�Sx�d��Y	�S+�f���F���J8,P�d�ڽ;���YG��a<<��d���
���ⶢӤ��i`#\�=�م&4
���w�N��lD.�V�D~�q�N؈L�yNz~e�ը6V3ͳ��̅��^�~}f��޼�dIi��pg��A]�}!*�ɳf�'�z��0peL6��}��:���������Z�$��[�7�*�'>�(������$@�|�`��:o��4��K�$=F2 �]x�����O�l%�!��Ѱo�A.Q1/�ƞ)�����*5�>)�r�ę)m����� BI�nF���Ή*�j۔�2�D邁?k�x�Qk2�4�=?;s��U����am��5�*5�	�jA;�tZ���@?������$a�O��1rG�H��G���=e���T�c�K+��^�޲�㏆C��_}�k��O��w�9u:phh��+ۛ[Ln�	~g~����~��[�_r�	������=yB�T�}xtWf��ujfFP�f���Y�N�0�#�i�Y>��m&�&��I6ɍ������0�7e�#����O|�~�����g������%��co�Y׬����pH��Ź�9���8����bGh��5��;�`̬S�CAՒ�Y��^��@��)�>��q�
|
���R�%~�p�M�����%<�3��!�[ة�O�w����U�'�(gne!e*�Fƨ<���^��Ap���y5U�gU�VQe����MM1v���me �t������6���t$�y��������,��WY�^�0�>���G�����[Q�t|ߎ��'_wY��lы���m�>�C���Y�U����T^��ܪ8Ď����w�Ӊ��ko��G��_?�[����.sX�[�ح��a��
L��#:�|�5����	�υ�=�0jA���2�&�'"���f�J����o�E�˨�I��F�(��&�V]��a4K��/Imq��u�9*RJ�Nh������.�iYX[�ϑ0J}=�u��#g�(󒃦i�P����3����5wLUy�x"��f�f����w��b��5��[�76z
�uI�q�o*��;
,!���R�up�E�,�y��!�	����FЙ'/�Gw��B;�N`>3,
��i�J@*��,na��d??l����.�3e`u�/�Ǻ��/)5r:DI���-����Y��Ν�0���`<�D0j�*��.�k+�Q�����[2l�4�(�2�ɭRȍ��f�績�Nm�-�'�������[����)S�XS��jɋҎ�z�{w����0����A�?��C�v�ó�>���
:�̴KK�%�q�F�	zN���dD���Ź�Gk�+�����6��s��מ!?!��6��޻w�V����OH���nw���I�7t<��Cws$��ګ�P�K�/l8�PGt����S(:fk�σV�I�AYS��50���^���__ET��B��!�e�ǘF��i���`�kIIt�$8���v�r�+�)�D�E�
������K����.�Ĺj�o�QQ�|~�ÂxE�iDSH�<V� ���o�>gj�(ˏ��1�̐N��9����Gh��{��GF~~_���!<"��h�R��U�#61��އ����À�4_�.��_��}�*R�Ɓ��=�7❃�>��ڇ��w�z��F��;+4��� ����i��IV���HX�R�m����L�K�uf������^"�zB� �$)�m5�F\�R+��P�tB_36L8�+X����� ִ>Oܶ�ѣx���s�7�R�$���H}��G�:P&<l�0�C�:lP��ԛ!�Vē"�/nhBO薐;�C֬dƅ��ɸ~VT�I|wX2���Y���Z��֡ȅ���VMɋL���;+Q~h�8��VER/$��E���vӂ|������=�AԐ�l�Ĥ��RNs��0M4VB7��jy�v����Rވ3̊')&(M։'����;�V-< �zxF����& k�o�|R_C&��ً�x���h��x'O� ef���;�Ok�R]l��+WɁ��sMt��%�R���ҏ)W�|I�]��V�c�
�Y!T�kf�{0�|�O���>���E���nԄ\�|)�pvW�(wkw2��|$}��u��//�h�*ca&A]�B��1S�����{�����(&�nNQ�o\]~.S
���L?sM�C��f+��������F�On^�Qd��K��!��^ ���/�����O?�]�Ɵ� 0JqTو���8�W�\�y�����	���Ԫ�Θ�/�-����~����<�ދǵ�oG�U�U��K��r[Ʊ��&IΜ��$�TF
���7j�fUi�����Ji���Y��6���"��t(��kJ-:��%X,�߼�LUs4u���%�V�`��:2REaAO�[���QfZ�k�i��}�s8�����F��
$�G�����kU\7�fJ�Y��[*��QԎ+ߤ�U���簕�V%�z��W�����h�\}�탎|�)�!r;G+������MM6;5������T����8.�koNi+R|��W���SGՑ�����q{O�BWf7~8�\j��5$Gi�J-�U���4�P�Qy(�l��u<�)�=�`v��YY�'�����&D�+)*}f5/H^7���N�D��ƔGq��BK �x뭷�<��-韰��W@[�i���fZM�x{�'���D>���w��XMWsHl�	+`��[)iUʧ1�ZlT��Ф#�t�Xu��J6��,�e%��Gm}{&yI@�݉5-���y���Ӫ�<��
*���u�ٸi���"�Pa��3�ON�ԙ[���B�R�j�Fj�.o^���d_�^��'��!djn]4�@�oc��^�-4��
���Ph"3�gPvߙ��(Q����,����kɖ���\(H7�We ��IäM�2�b�4.���O��G���_��W !��y��I����W_y��ٳ[[[l���{'O�\__���qC��9��iv�4b��JF�7�qƿ �ϵ���p��:L	��UV�:�g�={���S�~�qoK�\Ǘ��?��t�D!���~^��{nnA���J9����s]Ќfj�$/�1ũ��p+,h���e��Q�ۇ���u-���)�2`$�Co��g���G�������d���%L<�$P�q��U�xԹ]S�<+�]i��&(�����؅�!��׫z�U��}D���5���k�#���E����&W�[p���K��Rf�,��z]q9"�w������Oj]� 7�FHߩU��aQd*@'G�0 �:ypxR\M���Q��0�U$��1�����"��W(�OIЊ�b�������퀟d�ѝO
u 	��!��H��8�'�E�I��*Yo��&ʙ�П4��k@N�A�7<WPg[�ԡ80F�Τb�w`uf:��<]n���|��p��-׈��Q�
�3���-����j��]]>љ��E�0A��a*hR�����T�v��2�����C�Z����xSi��ғ�Q�r�u���)xDa��Qw���#�����~?��,�Q��<��d4���
\O�Ƀ	�ʡD�Nc4�*���L�GT�=���2��Q.��d,Yc�]��0�8l4[��i��O&iY�L���dr��8jw�F$�^Н[��|�om�>p�<V:�Un*�㹩 �R������7�>5R�Q��ץ�$S�(ˠZ	>l�����(�}�I�F�[\��IO����vg�wF˫�.I����[��n)8�|:�k����9K���Tp!�%��%���l�ĉŨ������!�Z0�0��%��l@:�9��0n�n<G7�t���E \)�c�~3��h�]i���$�J���*��Yϼ������P�|���3*7f�$�LT`�vmm��/�Ӗ�[�"�%j�i�dqP �wP�r~�mU�G^vN�i߆�_Ԥ~*-���#�����4�Z\̋>]p6��xP�2J~�qshII"�$����/���&������4�	|�����]���*M._[��T�9nL3��HN]�k�S��l����o�����*FUTE1-������TA>�-�ky�y>MO�)f�A|43���e��3��(u��V.-f�Vi;ݗN�a�S��r�������y��3GD{�W�;�ԧi��N{�O��[KF�* A�J�r�w�̰�cO�Ǻ�H?l�D��P�ô��Ur:>S&�2 ���������q�tH^D���g�y��|� �D5�-�e8���5s��ݻ���j��e��yo�.]eK����
��1�g*gش��� �Y��o>���ZIE����_!0fZW����� lRN���GH�^�T?e���S݁�Xnv8��Q�@~��QI��8:R_�̢rD�85���>�<w�h'9��SsD�W0eU�!'bb6{Uڼ㖘��M�5����S�d˱����A4�3hG~���T?�|��Of�C��\Hީ�K�{���G@c��F-���W���;�||��-|$A�-���Y�)�3����ơ�t��V�1	�%�����K� �t�A��S�A��3Xy��D���a��6=F��/}�ג}H�'�|�7���������Ǐ>�4�ӧO����0��u�8T��eCz���0CNg\�Tl7y�ᇯ]�Vc���%�k� �ь�I:с6����`�gff[�N��)D���㓩@:A���3�� jV*|9�R
{���&��2-S�p�%���p3dt@�{�������г�ܕkαB�
QZ�̺��e���뮮w�N�+��q�o��>�P��z�N-;�l
��<`�W�2Ġ��,Z�����_#�a��0a �9*B��S��U����O-~�����'��6�T<�r|�a-��x�ͺe��O��sL�5����V�p�˫Q�)��I^Y�#�d���R@C��F�F��nAH�W��x��@�onl���'��g.��]2=T
�ơPJ��p��#��CQ�D����<�'c=�3�+��.\yR�	ݼ;�܁�bO��������-U�1�\2 �{]��i�;��:��!{\�����PV��Ú��������N��V�6�
�J�z���`�g��97���Wŧ�9�*/�r�����q�1Օ�*Wû��9���V���`F�Ƭ=1�a���O��6���-4����0f�N��VY(�]�Ų��4�Sz�K�ꪰ1����d���TJ`$�Ő1�I�@�@i�T2��l5hHw��p�&��3�Ę>�l睮v)���/��G}u������R��LK\��d��O=�q"��|�W|���OZQ��d�����|����v._^�����	B�G�'^���t��A�t�~��Z� 9btR!ܝ����t��qu7�$��>���t��g�����-2�o�����z�����w�U:d�4�	�ǩ������X;wZ�h�+���hi��=���F�Q�@?��������W��={�O�'oܸq��e��߾}����˴ɓ��R]f�w瘕UTQi��z/�����FR�W�/��Ö�q����>Q��"-�-�*�+��L�T�:�Yq��~w5�M��=��d5e��ej(��=䙄��*߆I�f���?��Q?V����Lr��wmVU��Za�񵢯&��E����Y���-�)Tz��ʫ���ק����s,#�
3�F��葟���g}�*{�T������H;�FW~, |�;ԧ_S~-���;0�+l��Z>�T
�+�1(��#w.*�}�[��gU�s���I�ǵ
���!�׻��DyuL]k�=i9m铢���3��Zz�V�x��0���y@�?��/��G�
(K�ۍ�IX�U�`=�q��5<g�yS�\�r�_��4a�w��]SAt���kY������VLGh��)�gǭ��-K�6���Zƻ��-3
�s��@����,Y����
Ji8�c��[u��:B�EU�9T�8�khZ���T�@�X�Lԅ��ۋ?f\:�,>w�8��#���b��*_d���9�͆f��F�p����тlzR"/4��_ �W;����4Ua�N�c�E"�Q��mD��z�p5��a����S��ה*��0�Uf�#Xm���#b��`����/�y"��O��A�0�766���	�m �륗^�D�W���_i������t��zڋ5�B���ۻz��c�=v_��ͤ�=$bV��F�E�(b�yw_��h�����,���Lw�@�&��z�y���y�O�iJ�L2�k*p8�I��x����(X�X����/��7�	���tR$A10��fk8�]�I���0�x�uRJW�-���i|Dp�2���톝�H�*W�>xj�~��6�(j�N�LG�
��&�`��c�����1�>B۝>4����&̝I��q�k6�!���:�̴�3��dq�Zi���v��P��/�U)�1�W423өSfų����]PW�F��.8�����>�)�0�u��:=6JQ��&��YBf"�,8/�-�qTY��� ��Jœ,�v�3N�.�!�Q�.	Z�7\a[�;�H��S�L�ҩl.*�׸5�	����^�� ��Vh���,�'i3�.�Fvh����e� 6��^�/M2Xxm�>51ذBj�5|HO�uOq��G۲x ,ҽugcnq�C�J1�o�l2Jz�^�	��@L���o?��N�I�I8�F�
$�V����ww�$���F���33�r�� ۿ3����M�Fg��w}�I�-�8k�'Vf��`�i�$��0(�q�߻���l��q��0����&�8�<kŸ�y'q�uNZ8��x�?i��{ݳ��z�E�PG�msu���Jјs�������Vݎ�O�v�`(а�+���I*1N�8�Z=�h�L6c�7��q*A�)�YM��e6Pn 5~3S+&[�����`���S�'*W�a�6���q�����N��u�33��&;٨�ۙ�.�"���5�gtogpw�w p��ag�����J�8��h��t��y�T�E54T�D#�z6M;�$�P�҉�VUb8�J��a��m�18��l-M\���7�� lz�?JFi��͵�����CR�@��ɓ��m㇩#f6T8��eM��6�
��	���x,�b3/�q�B����4�u��y�-wè��K�ɺ�s��_����<{j�dP�q��n�h{{��鳧&���7rO����&�ް/N��@d���m�"�����Or-`�x0�n��4iO�&0-h�.�и�$��i���uAE�I%+)מ�N����h���`��w3#8oRN��4돓م٥ե��f<:�f��|q�{=A�͋���� ?�!eĊ~V"5A�_�x/��C=�~W� ��~�m��`���֠:J�h`R�|��B ��-X٣�^:�d�<��{�����@_w���·Y�D���{K���U�Vs蜪�Y|S�%n�k���r+<�I�ط�`��72�� ][2�#�WQ�ի���|�7��L˾R�AkS�мU^ks�آ�(5�H��Xl��������*T�4i����H˟�Ħ>`U��ȥ��Ig_��3Z��7��j� ����>K��2��Y[s�~������kxV���8��Ub�qs�~-ѡ>�#����t��N]; �wE-:p$_��u���&�E�.S�&j{Y2�g��e=/4D��*j�~S�h����\p!�	̦�=1�'�ۈ�#��Yn��I[P�y��Hҵ��T�b��hz$uX��6�ܼ9���sw]{�
����KK$g�w�m_1�]`�ez �Dlb��2�\�d�� ��Ը�#�����~'�!!v��S�+�	GL:.��iP~�#37�Z{���`�g� ��k@E�[;}����i��bv ��̜��z���寽qƆ����]��h�݅�)�K1Ϟ�I\�?x��Ì��t�سy����i�6�Ϲ�9���,`V�\��O-ob�4�Y��T���@����^�DX�
+#�LR!�e���>�>"K�ZAFyr��Lbf_��h2}��(]�r�d�V�Rw�kj'�(�����@슦��@݂lQ���I6���:~��|F_���ָ^#������Â�l���/?���~xa~�e[26�a�̙��e���ݻ���xAcw���W��S�N�xp���'UX��f��w^������{0�����gh^�^y-���z�LG��S�Hp+͸Z��{ԮD\�B��d���8��`ؗ��P��NW���s �Q�����|{d��Y�?'lق�\2�`�T�7�lHW|��<�yh/�i-_]�s��f�B5������yA)�ġ��(���DB�)lz��8�IhӾ"�����(;�q�eq^C��'����p��z|�:�꺂]S�}G�M]M���w�W]!�?�_��`L'k*{����r���R��b��)Rrj~c{�3r�#��bۺ�-6a�LM���I�n]���
����4��RT?��$��	���2��v`�L����pkkowG�S<�dÁ'Q��4�Ve'����}�f�@{�1��oN$��3��q4��$$�̥��+�u8�����v�A�^���߻���I����m����E��V�rѳO,J7
/�F�x��l�77�������L06�k~g�h�D�	�#��
���9��|3��y������ag����2�Ϻ�i>Pq�)�
���Z�6쏝v��4_᠟�!y\p�������f��m�dgh��vԏ����|��V`�l�3���	���=�i�Qg2�rg�=c��2��׿7N�$ۗ�,m�7�F��NDB�^6[���=&�hE��$�N'��#��X��zAcf6���(j�TT��(�P?Y��xY�S[���E�L32�A��쬙����;A謮Μ<�03;t�w1�䍍��0p��&n�\6��D���4Q`>�1�A��B�?6E
�/Rm��'��\�ʤ2qO
��f'�D޸�F�h��q��Տ�� ��4t(��z�;��7;�l7�v܅oiQ<z8LA{��Ѽ�hN �̰���f��%P�d3'��3���������H���l��0e����
�S\:#UU��{�.�]!�_y�k����~��	���[oAٺp�Se!z�1i6��z�)���s�VWWo޼9??&�?��?�>�;�����UT���p0�b���o};R�n�gk}�qjYy����$p�Q�9?Ev�z}�=���N(e�ү��z_�3]�d9�4ew2�2�qs�1�3 �*�i����ʹ�G��t+ �m4d)Y�E�ԇ��tS���[[[��ۢ텧X
�����Y��P��W����>>����j�Yù�UG;;5{Cݝ�띩|���RX�(f�'\��f#ZB]�pji�u�hj�ݢ����U�7?vD�ۋ#	�)�A]��ں���1�s��:婷���4"x�-H���6;��9f.xU7��ݸ��R{�9�L\gU��NU#7n�:���@R���	��Ǵ�$p~�+-�z����ֳtg��a��P�Ai;ͷ�MWl,��v	��n�5�v�c�%><0&����z��4|���=x�� �&C�x�j&��A��[��p0�S���1�n��{�V$Ň#��f�-U�J���k�8	C���6{�U�&�95e��iU��Xt�8���iD�sa�xL,XH'���8U7��＃Uʋ|r�c�l׻�~W��@�<��6�R#p�̲���ө�8�1�S�}��@[�Yʜ*�5�MK޲����:>?M�
�Yp%�|W�yí.�*��̼������jl�O��E�7�Q��k�d(�]�b4�_2>���З����K�BU�a�ëfcR��R��fi�ԓ��2��yi�`���X�HUv�P�Z^��Ne��=c�e�-<�I��ȳs��3�v�f
��N(8x���D�w���I���ׯc�gϞ�^}�U��^d�F���"4�=�ٍ��t}��U�7>&�Bt��<����O�����׿n	�~};R���5}�8��1d$	ӣgiyyeaa��Q��,�I�#�VM~h7���͝f�#љL�� +��� ���@�xӉxD�󙌊8���J��y�C���a�h"��ҽ�����X�q�}��DkS�
��0*݄���H����<�'�*�h���C�Ô�����P'鬯��S��cW�L��Z]�x-	���������tTLW�gϩV����F�U��4.��/x�<A!x۠���h�9,Պ
����K�Nju)��|��mRr�l,gIU[�+Ql�q{��n��jzt�Q~b�+������0Y��m��3Ӫ>Y�,���-����b6�l����U�]��6���f�P����N��f\j�a&��д;��l�81%���'D�+�m�� ��c�LZ_�0RiC_tg��8%��莰���|ؙi4"����^�ߛ�ϙ�=s�=O<r�̙�f�V��ߡ�W�>$j��iLϏ��㰐 D�jK����s�v�D+Ew1ͦ��ǡ�<������Wf$��툛4Ȅ������5��5ú�t"�e_{�!�C/SK����cOv���.�ZG�Nw��K&G�j�e�>�t�����'�'�q2��D������:�8�[t�hӊ�VwA����pr�3%m�&z��'�ѦPZ&�NF�^^����`	��!8m3Q�XV ���P�"vL��&�37ם]�y�������S�W��]<=l�]o�َ=�z�6%1�3�	��P�hP�/�V��C��	"� �w�ɮ�����'��d���p �J�'�(x?%V��ڤU�����lϸ-�}�qc������т����ki�-����,ݨ%���<��~��"o�pc0s�^l�T]<nn2C�
M`2�0e��"aHC�<3�R�p�٩v�5JU0-ו��� [Z[!�i�Pf����s؃n�޽{�̇qO�>{Z�=�е�!��1�&����rV�5�Uґ�ՙ	�ȹ���ߏ��O�9�ӵ׷���8��I}������2��Q$�F�&��[o�uo�m�Bb_�Q��d���GϴhR��@�s�γ��{���kgᚭ}o4�[u��Y�L�&/Uf+��Dĵ���s{p -~l��GMỲy_���H��c�zA�c����*| �Es����up�(oQ3��E�oS�Rfϕ�՟���v��k�m�M8�#�I�-���į��
��e/�!��O;5s��P���U`�*���-
�s����%�w�v�=b�W�=L9BrS*����4ƓV��&���u}�j{y�Y���L
1&Y`jPZ��1)�*H<;�b����F��8��DX��R!�7K e��v��8��ГPbb�ɤۗGG���%����|��O>����Y&�47WDw�	�u�_u�㶑����F]�Pr�a[�&�#وܗ�rW�Z�$��h�;)�5����|�X��{���FWP�F��ڎ���$H�?�4��i^����_yv4|;���4��[��t�рt"�d]0����zP����N�n�ܹ���0��D7��D����%>WH=M��E����=G����(�����6B))b��d�8��>�]�.^T�Cׯ�4�`t&��T�q�C��>���Νsܛ�S*pB+7�䏨�1�k3C�6�4�H9������|�&����X='�r0u9h������
�����x�-E:��Ha��.�ܻ��{�w_8#����'#�Չ"�暺���=��T�Ѿ--��zGd%5��
�_�ڋKtH*�o���nm���N+��?�������<��#���'�`��)�b7jZwd���c��7� �Ц���9 ��"3oԷ�?O'(��J4i�t(pI�)��2zz�{���ޒ�^��_���<��T���KP��4��5a>h4Ϝ{��7O�$c�%��drx�߭��\e�U�7<؏Fø�H#Xk������p�4�y�������o)X;�0��˨���߫{�x������$�-^��
.U�蚋��뎱-�v��%?]��իw7��8{���J�s��-80V��KDq=�2�|�ȣ������z)S;f�/۬�0��Tr����˦�HSK(Vpm�s<������}w�o�n�n>N!�-]*��L��a[{�.�Ӫᐩ�w��Q��O��s7=�i75%sLE���#�3ꎮ�-�:Ǹ�8�����`��%��NF�VN�̷ڬ�j��%woS��F�����5�[�$�sQ����>u��$�S�_\�ፀ�aPAb/p`�&om���g~ؕ��t�f���;Acpj������`ߟX^°��$�M��7��������ٳ��N!_Q�h�s��W#A�	�L�n�+%�Ƌ`����j ����C�yxb9<�r�������@�F~���]�I��\�S��\�&FW�xAA������%�f0(�i&�#�E�4U�$[����7�0s��x0�cS�d�~���쌰�n�ED�:��X���+g����n!��"W �Z�,��N��bJ��g��y-%,�C:0ˬP�Uvwu2�h�!S�oml�,�2��ݻ+xc���<s3N%�	bZ%�fF���|T\�N*�Ò�C�6*#چ���<A�*�[�fd9��^��_���$lN����z���Kec��r�����NM~���@X�Kđ���@�[��v�
��x0���n��q���ړ(�����Q&�^B�>͂�h3�z���?#��!M@��)gk��藅������˗���6w����R�u��7A�P��Z��c�=��k��cx��u��ɓ'q��ݻ'�g����1E����M���[֝�&�����~����W��x�t��_6_~?�|raS����/Ai�i&�g����vǽ��O��f��R�)b��lbJ#��
��S�D�â�`��R�R�b�a�*�?
Q�������~�G;�a�w��:�vn�)�~��� w��J{F�7h�N�b�G\Ɋee; ɧ�w�͜?ީ9Ƌ�����<o�L�fv���q̑�P�*SwR1�"�"W��H�!%Y#í��ձ�-�3L]x�o�:���L=�ɺ�75g{^�R�U&<G[v	:v�W���s8�>l�ӃE`ַx���ݑ�[[?�������%]f+y��MG��Df�T��V���2�[M��`ܵx$.�J�B]�)2v���͵[]#P�}w�t��3�<s��y��#xH\!��wo]ҏ�逮�B�tj�8���F���wBZ]o��f�E�2%�m;`bb�n\�тL,	ޡzZ��oѡ1c��F�U�[1%ʛ�!�t�mwEzD��'|{�GDS��J߆���N�/gyn4J�"Ss����0��MQ��]Y�-����j҅�0p5No���n�$�UքR��(�_�}g=g�Ѵ����3��k%�(suͼj�)��d>d\aq���p��ށZ�CIj^�[�&��{�S����L��u�����TOJ�����jC3'@S�O�3e��.�(�����΃�C�̎��N���rC�3�4d���jo	���0�@��Fp��!��/���+���I��F4c�OQ%-9ڣ����^]#/kCJ~��VZ����YV�`�8K�+x���~=��ŷx��z뭯}�k�>��d�߼	��L��1w�↋�KX�_|��ŋ�6����d[Pc�n��[��C�}V����8���+W���>�z��l�:s��:��2'�W�:�sL�L"��o��ĉS�����|i�fziwv>�v_Y�e
�i�:"wr�uff�!��Q�ʝ$�h�S�1	�E�=��hf^�@?/f�s �V�]h�.�1�	Ξ��%[h�e����L�~���6���.�{饗���2��j��h>(uee	+0�fqq��]�}kk������~lll�MV���?�-��8�ń	\�3u|b�UW	JQ\��ъt�6W�Xu��U��P��.���7�$���@G����m2`�� ��Xo6�L��ֿ���2Ǹ�"(?m�������\�wf�f�x�N$n�f�P0DEVJ��_�C��^V�6���rk�Mf��h�15]3���{nD%�sę�#pA�ȏ>�0n>NؿQl��!�)gY������|m@N�x�D�����M|��9��.� �\��Hsם�[�ER����^�H����'������T��h��Ԙ���hމ�ꅾ3ӎ �%v��|wvo�k��<����l;���z�[��.��e&��������Ͻ�/���k^�Y�\
�W��8���nw~gwki����6&2�w�l3����9O���n]/���9Ϥ�^�n���;���k��;b��m�*�gJ�D�r/T|\B�iv�4\C�<��_f�X�3�7�5&���O���O.-
���W���8k���n��'T�hy�؉'/���Oz�����|i~ɦ��̄
�h�9݇���Ӳ�H�4[����̹Y!x�a/��w�����z�)hV���ck8��r��4ssҘ��B�2�3�p|vEbO�D������Si�A�h�E����BY��B��gF�l�I��^o��'����.t�CС����|�{3y|r5�i����kf�u�OƁ�:<..TK��a#l����v��W�����k����l�쭭��q�e�h{o��DY0T�������)���۸�����\-/_��sMc$�\�~�qf�F��o]�g>6�?�A�b|���� g��ɞ�a�������B�KKK��'O�L�'?� ��ض���P" et2�o��Gnc_ߒ�oC���hi;�������/��-~�Z��3g�:"�A%�2��`yP^��0{C�q��MQi+[�������j��Vz�A:U�v݈�Wp�w�y��V�<�L?�^\Z��XAG!���Nō7�]�:��c3���x1����2+z�*5����)����嵾�^T}�)�KYH�B��[F#D8�	:;^`�����	:&�
~}�GTfg�'��g7�6@�ڎ��lہ�&�Kl�� �V��W]nU�w�'x�6�_d� u��\�(%����2uJ���vF�*m�W�rR`V�Y������B�p��$_H2p�Am��!�m���F#|��fT�_�z+����ӧ����[/�����]bD�%-ۋ�Y��cR���A�d���$n4d�5�WZ�a��Xb�f���23�vNr�$@U��� �T�^���lI����]p���5P��nL|jw�0�����_����bs鄧|��&,����S��?����'�1h�n��u,�ٳk&M̟v��4f��n-�XL?f�Ւ|#��7y\fJw&���M>_����e���z*��:����6���M;��j��U�3�U4U�"�7dU�R�s��N��\�׭��[���R�Ǽ?�ږ�c�8}�B��E�4;'e3qe��b�O¨�#�ˑ�P�9��N�ʏtaUH�֦-��՚�1Ʒ������S�����o>��ȑ����)����Xn����paF��W$d�L[��8�����	��:C�B}��Q!�q*i�@��Z��>���8bF���_�'���g���Aw5� ً�:�{Ӵh��(����A*=�ЅV�Ye�E�ϒb�f��:A��}v��*|1c�U��j4�j��ޗM��K'��A�0��VL�����<���������Ϡ�&��ٖ,������x�$���L�P�n�ms��l|�ʫ��*i/ӱ5��W�$��
�Ɯ�@C[ۛ��]Wǧ�&���J����r�[A+���~�`З�s��>�g�ФtlK�z~�&5�ڊ��}��
�\_	�Q-�C5��(��j��|�[�1<�>w���Œy�N{��FŘZ��%���l�gKg����y��Bo=�GD�|�s�̎�#�u��kB-�2�CM=��"y[����Z��Ȣ�>�.��*��`S��1���;Z[o$+�G�{����{���OW�|
�=Ν?�?Ay����pv�S�>�=�/�;הO�.�$�Ӭ�
ţ�&��7��}���v�p��2J�i�dI��\���ڣO��;��G�6Y�%�<��lߨ�	9�òs��`�}���{��$�377�7O�`,-�h�,����q�����^����yV�>��R��w�;^.iA��G'��r���6��g�s��O&s�_*@�"&3v��]��S�P�{)anm<�J�L�U:U���w�[�����ݔ3��������f5�5�b��T.�4�M��^/��\s�MYȢD2d �������q�������Q�DtȦ��q�u3�1VմS.�=�s�VsS�KP��R�gN�D5�X�1h|)��=1�Dʗqj�$�J$�N;�֣`d��nk��P�K�����3�T��}|>4�A�u����O��z�|����6'l�MGjSz�$oX�g�(L��,�E�������������7������&�j�h1���Q�>���ّq���W������`�сt!P,�$N!����zRc�ϑ����"�i$����F�G#�m R�x饗(O_�u�U�0`6�-����������ˋ���$�(06~2J������y�/?�����oU�[��!L4{�_���5��`D�<�ȥ��.]:�D���G|����_�6����Y<�6M�IgL�:}�[K{.�wJ���*��ܜ�mt��*�|u�U+'�j���6�ͷ��8?�яE�fj�P�D�g��Ե�(@_���[Vu��P����S߃1e�4;���=V��Q.�c�z6�:H{�ަ8u�:�XS���gϞ�{�.Ys,d��A.���ʃ��`}[�:U�iֺ�^J�#d �J�bkk�*�%���%>��=����E�)��%DD�,��DZ��0�y�p�W�u�_T��:��j��Cō(*�+<��җ���)�hzs�kq��0����g���/�u��Or�� �%Vb�;{��z�K���y�IR�=�+�%����&aH�����I��%���5PH����e��]��D".^�R��}G�š������2��ع��d�7�פS*�-`��Fe6Z�rJO�'� �%^��<�e�a���q�(�k�#z�)(��H�����o�0��`�W�0�n�j�+��Q��̫81#�Eс�#���S�%_v)-�ְ�x��j�bZ�ˌ%�d)�vP��<�v1����*��~�1<R�ֺ����p�jY,׫K��$3y:�q�q��0�!(�8���H��*�٩�"�76! �A��{��>���W~���g�.Xfk�b��:��/m3U����9�"V�f���9��^__�<���-��Ot����e�&���_�Xĥ�/�������R���F���M{	�N����s�*^���t�Uw �{};R�"�qM�J�G��>�������=H^~�խ��3g�<��w\�|���A��w�#�&���_������og���D�]K�/w���ǚ�!��Q$|��G����y�����4F<PM�ԧH�}�6��o����c?�cO��FS�D
�&�{��Z�����������_�|��{�sB�zh,�U�>��4�P4�=��8��*�[�׺�2wGQ#�Y2��A���ͭ��������2�S��XO�00��/����i�	�f!���UV��պ����f���yM-.�k�I�J`�ɹu��ݿu�'[ט�[av���x�ğN�>5��v�`$5孎��cj��tx���[�������X�5��p)@��X� ��x����}��+�����x�A�m�l�+��x������\����hj\]E�|.$޺�g��rV=�	|o�q�\|�(�F�q℣$��Ao�G�"s����>�q��Б�F�Ӏ���XS�}��e$��:�<?����w:̜Ea�&�Lbl5N�Lg[���'і9��U�s��\�Ʈ��\�r=�G*��:q��/��*��S��?��<;���8�}ͯ4�,����(�r����2R��ؗ˸��Z*.\E����ø2����+[=�h�>�v�BW��7�0U�
�o�7�2/UTi" "�7���zbu�w�
�B۽iϰ\����W8�J��,(���|�$�QnF�,�m�sC�ä?��ߑ��*���g�]�N'�(K�dV��D\>��*�P�R�'�����p�R�ԽB��FX�hM�����W�C�_�L�����i4�q.KJ���'�@�
PYd�׎�X��a�`��ALɍ�h�����w;a�pb5��bp�t{c��?t���ϋݕ5p^��z~0:��\e�8�(��>�P�R)�6O��B�L��_|*���*�'!��XV6���?�1���~�2%�`^�7`FB]�Q���
Vq�G(b�9���}2�������Ӌ��${�B}��[w���C;�Αo}KR��x��u�Zb�"��Uh�[ST�o���s��������Ї�}�v�m�}xj���;��߹��Ļ�u���O}�S�?Y��#��^�~��2�O^C�j���y�k8�P,9�<pS��'��8&{��M(_O<���>�����_�ס���.��jM@�_�����'�������:�O��j]�j����J}+c��C5��T�2���5_K��V�F���M�LC!Ë����'~�H�`��N���7,��������w����F 6�����ҵ�^:�2��aۓ�Wɉv�3ɤF�������w~�w�j�NT���j�q�J�B�X4�m��[cE>�ܿ-U}.vv�5���_陦9��d�l��t�P%Ǿ@@�S���E���lo����?�y͸�}�9�zz;4'�����Qa���QT�CN��]׳n�acVW�^���g���=-iP�����aEbW��	�)�,��İ$��hTVp ��]�(�N�65�TZ{�4��5��Y°��q����K�����WM=�b����>���힣t(jQF�8�!��tj�W��'��-4�O5Z�X�;�/�G���A�2���cJ}���gJ���p���о���u˾<��ש�j�S��v��\I_7��e2jN��T*�O�Z��Ú���~�c��7Q�U�ʇ��Lv3�ؤ��^��Y�~�ĕ<�dS�N�)2;}�Y��he�>w���f85�w�+��6T�;w�,D�8����|G#aw`/��{�����	1⠥4u�WR�W�_����>[Mj<���˫4�"Rw��<ݹӏ���?��~�k���g�~��i��Ґ�k���;����8`�L5`�9>�>aG��-%�Ps����\���K�/?(�3^x�Йo�D�L02jƪ������:�pݾ/	��7$u������'WVg|%�L�Ω{{3�no� ?)b�VO�s����ٿ����g?����5����'��C����V1��X���զ���'���a�!,�\��?�?�?8;'��lKϰ��c*���׸�ɓ'������|�w~�w��v/]|�;;{����.9�`?~�����<�����pΈ���EZ�O(�ᜲ`<D�SO=����������ԩe�	l����/ ��>@0���K/��O~����&��I۷}���ۋN�jdh)&�ĸ�N�K�&��w�H��=��3?�3?�j#^v��z�R����{����ܹsTSp���䛚�7Ŕ
�:��ZOXsX���ő?�,�)�)�������|�#FB��l+���B�i|����=�&���:�-��R�S������������.;�B�kJo�����OqN��Kn��P�As�Fqq���Ï\�J�_k�c<�w ��v�+E�	C�'(�+&u�g���WwEa4t��/}�rl�4 �f�4�����ٲ�ްH�V���qC_�D������aw�bm �f�H@^�+�q�?XYY��bcc�������0���:dh��'�;��K� �~y�P_���n���#c.$>횲O,Q�V^Tƪ�'T�1�_C����EǕ��=iE�����4I:�?'��KG2��&{)��$W�\�J[{���%z�?=��z�_M�MS���򿼠͒[pY0�\�\�r*�����1M� ����ȣ�n���.�z.X <eb��vl�D�{V[r�2�{����dUi�̋)ez��D��Ȫ�`�;�ƘK�F�����:Bx�Q5����������	7��>�N�4E�c��}���g[�"Bt�ģfk�Z`M�*�[�����W�!�W�v[��\O�׸G0��q�� �G��Cψ ``��]�����5�� ���d(tp����9ho��&X�4s��J(�·�U�9vQg
\O��u��7�x��=�I�t��R�TH;"�Ee�b��Vhm}�R�'i(d��?pn�ˤO�W��+VhF�8�و��{����p�e�f��������������� �����Tf]Y��� ъ�.��K��ZIؠ'������.-�ٱ�gY`�s.�\��9�?��7��3( �
��o��o���+�K���1�@}�^-K6?U�.�6氮]�Q�@�X��������������YIH&�n�Z=!��u��w����'ww�nܸ���������ӟ�4H�ҥ��������#�n_�:"���1�Y���U��cS��f�nHa�����ӟ�	~�hՂ�*L�O�+���?�������/|��~��O�<I�fA�jS��S�G�̎����y ������+��T���xㆴ��Ї>��O~�̙3���:�4��\fr@������7�|��_�*eks�TI�nU"χ���"�f��ay�]��(�5���1��E�]mA�((ҺF2�b����ȏ|�{��A�蘼)��$�sV�+�����8N����x
(��#jo&Ԭ���n�ۗl��:$/�i#��?e��Vy�_IW�ڶe�{Ǝ�8{'HH� 	x���F�-a�QVY
�e(#���A�މ�%ے����w�c3�_�WM�,_���3~�<gh ������U�0k����4'7hj0�&B.L���	ᝎ��p�ϤE�in�!�(!	�_}�ck~��)�n��ϑ{�_��9Q�5]1^
"��U��[{pI|�$CB�$M)N�4��i��dO�~>_�~	�i����v�XHK<.׊_���D��&:oҲ�'��$�������Խ!��Ѓ��������a0,��x�^��PF^)�Ϡ�>�Z?��_��(�(�I&$�� $���Md/%9i��]b�l�g�N�hp^��i�¼bTו�U��G�\y����g��cfFc���#�"1��TYC�S~��_!Z�Z�%k�ԩ���d��S\�q�7�]�,ǎ��oSSn3d�bR��. ��[�e���o��#�;�{��^0��P��<��k���+�Z?9��`4\2���F�]]��6�^���hi4A�IIY �~��Hj�1��=n��e�|�i
���?8+I�������ѯ7�s�mm��v��N�Bn�իW۲��Z�F�A���E���y�F�Q��(�cN�0�Z�����*r�hqh96�ܰ}�|���7߼���V5��`(H'�*9MۙV���x,�D��,�a,�i���Ǐ�0��{��k֬�Zmin2R�%�z#��,/�$�%O��� 5��x���+����$V*maQ`->|��ϟ�b˶���d���e��=�8�����׊�;�ع�s�Ŀ����g�}���ٲL�<�^SU1�
P�Y���yÉ�W�(ib�p4�%��u���}�հg�������û��k��Fd���.��"�0��G���wl�v�Ե?���/�����
��WUV�L�=�f���pZr��2>�x��~���
��ǚ�,��"�.C������_t��e˖�7F��"T��T444����㡡��ئ��3@��z���}�ȑ`�33kȞ���:A�xD�' :���$QYY��т����ʆA:�D������d�>�$�������T.�4dh�j��
�w�pÉ'L:�s����A�AQ����Z�}�Μ�������[���5n�8�A��D�:
�Z��i��3z8e����^�C"��t���2�y����l������;0e��$CfXT��Q��!9��)&���T��d4.P��(�S�Lk����6eeB!�%���=�����$�zH3�B�X@�Eur��W�ԓt!�yN������+ۖ+�����y�ABRɔS=��-���d�Ȫ�?�Vt�I��n�7�p��Ojm,�x�`x�AO�5ӂ;�t�u9�Lڂ�No �<.�'�����_�^ғ��ǤD@3P������w�T����&��$����&���9Cw�iN*�n�hi����G_�{,���_�	X������#Gkk����������� ��<+u���Y��T�,	�AoES~�%���YMF�&˦���QA�D<Qk�jjf�V+��Bz�a�K�LژX���{Lɘ�7��+�v�L�o,����
�\��!%��$���A���&5�"�J}v�Qc����y��!�%�u\"��bɒSV>����Tn�&���B�sǝ�FJ���h\ÁSq��juLVK���
)��*���{{:����0��}~�����M�8�:_�{b�lcc#��[�@��5
mmm��������C�q��A���t�S`� ���e��	n���1v�X�m\&�aR�"T���Ca�ݪ7��NW��k�:�a�ޠ�������O��~�
��!]���A���x��b`��i �q�s�-�a=��s�~���m����Rqq�����u�^�Ν{����ƛ q,�5�b;�A$��T,�)��b�C¬�>�Q���jB5`�����.��2LL�0�1:�Y�6�1	�=~R�� R]�.L�j�e��պ\}8������}��w����pC��uq�U��ن���,�� �7	�#C��\+��_ �={��F���������[L���(���`��D���0;?�0֭� :��%g�y�#�<�u�V��!�QhI�K�.�&�W����(BL�����0��~�	�`F�	����3*i�؅g�ѭ�h21P=pĈ�ƯK�޼hѢ�o���/�����t0��s��D mZ맽�i�(���	*ₗʝ�@'����s�i������[����P;�N�ƃ7k׮�>}��U�^�����
� �3C{v�c����^7��\y�U����q:SEEE9%�Ըg$�
#�k֬��2�w�Λ�h�9Q�Qc �H��DD��^V���������kEYY K�\��6��!J�K���M��ѴIC���`PG{�)uJ-Q3rM��,�_LzHaXQ%W���)������~�ǰ<x�`ff.��A1���=1PA���'@�Q��
��Pg���d.�?��`����˦Q)x���q=w�3m�q8H���zZq���%b���^s(�d�	?�:��0̰��]�A�8��CD�&��nZUML3�fzH�����+ �DA'��&FX%*t��������裏>���LKv<�O\�qa��Pޗ��C~��2S��Z���}wt�O��sϝf��СC'�PG('��[rg<D��(��):�HP""��
�[�0E��.5X+���~E¿SĬW�K��0��LP����T��`TǏ6fLJ�b)Z%��
�!Qi6K:+����ۭ�P6oj��(�2
����D��6W���բ��_�3A��d!��/���*�l��)	���b+�Jz�0���wHp=�||�|��ɠg, �~�c���Ɓ�]��˃
�.TWW7�4WTT@<�[;x�]�`Np�X������~j J��)Z��_��?܋}�f��������i\��ic��`QR�����X��OBw��O�K�R(�)[�<�����_|Ɩ�9:;Y�m߹��/��%�����z�*�J�Ur��K8��9Y�1IL����裏B=�V�`���j���X]�o��-h˒��ƽ���/ X�w���I'���O��$�h;�iy��"j��'����@g)��͖�[�n1�q��/�7o�����se~!������JJ}}^�\-[-T^p �z���L�����䓧}ǁ�" #�w����Ù�X�Q-Up��8<�O��=�s���X���~s�����~�Ѡe����ʊ��9�(�.�ꏁg�e��詙�9�I�~�Ϛ��?H�������={�h��=�W��'Lr�;���O�S��V�x��/|��'���b Y���/�\�v�v�s0�Y�Y�a������)�d����x`9����.j�w��6�WH���0>��c���n���+��~�)p@<FUQ32(�R��5`���F)��I�a�������/�A����JN^�/�d�%'���F:�6>ڈu�����u�D��vZ���\�$���I������������zɭW߸��%7�����%�X�fUZ��6�+�W��W{�Q���ħ䵥�y�s*:Y���(�,W4���3����pؚ[-�15��z��\���`N�r~�x�2 �A�'��H��hs`Ty�T�W�T�W��}xʔ)�ܜ���O�S���nGJ����E�7n�� L���d`I�֧�J& �mB��勷�Z�U89�"�u�)PԠ��MG��6�j�-��$S��c`�dB
��bZ �ʶ�woo?�l��9N9�I�w:|j�,K����@�J왍��l�JÍ5
i�����@��j}�JOEZ�Q�V+N4(�M�����>���N�W��\\p��Y��)@l�0�` y�F°y����{��K��|G�Ϙ]�w���?�O��S�[s�\�͡�l4���k���Z��i�E`6pR��c*�"ke4��W�_�W�I$E��$WD����l�0�dd�Q uw,��T��<G_Sy�g0���m��Bg��m:]FLr�UZU������ �:�FV��T�gZC�	Y��uj��-VY��US(@�P�P�� ,:��`Io��T,���1��<�"Ip�zh�a�$���՜_\dɴ�u4+z�Z���㉰V��uv��{|�s���d�$$h�	&�'� ��Uh��2�b�0~:&����o��Oj�nͦ?g$괿����~�N��G���տK����!� �[.�:s��^��Bmi	��t��O��8�I`D:կS�w��e�j0I,Ї~�{�>���O?=n�8X���)\d �O��q��)����y��~��V_Z�"�0����fZ��M��AmHR	�#G� ��h�c��C*+o���믿���E����쩸i(Ӛ�P��
7ihhx���1�ɓ'�����=���I�Ρ졍V��꥗����܌r�A�l��`Q`L�����W�롓�oX?�b�{�7�\���p�F˩�,U�fC�������t?�2vO>����p�,��5j�֭���R�R�c���qm������/D�Υ�)P�a#��'+?���z��,X����ͫzoK�� kH%<_d�=vp|eذa�
���3g��+��v���=��hC���>��Vj[�?1�	�f1��6ך�;c���Z�|9�v^�]��Ž�'&��c)��h��l�2ǝ�H�V���yL���3�lذa�ҥn�X��vaC����^D�b��� �3���\��UxVJ�)�X�(����(|��/������1d���;ځ�Ca:�-�(a�-|�G�-�ͦ�k1�Ǟ����<p�޽{O�T#*���n�ta/�����W��Ka#E�0�I��H [6ps)�ݑa���"��#c��	A��"�Ad��h8PIy�a��1���G�]@�� 	"0��X}+i�$U>\�DR�L�������)"JKR$��^���&Ej��W�Q��l�����8VR:���+V㤥��l+�W�Ch�>|����{��M�'�}aŊ���Ӳe�c��2."ƙ��ɣ���AxM�L�^i������p
{MP�
�,
FŹ'��JV�� x׬�<bD���T7f����']]]�l"CL�(������>�3�Ν���2y�DP~�߇�����=aeR�����vJ33�`Xo��^��0
i2�G���Pr ����q�P�"� �� ���mv�/���2Us�� ΒB��͛�N��/(���4�͡`�j����ukZ�Z��iӰ>m��'��6L�z���p��Iq��9N��1j!sԢ|{��v؄W\{���������ȑ#�o�#��
�.����F�������{�Dľ}��t`	��o���ꫯ��:p� ��v�߅e����$��X3�p��om}������b�^`a��`�_l�r��ȫi $c���A�6:p����I:�Q���_�A��_Q%�X�x�o��_<�WfeA�9�շ�|�f��@��ͽ`̘1��ߠ�`����@F`�h0��H<q��_䱿.]z���_�ſ�]7|x�+�>[I�zZ �nXMV�������o{��/.))J���֘�&:{�Fa,@�K�o�m AjC&����/��2�d�ʕs�́��%�u8g̹��vuu��ƍn���/_p�M7����bId����UIQOɾhԅ�C�����I@��xa�����]�47���� V�l�b��]����/@F#F����Z,tF��8阦��;5l�P|���=��E�o�������?aOǍ�`��O3<�(�9�t��ݤ�������>d6��_~����j2):�� ��|�mB�Y��k��sJ�æ��x�:�*(��`7���j�[�hѪU������}>���G�F������/0��kD�O�H�@O�å���� ŦH��2�����^(l.k*d��ĥ��"&�7��
عs'�e�ԩ[�n}��|�A|��"t�˅D�^�ǋI�#�z�}��! O*�gP�&o(��ܾ�^���ʟ}���#F�ݰc��qiV���Ƽ���p�H���+*m�ٳe�4��6V��lljw��O>�������뱇��2�����$OFR*����=u%KR}J��TP��WG-�ea�I�6�������sk&U�+�d�Z])E�щF�ƢZ)J�}��#J$����D�K�3�uj����2���[R2	W9��M���e�giZ��{Ѩ��Y���E��!��^tӑ�ٓ�,�X �:���߫8��ޗ�c�v)^oWg'e'�3z]n�>�p�'L��SOM�6����{<��n����SCe�]]�d��CkO³���HMM�#��[��ܼ��W�Ҫ���\�H�L�F&7�5K�>��t�;���[���� r��|L��+z�̘R�0�;���W~�噳gC:��v�"O1)��N��VaY�&��3�� ���#���Ç9� {m�:o��zvU*2ND[0��L�z��TP��)�<]ЂE%�t��r�_o��/O�"�OLJT>��e�o�VI�"�?b4j;��p"��e[5Z��ٸ��ޓgL��}m���LK�`��L�Q��{:��pIR,fuR���j��$�թD9J\�^�����1�Re�d*
24*� �C&�R*�Jpt�Z��d�����t9-���8�\
�ٶo���!V��6���$�<~��j�:**.�Ģ��I�b��Vx��b�Ξ={۶m`�iӦ?~�&� |�q Op��{'DvCJs�>�B�L��WZ��M��C�����XR>4Mc�[����|�a��Ӊ�Ν�``> /��)S�P\*���{�3�8��T�.j�d6)�g*�tjo<�������d������::��f͚=|��D2�>��!�<B����U�x�=���?��U7�x�Nd���~s�=,4����a��0z�p!ߣ����aGu��ݻwc"x�}���o��`���c�A�_q�����c�\8��N��Â����Kz���v�O?�����ϙ�P����*�����ϻ�{ɒ%YY���@�$<���5�#srl�z�x cǎŮA�}��'��>'���cw�~��zxV Mt۷�b��6m�ӟ�FǏ2ͰR��tfyj +37A�(�wï��m���\VVF�q y&�V
ك�uH��F���`�X���7�袋���i*l��Yr+Ph���_�fP6+�Q��`(5(
�̧���-բ��eo'�zٲeP��->�c�	��`6$�+������z�S\�y�=���F�M7݈�c�?Y��С��:W��>x#*"��왋�F-��^%vN�lٲEVt�>��������0�|���wa%�X[�!M��WsK3����% ������իW��X.���K/���;����1�.�(Xm���{E8~�#�*�$NR�MX�I�dW�l�N���+Ir�E�q\�� ĉe���vʢ�x	��~�^9r�0K
ွZ*.)߻s�_|����b�KJ�9�\Am�d'�7�ĉO�<[B맗4��-�`O9�2!ڥ�Y�����f�v:i� ��> ����F���a.�KN�2C�a[�DG�y�i�~��㏷�5�j-{}� � f�$9z�K�)Ut|���dx�Lpn<u�U�܉;.J���H4����u7;|�������������ò��6�P�2����C�_u�U[~�P^^އ%��F4�m�ޞg�+S�Z����1h}ЌI����Ɠ�f�X8+.,/��3`᪝���)�(dH�Ȏ��H[�au�N�bj�H=�'L(.R��>�}i<��;W�*4�0Ó+����&I~AhkT��+)v����W���������a���^x��C'���V'	����ʛ<y*���۔d�t����Vc}p%�k˵u�+d.�A���>�/B>�ڵBc� $pp�1�'&&SI�q�ϚO*��:���ږ��x��h}��b9(��MQ�g�}6��q�&
�B��F)��+�+Dl�R�x�O'�*)~�С/>}�7j4��qt�+��<7'���ѭR�#�h�U_�o3��7mݼ��+��P O�� )W�.��m�w����u�>���,Z��9l�0������[K�,�>�D�´��	G����ӳ����������O>��Ƿ@�3f��6o޺iӖu�6@���0c�
�s��������7q�D�-�p��嶬\O����A]KbZ����_|������/b�z{�rr2�*l�՚�>
�?z���#��6�C���	��o���;w.t�U�@yXP!g�p�۷v�z�u��;wl��wo����bGcv uƞ�J�гT>V�����s�́u;r�p�.e4�p=(Oo b���5��+((�� A��߿��h,X�%��t�I&'�� ��a֧�z*��׿���G�� =A_jP|(�!y�\cv�z(�GQ��/ $�Ͱ�͕�I�p��2H��'M��o�2޸q�̙3�;�<���֙�.l:��%Ű������S����.��?(��nL��w��I�ΐ0�����R�/��Y6o�#�5�t; �D1��FY�k��	L�I�u�����g�N�*e�0�XyiaQa�h*���1��>wVQ1���;G�Y��?N�>4�yGWnnaJ
E�*#MP#�"gWqI%��Ј-�*�P�JCB�S\����Qړ��ʚQMj2�'Ť0W%�z��L��֎N�Y2��j�QG.��Ϡ7�N�.a��#7i����:��<B���S��v�w��Z�n��� ����̶�.
�H&$�	[\���q�N��k��J��p�7���-))�\~�B�J��=u��R��%�h��-//v��2xX̶�:}�h4XPX��V�����b��ag���������������!�d��MC�$E��u{z`z����>����*cfF�^��zz��)��j�޴�:�YOH���8SD�M����z�Ԗ^p�
R��iժU_�Zs�u׭��l_H�dU���1Z(�"ܐk�<�=X��CRWG<��+�uz�wA>���V~B/�1�nm1�a'82��B~�З��MƵ�נ1-`��,˱��3m�H<k�����j�NJx��-�̡X�I-TZg\֦b����
�%E�; �Հ����N��Z�!����JY{�27L�)�����uS[K�=��?~
���`�a���<G��v�x#�_��mvQ�#������]���'��� ��0qNN�|�¯v���7C������nXA��L�?|��_�E��m7+�J��*zA��W��V���ϵ���O@�XC���#�H���Y�s���#c�OG�I�sJ�<W~���o�y�=K�w�	D��c*��9W��Gy䤓N�2y��`����<JX�$��?��rHewO7�������O��b"6������cӳ�# ����U�^5��\:��co�h9x�� �g�ʕ���:�,���ˊt,�
̀�X�+����믿��K(��f��P�(�h�����=~�(�� T}}�H���K�׊!�����?�x饗}��G�+���߽{���f��s��Nƿ�k�u6q�uX�y�o6gb��\P���+�X ���SO=��Er�G>qg��a$@3X�^x�s��כ�F>�Sm�0C�����e�u���_�
ǎ���;F :X:8NE����0�u<�;vc��{�.]��<���cǎ�]��0_�Aj���q�M7�s�]i��^�>��r��u�ρ�Pи��.���?�y���cI1�$x��[xÛΕ�0�~��s�����%,�
؋3c�B��C����!#G�8�+�������1Z�X�$��b�H��`��z�ul�ҥ7_z��Ϭ����Eb�P4�N`���G�>�9�g͞=��i�H��f���/��'UF�&�2�ca��/�J#��V��}�/�!��Q�H�,VX6��^�#���)\,���b��{S���驢�oV�>s�i���ēO<���{��)*,�Nq�Q,J+��7��}2��V�,�8;��z����.�&MI�(����X`):�ˤ�N��5��^����0�qF�s������� ���[�,;Ǌ�ΰXӑ��@9������d4��S]t���o�}��qX��.��v�3\XvBIA��T7��B\�n����!w �'�X�ٳg555޿��O>�d4B��� ��mI��@� �����_66�ǳ�X���2��3��F'�̤pP{C>�7�-�5�=��"iX@�Z���MZ����1cƀ�ݡ0�5����!+�&��$�`L�fyA�L1��Ux����1�^͍�F�ҫx�֚��O�9�KSskkk}�����F�������npJ�Eֲ�f�8� ��{VTT�2�l5c�,v{�	B�m۶a�@EԜ�l	��h�e�v_��\���Q�!w���%��CyҌY�������a�%^ÇS��i����;�G@}2�E���en[g�t����ކV��n\���sϖUR$j)�J�Q����o()�%c��3w�zvn�<y�\{V]�}{v�ޱ�uhm�^��8ߞ�����/8��{�=��g�q��3�M�4P
w��S7}�6s�Q(!�.�	�:d
vs�Zj/V?��«��
{	F���oa_v�e<V6�=�x
�k����7n��DH�� �[�v-`�8�'�
Ü��D�a�_���pii1��M7-�N��9�<}��;v�-F�z #J&�D�� C[�l��R';0�z3�Z���tB���~����>�ڹs�aà���&ؔm߾����� Jվ�� D�U�CY�R1�T��^}�UhAL��1�/�q��g�y�/�4kz�8%���c��b��)|����^{���r��X;.�ǩ����A��04q�]�0I%�:�zɝ(��
�X��?�x�����ͱ (�g��;����|��9r2����kk���[�n.))����d�@�H`J.��:>%�tttA��K$�}n(n�/�6}�#�<�EN�(��--m��.W��f�|��}}T�{hEIVNΎ-���=����^u��};���&�����VO�C���_��!_v�q�$����͟v���_c���S� �Uz�֒�z}E�P�RF�\���TR�4[��&� ��ꉙL��]͠=���T�.���aф���y��'���߼u�b�A�C�ʇV����x�\�,[v��7b�X,���ݲs�՚���ۮ[�+�����╕C�J�%%M[��QPZ ���E�"J1��6�������쏗bS*+(ֺ�����b��x$���]*+;��ѡ�k�D�u"�<j�n+*���>�}R��z$Oܑ�6	Gbז?����/�
�m�έC�V���r�h	�P�f~~'�p�a"?�����}��m�F�����=g6�z�h3�[ZV�����(�UlkQiN��F`wn��N�+����Wb�XdaM֯�	o�{��%��
����O���)*-������|�/^PR����˪�mz�US����3Q��4z=��v����+ߐ��@:���6��M ����c��	Y�����D*��Gtr���ɞ��
z{��:g7��\=��0���c��O>aJfv���0��.�*Oj�A�Ah/���q���� lBa/��l��:ۓI�^�Mh��P�d�R�n+D���� ����}֬Ys�-Pt�>�������,Y^ZCޅhJJ�������Ύ��F6䊊�>_���fr���(
��9�C�bl���ǁ�T���,�xy��'x�N��L�܁Wt�I�*�օ�\x\�rߔ)S(9�CѸ����/����,L��g�h�C�`p�VV�U V����4FOH"� �%c�l��C������ڬ>���s)�ȷQQ+3N�J�ML�P-�ٱc��Rv_��_"�������VJ^��˽e�.k�t2 ���.��:�H���r�x�`�q����$,�2bq����t�*'��8̳lٲ_E��+�+/<����'�0q�ʕ���_y�����^�?n����6����	Bo�q;v���Lk�g�y����>��Ҟ�'�C�@j�$�!{�!�/���w��	���GS���w��/����+�2}�����06���7�G�Ʒ PZZ��)^s@��~@
���+#�
r�d�jj���*L+($HOf�,v\�!���x�5�\���C�f�{�;p��h㧟~�@Z�ݻ��w�ü���'N���r�9�#x��y�3��Ky���^���z�ؽ�Ŝ0aƶz�j�p�޽��e��m����@���
HU|�����'\���ɹ�X�ݻwc%qO 3�?��XR y&H� �hӶ���g��.���/�¡�r�	���`�`J@p�p*AYyyC�! �?x�j���u�l�����ϟ��\�iʹ�h�z|t4�����MDcDTG�`�ں:T��0!����㩨�2j��`�e�.���թ����m0Ć�W��e��:��d9z���h���e@f�L�x�r�0z(!6t�N7���J��=��'�����1½۰��M��^���az�L;q���=���B^oݺ����XFQo�(�&.ƾ`}��wo/�n��Oݞ<�d��~
��c,Z8��i4ZЌ��`����B������	;>g�9�<%FK[`�¡ЁRI�Q��sv�:�f�jjjF��cǖw�y��˯��o������;>v�3�į,���(�{��� �ܼ���~��+ɖp��a��D�9�QRV����n��	��rA[`0x:�6��u����g�ţ�Z�' (\��Ӯ�?���ς+ׯ[���G�D	E��)��E��@-*}�����WJ�`�Ǡ�c�p*A�T�"=���`3�Z;[{�I�"ԧ
R�Dn�-�98� ����GBa�n�j��*;�S�P56��*eeZ]�I`0���/���·��� � �±���R�������'�G��O�칐�m���J"]"�����]�L���e���^o$L�q o�FMX��rg �8i�3#��p�����8�[I��a;`,H��	���X��ͼ/`I싒��#@Z�=ԗ���O��H�T��)�?�@�g�WJUi��%���c͢X0�!�9��dP�W�о��J�FEKv��h�i��P8!��Tz�YߤI{����?���8}��t:�j~#)Z9����?��y�Np �3��P��o���F���V�x	|�?�i"�ذ��y��Χg?�8�MD����o�vw�ڵ�C�_~y�
d�/S*���%Q��_�x��{�c��@�6�57���ڲ_��>r(M:�㶳S�N5��o�|�C�,�����j�ڼ\��,cz+٭�f�ر��/ ����Ed�ffee��G(Sў�OD?��ӑ#G.Zt�̙3�����s�Ν{�=w�ڨ��(�'H���'z|�w�>���:����o!���� 2m�r�.��}�V����v\�p!�@�29���b�~N�v��.��K��W�X�ß����O>�e������V�0RfL�-��Xs�x�!t����7`W�@�P�<x��56�
&��7��-z!�1e�<�������l/��5z��͛7?��s0�}��(=dŎ�Q���/p���ݰp�E�x�)pg+:����k�l���T5�j5z\��|��;���?z{��ڠ3�i5��Y�,���������c�=6�dRu���q�Ksl��SQ0��:�tu4vvw�Q��3D
��9���D����:_P�3e��|^:���K�KJR���f���ʶ�z
�LD�d���cxMMk��^wp��
�5q�֘a26cr��?M��9&fc���~�W��nVYi��4C�K�:]Sƞr���d*Q;l(�l��ػ�'M?�租v�7��~t�	S"1oS�,���ݻ(�؞S �<z�U��tB��W+�M�f1���(�E/X4��b�)�		huҤ��
�T����x޼�g�8V^Y\Rh�R8�Y3���������߻s�/���jr�۠}\v	�]}��4����:ljn� �vvQl�U@g�h�t�������u�zp�[�<�@P@iI���Z��
�Ԫ�|����JmM-�k�_���:(����9s��!��#<�%;���V��lR���e�؆�Uoز��W_]z󲒊�`4R3���o���:�������vm0,w9b��P0Ch/ґ��9��$R&�Ū���9֯�G�93)����_r��w�dWUU���0��nP�������.+�DBe�뱂Ś����a�� (5��x#�C��U��=���JN��
�pR�U�h*M��q)�R�:��M$=��76�2a���e����,�y��v,��ŷ���=r�00E )O�?;�N��s�Ky�W5r(��#�{z�'ϜY�e�^�WO��y�l�A�c�1Z\ ��k��@,٤��6�-'{�a@�T-�� ���,P�"�K��xq�g:һ�H���[A�5u���Z����I"~�9�ə���e�?X��`�Ú�8�{�=ȑ�O�hX���-GS�I���0��qqH����H@�=���BT1zP�6Pq�5k�l߾�����<`j�%�8��|�J�Uz��B��K��h�T��d�d|��/��Ɵ�i3f��G("W q�<��=T�mb���0���-饗���ŋ���B Bv��PWδ��B�%�?�K��N (�3���8�}���z��߷� ~e��	�l�2��\��~�tꩧ������X���x(��<�W��0RmqҮ]�c! 靖�A�Ȓh�\�d2��Ʈ��A�n/++imm_��w�}T����\G��%xq0~N�=z4@4��p�e���ϱ&YMr_K�p�Tܼy+������{ꩧ0�����a鸴 n��!1(l�
z��K�.}�g d1ZI$p2p�3,6��;����+�����2����R�4lM�`��\�F���@���kѢ�@x�R�i�&0�e�_��c��d�l[6�d�P��(L�UYSd��3ϼ���J���U��blP�fs\���s��W��v<�ԙ����R�SlY��9)�E��%��U��6�ߋ1dfX�)�j@�7'�!��y���e������u���Ӈ*�nO�6n���b2�3&��K8�e��vH�Ḥh�Z��/�3h�99yd��m6l7�\�Ș1T���KѸE"jՁM��M[6��Οs>t��'�(B�0@1H[�/7���Z-v�}T���ڽ�z��j�lpc�^B������`��/��s�y`|PHB�B�ǶVUU�|�«�����6Ü��Xa��"q24CA
ZR�Z�0Y�?~�+�x ���Z��Ǐ�,T��A�A	�O/++��{o��:x���`ʘ�4�F#��Ye�%�E�I96�%0��}���qΚ5� `d��{�[q�,����r��v��-��7.���ON<�DC·0�o>����Ԣ�&���esfn<�5:��ҫu9����M8-�l5�숦�/#��['������3*�k�!'5�SQ��̜���^-G}��FP��0�ɷgfeg;���^2�(��)�C�8�MĦ�b�Im!�r�x��-���+�=��S�� 7n���b�I��b��VT�t�:|kƌ��܀�H}��]X�ݻ�.���*�o�%��baE=>���h1*�,�#c
��@��+�:��<
r-?�5�B�j<\���d��+�NN�n��D~n���������\to���]��)�qp�v~~!D�w�}��GA^/X� �y1)������8��J%�"� ���[��P�"D��*M���������]�Uv��z�t-M�~��.������Q�v>��|�ZY���L6����ڊ���Q�:;:�\�Vjhe�^O�����H0c'0+��IjܮT�bq��@�JwUT�A���z�o�]��$Q"�(�i�?\)�t�ή�^��@8B��XGSRB��\�
2t۶��sHz��9�T�(��u�ꎎN�I�A���A����������7�;�n����zUR�l1UY*=^�����I&�QcFBL�;�����n��|��C�_�N���1��c)|�+ �>|$����y�L�����ޥbX��0��h.������� ����;n���O��gϞ�e��qXN �0??�UV�rt�ٷw�SV��}zף�(׻�����?��==�T*a�S( v�;�;I�ݨ�<g�۽�E��@N�5��`�I�&�x�E��7��u�]�
�RVV�a"�G���JJ�(W�����矽��+��~���n���/��/�a�y�d�ɶe�����,sK�aLdܨj&�w����[��
�M��hШh����n���}��Լ��q�9erÑC�]s�E@Sj�
L:ɔ�Oă	#Y�fK&����:z\�UVk��ux"�A1�
��l# N���G����ڜ`��	B����;�`��&]2Zd�J���}=m۳rCF�WK9a�h2 �uF�,��/CH��7�����;~�X��
Css�Nm�)̋Iv774aF������������o?����ӟ����z�� � 7;������x���-[���	n�������e���lu�gyِb�V͚ի�z�����2#�8�c��I��v�֟��}p�ygA����/I�xiIU�}�dMF�=���۹m�%�:u���V~ ��O>�����Fe
��
����;��sO�v�8�'�K���zɵð4>�G�y�O�<� � ����q���tw�����~��g�~��nl��E�pO !n+�mT1�.�s��a�0����vt4���:��W<s�m���/��Riq��]�j�b2-B�H:%7�{c�DFFf��\���n�p��VL�&���T�@��@�Wͳٲ%����l��,������1;te�f��n�$��F�^�������XRni��qp^M�IԼ����u��Nae��Y�]��M�1{}�K3M&s8bh�z�t�p�ٗΛ7O��xl�-�+#G���-�T���Bh��}��ISj�+*�a�����e�����'��|�x��3G.���s�/I�;�Gc�h�"�D���P)�v�:�ZQҊ�@޳M�G��	�Y�u�}�WA�3S^�?9rdf��A�&DjPǩ���ُ:��Y/�+��E,��2��ڵ���d���h��	��$�gʖ=n��ݰ��h�&쏋u0r~Q��!���ǌo�ٳ�A�o��_���_����������b�D�.����S%
q�����o��� آ"�<
98̖�m��S� ���=����o@GG;�7�oh�N8�Z�jT�7�p�-�p`Qb��Y�K 4$�5��t�x�q.����ӧ#�����孷���0%%q؏�r��/�Dƥ�������#]�p������:��w�y��_�x��m~��u�L������&vvR�\NN��D8Ι"ZE�1��~�-,XiP� �r�l:��;Va �sӝr8>���h�?���Ǘ_~�-�6��B@�< j� cL!��=-N"t��9�b�}^P)@:S������⋯ 5p�]M��.�|xƘ5�)ѭk����x�С��>��/(*�Ut
Ș-|�㩱�� MM���·`�I�߃�nO�)@�Za�->��\�s)R*���?��}̝��1<���S�"����+��`Y�f��$#�
���a��ˮ�����%�R�)00l�ha>���;���ʸ^d~.��R'��C����{�SP�~0I
�I%����h��؎�1�vt��u��hh�zEҩu�4�L�$�F�S�Ɋ�2��qݏ ���j�OI����:siXH��	��N0ZȻ��|뢋.��[�v��^��x�������p�F��cH!�D��rxĈ���}{�>���o��VJ��@��Az=e��6�	��lݺu��?�������O�-s5'<��_�4wtun�i���^z�Щ�ȏ��Ôܽ{7�3m�4@�3� 3�������b)�]�~`���,�0q��&%7n���Ͽ��GP��@<�!����U ?����{�?��1c�`7a��E��5�Z�j'�M	ݾ���g���� 
��UJ���b������xa���GCA���b��I�Dƹ�C�)�K�tw;�6j3cU���m��&�р�Y��j2�������YE|}�q�� �`=~��d������a �0tI��Ȝ��U*,�y�+1�[���e�):Ҿ�ǚ������}\Έ�����!��Q7B%��>�Úop��fF�� ���a�Ȣ��7�N�s�N���	.��B�V|�e��8x�����Ax�S�L`.<�\E5P��k֥_l�q`e��a����	���8�ݟr⌴Q�������x�*3�M����_ �m��?�1k��\r	�R�:�[��M�@�F#� �n��-�&�b�;�;]�H꣆��Zu�L�����������5������\�e��EZ���s�9�6[���|��TX��r�#! O�Сr�裏B���=z�FM�dTt�b�j����B:�x%�)��'���z���m�~�ذ��kK��0��O>��u�n���3�8�g\FU��p(���g��U�+�͛ 2Ə,�L%�|�;���1�S���(�%����z֬���Y��e}~�sո�>h��W�<c���.^�d�x:��;���Tr�pw��N�|ꅨ�{����*�x�رS�ꫯ@�P���r�랊%ͤϰ��
�`��և~�nOԫ##����{�m۶+	��U���R�6�ѳ���W���+��r
>��{��O<�9���`H������K{Mm�#R% ���A��Y����� 9nϱ[D�ń�M���#�����O?�8UYY��B�ē	蕔��rt'�q|+��|R<����W`?�w盯��N(���#F9���N�cY��~:Y��Z��ǱH2�(�I��X��l�=O?i
P�틯�X�'��R�Fo ���mJ* �Oat�P\T���q�:j�(NQ�W�d�����@ss��Rh�W��-;���,3�*����
���޺�UL���Pm�I��F�YRUI~���5݆$I�S��J4*r$��C̙J���q{{W�	;�Q�k$�ŤK%似BEK�:�nl����b�?xoeqqɹg�3s����s�Z_{�u�(맽��i��pts^b"��=n7�H��S%u�-]���~��goQ^i4��t�-�7�r������[�Qrʔ�_��;W~���߮޳��UW]���5f`mO_H&Ú�m��@/�+�C[����1��O?s�E�y�/��r��I�]wt�NQ�������q*�M,Π�6z����}���F����p�BX���!s?t����d��ܼy�ܹ�v���{lܸqgs}3fQ7��g;�[!� |ȳeT��6��|�i�]z��g�:s�s�B`V�m�lULeٹ��bIm�hmv����f(6KF��X����Q��TZRst�f�an����B%�"�N��"��R��>.�u�|�o��E񰳧��q���ޥ�M����f�δfa��6 3 h��j��ʌ�]�d���Pv�R��*�0��t>���s��&���������<s��7�\S7�s��z:��A*o�NE�7�(p���y�رee�X���v�*#C�j�i����0,�*�i՞|�H�+-�3���- 
�X7����T���A���垨�0x&O��FA�F��,&j2r9����|��t�n�
J
f͚�}7���������"/�!��S��P������A9m�+�s��\�g�,	+���?m-q����릣VC6�dr)"X`F����ӋY��7�ƁY	~�M	)�쎻G��b���X2�&ז��<��ï��
9U	L�wE�(7:���*��gq4�ْ�M�x.�o��N`Þv�R�l��ɂ���كU�3g���_?u���V(!�ɬ��<@����g���[����D X��E�U$�Q>�L{��1�\vR���>�a���&�/N�4�믿^�z5����7���b�TR���[��*@�_2c;����XX�*���`�k׮�:@O�'D{#�B"���n�U)��J�G�� W�`���;L�4	���o\�r%T5,�1�DM��L|Fʌl0f����s���he��2���d7n.�~1z`��]�8����P]n�{n�Q�s��?����O��ǿ@ �V)��Vb��a ����;'L��dP�B,NN&��z�w�5AOW��9����NXuՕ�r����-����UJ��%��.�2�es3��2e>�����~� Ͼ�j�����T�[�~���c�C^a�,��5�=	<�'F
��N�8���:���Jh9z*,��pYDj�(�N5(���H�T<��X'<�;
�b�RU)y��}���F�^�3}�t��CL�ও
lph4.��5X[���n��&g/a��oQ;���1����y�W�����?��ue%e�$�Pw�$��$5�z���<5Y�9՚xQQ����$�����/�X��Yf�ˑ��!�!�C��P0�{,�)S^{�5��&L l!j'`w8� �c�wA�0�0��#G���2��~�m+V�v��P0�k�
�t�hq��㦛I����d���2@'�>�l�hZ��p��I-.1���j��
x@�@�57Ph��B���'�εg�u�YS'Sݺ�������T��#���ĭ@<���ĺ��`���6
��s�D�<#	q���,���W�Qs��&���|�¼��<�s�XK��}ܿ�8�XE�.������5��ɧ-]��z�=V/*p���k/YKnx�m�FXcܸQ�hd���&�TR�ݢ|?��KF�3�JUϛ7�vյW�͙��asw����3�A����3'|a[sr�?�Ն���\��rID�=v�|V�)):�%Mڢs�Vd���?~�oC���% )td��b#,��2L��b2�2W����_y�����`6 6_�����{�2�`pEVi�xOks��=Z)��B��b1_ ����Z���[�aWO;H[�M���`"���q)�P3zz�dmg4��馊�@$�Jf�55�k���ѻ�5L�zʪU�f�2M�3&E�l�*Gg����>��TQs���|*x$��
#Q�M����p��#��*��F"Г2�7`o�q3Q��=�΁�9E�@�dBv�P)����!�TT��[K����R�ߚ����o.\��C.7���������f�^1����˗/-��	����bl��B�,����R�cIH].C"���l�J}S�N���@���=�"+�FeMjHy%�/����˖-��j��ljjj��&}OwG"�F�&�����+b镓Ed��O?�&G�b01`�)g��D^Y��Ҩd�!�l
����jX�d6Z���Ⱥ�ȵ:m�Ό�֌�!��v�~�LXHw�qGiI1�&�3���+�-�jMVN&���۷���c��d�-���*Xn�豱X`_t�|r.Z�e!e��s�,i��i�$N���/�z�DoC�	��Y��u��Y3Ϲ����sYaQ��hZU��\�PP��%��>���Z�ξ��XK
K�=��� 7K�rlJ����}]]�.���>3�X����⌀ƚ�k�l�Ʉ�h�k�A���:�RI�N�QS�tJ��1�D�`�F�U�u�T������3�nl�A�2����梉��H���n3j�of�0*f�����H&�F��2�Zm��{34٘?@2x��͐�fu`L�d���?��UՀ�SI�Jg��T[-��)�+%�T��4 �JR-�4ѐרN�a��{��;�~��ge����y�u�b!���.�LT'i��������z:)�f�E_�⁌֣G �"�d(��� (���Z�fR=fO�E��T0�G�OrL
F��Z�3�Tf����z�E��S�b����������������7�����3�y��JU�Y*Ͳ$ۑ��8$�sH�k�@�&4�xҼ���5Ёi �WC�vC Ƀ�!ǎmy�m��y�j��Uw�����{�sꪤ�a�Y�ZW����������y�{9���z̝���f;hu*��I��ə��j�����*g8�/ξ�η~�'�&�c�&U��
����ű���O?�[��[�����D�����y�gRBO�e��M���rI�7�c����I�7��_�����S`D#�k�Ԃ�Ė[.���#��
�{�봎�;Ei=�c�$���/=ztxm?�!���M�Jn��֥�2e�k�h��
N������)չ�/Vz�7��]kq:�n�٤u�1h�^�ܬpM!�}%�����9wo&w��G!�����oU�Iˇ�V�:}�}���Cء�.,�U��E���y�B�]�m�¯���K^x��Ե�����v�z��S�tj]Orh���3_��ݲs���kg���r��)F^�T�V�2y-l\:�:�	B���tiΝ�<�Y������?�3�������z�C~�}�صV})��7��C9l����@o/y���ܙ�{����޾��a�܃��)�J#�T"�S�~ c�k�b$l��� [5h���w��Z��#�!�E��K�)��)��ߓ�b��O�l/�n�?( ���x�`�ʛ�n���f{��;��5==�!���R�(�h��;�e�i��}���d�BGl4���%|@�m3D��B࿾ UԘ�c!���}^{�5���� A��HF7�U���ƂP����ߐt��CL��C���ULX�(\��������X!)�o�+2��׿���~��!xǎ��0'MT7��{w����+"P�K��D	08K�g�g�����O~�<������BH#])5�ַ��ڹs;�������=R��l�"!����n պ1c�;��4Ԣ;�N�7�7��~��#�H��,�$�yI6��|_r�?��OC��:"��wj�r��/N��G"N��kl�oM� 1����n�I�P���`�*E  ��IDAT�����G?�џ���7L�����^X$�t��T��'O�q�~=�N����l�Dua��~�������L&%oG8�F��UEc6��X�v���ʬv�@�㧛f`�a�=s�_��_�_��oWo�}�w[$`�ti!�Ŀ���~�[���2u*W)X�12-h��]'�p�E�9�SS#k�jV6p��������W�qV��b�BŚ1�ۿ~��`W}���b��w� �{�N�O�+iN��(*AL��A����ǻ`]���'���?��^x�K�%�QŔ��:#�c"�_~:i�����⻂Z)�?0�9}���s��G��v�ٓ�d0g��{�%B�ڲ����ߏ�VA9��!�`&�;�� ���x	߃�`��y�}����?�cЉc���xꩧ��^����	X�B����,�������o�.1x(����-�攛�b�#G��B�j;T�v�,uTq��%�q�=�A���G��ҎH@���"wWz�]�~�ד����+�������p�Ba���d%�I���!����7>��3��WA�`����{��k��Oم���<�ljÆ�R0�/�y��Ż����3o�f�.J������
ӏ,�0s�kO�����׿��C����?���[ϟ9s��"�uurJjh��T#��}��T%�"Nt)��&�t��e�W�{Z����|	!��,*�0�j)�]<�1	q���n�%X�W���%�j�Fy�ر]�{*��|P�s�ȷ٨A�8������LP�`�R�P�;Sq�zj��--�3�%u�n�j��*�It�u���3�aՋ����2`=��"�bqi���r��	T���+?�2����� tO����� A� �<u������A�*��,�����y��C؄���EGХᅯwk<`y\|�H��JV��M�	ZU��(�M�X���`�A���>����R�/�jxM	uc7��?���|��G���o��)�Ȱ[����c��;�k<����wp����x-z{�Q��2��[A������~�����#�<���|�P��g��n���~����ԧ �8�OEkb�K)�m3r���p���N�{�,�'��2���5�DE�%_*!\�1�<�^�����:���}�c<x��G\�XS|�۶?z��H�Ew�y�ҳ��������'�"t3����Y�Y2���>�i��;h�6W녓�sW2f�X��� 洢�Y��0*��l>1�Vm�(nب�̜z��e�þ��e�҅T���hf�<{�2żLgffq���3g�4uJ끰�-����L֣�t_ٸ��J�t.Y4�T�<s��Kf2�j� �И�e�U`1��K�͕IM[t������]{z��WO�;�{O>�����ϼ����{��F��u���n�۴2rٴ�cL�{�l��<K5�V�����'�/}	GpE;m��C6��Q�l��N,;�Y�n9�6h�5�>D�ւ՜H�,�����_��O��o��o@��%�����DW���U����5ͽ:��sb��coLl������qP)�n�ZB$����_��_b̐U�D����rm�(6����FW�ե|�2EH�����?�04����}�k�B(����zqܿ�^�/�w<�Rw9ᔪ{2���������z�����KGȍ�m�5}B�0��@�܁=G�ӥ�k33��Lvp`�0�ԵOŜ�e�\�z�|`Y�r}fa�Z"��ᑡ�k�33������Z�~���3-�R�;{�q)w�cW/]87�y��~�8��羉9���.�y�5����5Hh�)�Q&�X^Z̥b97D
�^��$8�X{_�CW��3���3�?�k��m�����i��˗.��.����LM��k{�����"(Vj�q+(P��c�E1���'c9�J|�s�A�R</KL=��)A�������eUx�L��CIY�T�nH�R*�������2��P���(VAڴ����2����(���y�I�L�*A�����-�UxK��%^@^E���쥮,>�^[-|}_�R!����K�nn��hC�n>2�7z�%u__��6:�x�:�R (k�{�`6,��}��e��uR_ݠ��|�l�Ug��%�w�!�6�U�ء��ٟ�����~љ�� .�̃d��o����_�R�T�W��C�=�U^=����*&t�
~|~��f��P[RP}`�cT����*�N��E�ٵk��

f�@���|�� R�%��R�n�ю 18<$}��W�]7W�o�\Tl]r8}�4�����ٿ~Æ���jmY�=�/�r4����p��yh'�|���Mơ7@Ӆlc8���!��L3�F�e�.��1IC����8$�բ1C�P�K�����|����6�=|��޽{a\L�5nO%�x���X�����tڥqI��.���^,vj"z1�K{WG�t��&�=����QHls_����֭c���/}�����/�#Y�n��L��e�@\��[*���Ʉ���]�c �7秊�}O){�D���I*bj$��93Y��2��&l7�wM2[}�Q��{祗^�Ї>�?��P�,n�ԙSU�/��)ow��Yr��D���m޼�� y#�9��������l.G=M|7�4��JK�U��{O�^�y�8ż�N"29=�(v����n��'0x�,����P���ի�M�[C��j�-ʴX����s�o�� N
�DU,.�C��K�	�M�@�aq�
�#0�φad���o+�UOI��r���$biuS�P�',��4����~��[����/�)�w��0;�m##��sG��u��];w����ۗ�
ҁw0� �[�/�=�A�ӻ���::*�.�ʎ��橫�������2G�TL_)��[ 4A���߹s��G�+dɥK\"��^\^�)nq���T���n�{a|G��-	�qg���b�G>�S��$�9<�^(�7��q�+���Y�[
#���6��z4�����O'}O9�W�5ۭ+�Cy��D���)�}��5���Fsap�r�.u�xy��ĝ	����Mp��s��i>C��K�����h��P���e�C����6��
���	���H"�I4i^���������`7J�f��j�fP�Dp�b��Vt����BO�:~jRŒ,`�y�뎠�%�iF����[�������C�
��MM�lذI�W���Rb�ࠤm^���U#	mz	���o'�6�J3����d�*�0Q��|��C�B67���Ê�L9�U���s%���_�����-`j�&�}���g�p���Z�������ըJ#s8�N���'�c���TY�v�P$�C�@6��8���/�n���*����M��>�9q��wہ���������)u�}w�^���Ԭ_�cK-b$���H�̹	�J׵��P1���5�>V��ˁ�F�)sʾ�ːF-/h��:#k��5�~��䩻�v��-#W�������0,��kGΞ;t���t�w/��3��48��RNE��f�:u�`�cj�nb�2�\��&̕�Y3в�`"�v]#�1���j	C����}C�~HB�����d�/����c?�c�7m:y��4/��X��S_�$���{���%x�/~��˿����h���s'��Y�tO�v��۰����c=�#qr�}D�-ҭH�2S�zŴ̭۷�+է��֫�_�����~�� т	lߺ��7^�e�Tt`FqE���7�wΟ���?~�G[G�=��g>��_��.�1Kr�ih�v���K�64���i�c����b:�B�U{zj����۷ow)M[�܇?|��������[O��LjXt�zeyy�|����.t�F�zd3�]�=�lV��Ξ>mw΂ws�#Ȁ�{^]�,^ل�MǮ�*�W�'������:�gU�fV�3�l�H#M�uW-g�fn�B6����sͱ1�u޷�Z)'��33�[�����Δo��΄E���
���[?L��/<(�C?�>��?���}��/B���B9Ⱦ���,TG=�)���:YV��i�i�UJx���<��R���f��X�\"4�m�KK�7�|�O��'~�w��^�9k�?>75n9�3 -d�Ή��#���Ui�	�%��eb��w|X��p��奡u�^�����$��R�{���'	}t�5v&��M�]�Z	��rp.+����;�M��H��LF�OT�9E����R�H/�|\599)���Ppv<ECA�����|u[Bw�/���M�M�.�OX]�SVOo�Զj�8�b�(��n��е������l�z����7J궉刚����~��܉�����C����ϛ�6�;���cZ�N�d����D�zQ�z|�	ۃq�� ��Z�C�<���i�#�5�����͵��~���O>V���@� |x�7�hOLL��

f�iK�{
�{JP)4���E��:@ۉ��n�*y�*2���Z�XH7-0r��+�ւ'�|�~�0���i��)7����n�pO!ΛJR	����Pئwk�f>��1�֧%�o�RC�H�&I,#�6Ef��pB��[���Y�t�� 0��o�^�S�m��v��b�<_�݁���o�M����٭/H�;�oV�^��i4��H����N�kW#c��:�moC�
�)��!m@��(��(��'6�T���m��� �����y�_��_���=��(f�� ���TK������~���'O�>�<=����T=����B�LO�������R�ÁtS��zXq�)P��q7o��;_����|��?��?�G��#C3�r�W^Z;��*#�e������ݶ��x�g?��x��c� ��:`�1H��*U �0�U<!6RU��1�

�/���|�ӟ~���?��O�عsӦMo�����1c�6�LA������ڹ���ЬϞ;uJ�����r�l+A���piYI�NW���K`?R�F�M�فإJ����#��	i��1�9�I�2XY��ڱX�}�]�|�ʵY�%���>��3�-WJ����� Ο>��{���կ>����1�������S�MBc��+eS�f��$cN�u%T�Q��
8�����K�iO�Z�'?�ɇ~��[�޻o�0EΕI*藖��Z���x4�+n<I1�m��u��/^�J:)���$Vߓ�_�3wcYa.y�؃
��
���;f�خ]{����s奎��-,.��0�f��<۱;��~��[(M�LSA�o��T�H>�
Ed�FOo�X�sC3���q�j�*-Bt�HDw+>�J-)�c/�'ҋ�p�KB����ħEǍ!9ڭF7�Ŀ��3`��Yr�	�V��JR])ґB �+��+��'���Ǌܭ��M*7����;h�4��B�ԍC�q���GjI���4�b8��ϣ��^pbW7:P�|v���8����Udjh+����9�g�380 1x�¹�g�doŞ.aߊ�Q�D��	��;���Qѣt	˘)��LH����4#O)��~wI�$D�_,-V-+!h?��
�Sk֌����2��BippX:��vgtd+�S�g�jzj&a�[�^�+͖CO6�<�^:��#*� Ndȼq�|��ߏw���Y&�vy��Z?V��ͱ���NY꥜��B�+c�GFF� �z&��}�x__jyi�����u�J�S-�-XA<��m�v)u� a���
}�]K*ٛ��"�G/\��k�����F��iݰ�ԃ� 
,��}����<����
�3�B�Ng�����>��]�.\��T#�k�/}�[���O��'����|a~yǎm�SH���\���@ύz+�+�Z�7=���h>�G
ʑ�{�C.�t�u(�FF�	�rV�W|����������N+�J��\���c_z�����>�������~��a��X���	���?t�¥��+��׾�d<�S��P@H�[\~"�L�-v��֭U����.\~��qb�����/]�$��wߩS��^@J���ڷ��<5Fbr�َ�Lk�[�D��{�����7�1������N/�Msd��Xn���&1W42Gy�j���s�P_"���ұ�46�bM����؀f�ۮ����'pN�=�nʲJ�ԼF��.��:8�{|]�˯�A�o��[��X�7����b��w�y��׿����?;z�����Ri�Ry�ʥS�Za�ƍ��;�F>K�J�Q���©�o�LV����%{��wtv�s)&;Ђ��T���H�����ӧ_��'z衻��ޑ�ҷ�^9x끹ڲ�k�[�رCl'�\)ٗ��""v��Z;����9rChڶ]�6o�r��Pnd��T��!�ݍ.#;��S���a[ܪN��"�1t��u�;��kCA��^������t�"�'k7o��.]�����������Y0����`��b�1�����~� �^�ԏ3�o:W�T�w]�)�
B:�^z���[��W,e+�p���R�	=����T7d��h���X�ï"�\ ����Pr���`12�$]��]��'���a���6۱� �F�����^��S0L�d�\�!s+eNr�P������)��a�p��&�ܼ�`�X�&"L�񰱩��a��A���s���	�%�q�D�d`�7�P��e�N�.	�k�ۃW����M�@<+�����?F���szZw%!�w�\���Cwg��P�!����G�Z���L=OT)��v�ՁN�zz��Pjg�T�S�k�$�ɮ��T|F8Hd3v�E��m]G���==�W��okZ�яU��^p)shp�����JGs�v׮��>a��ݸ��d��T?C�'��g>�j��{�N��&4b�k�N������y�<�����%�w�09��n�ݔD�M׮MQ� �#p��D�l�`��l�����zP��0���{����מ��׭[�������O�9NQ��[K� e,��X�O�Ru�<	i�ˬvs�j<�1«�+�,�{���I�lh��c�=���c���w�E��� �J����.�N|{߾}�duqa�n>X�"{v�Ț5KK��
�!!�M�z�+�t���%�E�^w����`SD]o����P��h���S�!H��y�������}�+�����Q�\�G���C��e�������s�̭���!T(4�{�Ѻ���X���ÃTOa%���¦b���حH��Ѕ���H{[�n��C��|�ۿ�����{�s��Wm?�w�H���t�8����)vc&������
���v��h��EA��N��ߓ�i���flT�-poP[��9��A.W�Oyi?צ��e� `�C�������7k�j��?j�j6j��e�,�l� 1.��<'�i�����_�K��m۶�>}z~��D�c�l]�1�G�@y1s�f v����ʒX2!	�M���*f"e\�_�����=q2�YI �a��4o�E�KT�P�B�{n�Hٮxk��ɮV�ӾJ���
m��A1#�$pq$d��+�PB��Ebɐ������CB�&Gn�-��y	|�I�ץ%�E��T͑	1,-�RF�((�i���|�4�ʏ�-�B4�$�$QK�AZ��bl���Ub��X��S�֒�w��C��̪$Ih��h����٬�y�,"<����%�9�C}}}P��%:V3⛾��Č��Ry������Qo��R��e�&pX����a< ����B>,���M_MR%��;~ǵ�m�߆P��O��1s��&tD�"i�`���v0i�F�H��ڊ�8ߡ䎄"�ְ<�7k�;M�2�==�f%�J.�X�V2����ܹl�eTl�6y��I?��ʇ��4T`�wNk�ںiuΞ�ҫ�7�f���'���-\%����{v��wI{�V#�i�Zm컅�c���lתMJ�v=�E˴M��Q
�mR���HJ`�ˋS�Ú�5�N���q��e?pubF�E�^��&;?2���u�g��;��l��$���KvK�Y���n{�g�-�(�:��p�e,�zΦ\=a$:�U�)g2YKU�.-*���@�X�$�֙S�׍mY795	b�گ����������0I�r��%'pL HhfЄd�
O�(��D�9
S��y�-�\�pA����!2!�񙼏�g���w�=��4���㧯nY����\H��K�K4	��rkbbBe����o�A�Y�4f��`��T΀J��)Q���$��C6���:�dL;��Sg���t�12�Ui5Z�L�`_�̬���Oܲ����?~briiY;�-=p���V�����u���@�9!� ��:���./-Re�OB�@/a��ښi�ڶxG4ݤ�F�$>��d�� /
�D+��(��2U����.�e(5�����..�������_�������s"8��ArC�`��5ǎ�VOXe,�QlŴ����3�{ד)���d/��b�5��w��FNh�w��ߓԿ���*I2d��� �$��d��YAW0����Z�i�!���^��­ ���)�Y�M�NԨJ�ʹ�y̋e��*6����|U.`�5�Szm�t�n�Ў�"��'�ؑx5)&�v�s/1���-���}KE���rs�:iC,@��UIq�a�܊�?���3^EDc,}5����V������^i�D�{q#%�"I�9]�/$�,S�t�Z:̊����2�F�9�>C��@�PlŤb��d��(^7������䁧�<�Tr�P�Ī�|#�uVM��ד���
�K��}"�YM�E#��K�%7Gp����⿂1�s��b2[͎��`�k�*���Mۑ�`�q����4~W�B���۰0"W��2u��d����v�s"��v�2gc��w��'��D�[� �p���"4H+���$2���T�d�Z�
[�7:6��׾v�	�$w��vDץ4�����HDRM�_���w'������9u|�q��b�ε�:gk:�Q�*ߟ�k���Q��ʰvX��`$�R NPIY#|+aJ����N(/��熸��섓�fcd��hDY��+O����N8���
�IA �����'����)̙��cX9��_B9�&@�����pQ8��Gz-�^u~jj��p{2��٣�s��w"'-J�U7M
��v�E�-����09s%�:�XI1��ss�<h��n@�/��σ�/�5��*���<V��8Q]w����o5�I��	�}�ԩ����;wR�M��'���˗�p����ċnw#"oLش��0Lߌ��~����d�p��H}y�?�A��ہ�!�>2�v��T*C�s�Q,��m�$/}���)0x���p;�I��Gk0��SH�Z���g>H�l�	�����E�,�(��s��C�C�ĮY�:n;����j�E8L�h��`Y%3$�k͆��X��pQA|nC���œ.]���b�k+"*D7.���	�x�b��ݽ��2�A��L���_�T�]Z?t��>�1�Ѝ �sBds��G��=��@!z����������`"��Q��q���ED�E�"d�h��/����]�?A��|W�!i������T�A��P'�B���a#c@�lA�f�Z�)�8d;�y���X�	�_T�U�	�$>a�"���-�������y���v�\�C�����m��a&�K�f���X�i�����S���^Z�H%!MQ���2�;��W,W"��(X�&�2��\��~}2&W�+���M#�J�(}}N��H��.��b�#��1q�1�%~<v�NR����;ۏ�����'�~��ŉF@�{��P!��n�z�@ �k�GȱoXo�̡S�V'I�'N������ޘMk�L.�Vg#{�d�����-�^9|��ѣ/��G�`����H�ɷ����+j����<�<1�.:�X7Qs[h����(��	��q}��/�F֛E�D�b��mZ$5��$F�&����{6�7/h���8wR(6a�̤�(f3��xx�!�)�� ��6{d�[��J%|?,����}�m�J�����JN+���<�c,ު��Mm���+�������9jͅWƎ����\�8nO������"N���5�:w�\���d�3����PJ�5���#>V\ӣ|�܅gΟ�H�P*�=dM
�ŞQ�<^6�nB�����χST�9~��ۚ&���2�E�v��}㠊�.sŤAn(��"�TQ`��I%-C'��j�V��Z�����[��L�_��a�����g�)��Su�(�����n��U'�N�^��=�[R�a�J}/Nc�!Y� �G�%���m��B�*�QV�`	�M��zm.w�|�m�nO���ap�jE:J���{1�q+$?Bő��g��Xj�r:��3r�H���)t̑-ҕD������v�Z�t��r $�H=8���;�'��iO��uum����B�܉��uk7H��VR
p24�w��q�Ak�_%�@�c�mڴ	k,�7M��%�����c�Ux�/�<��ׯ�HHX�17K5_&A�QF�Zy�|:ͭ��#u���@H��b!B����b�r��M�X�f��D[,9!vɈ�{�L^VPV�"�,�rCl���0�N��F��A����P]q�X;�L�╣��>9G�i[�� rlT0�8�����ի=�>�U�Σ�S��|�&�?>�괂���gl��(�"�b�u��"�|�"�CnG�Y�*�W��b�#gr��wl�)�R]O�n�$�߬���J"�bklq��rll���I�	��"�p�ؙ�Ǐ?�����F2���a~�).���#~�C��kp&�%�_<Ur@4�k���|ː�D"���Ѕ�l�A���ׯg��:w�nQ(6.�d)�(�V�Z��52`�W@/)$��p��t:%]6�؜����B8R��I��iZ~%	ΒtzT��v;���axR<,�W�-�bL��W�����`@+uv�aP��|��Y!I5u�4�g�kl�y��K`� m _ś��LV~�SEw�n¹��.A��I��?�:==-S'Yr���\I��] n��B
/�y-L#w�А8w"m���
�Zh��o��W�O�{;`��N�됿���Ai�W�툭/my�ď��"�4���*��e�i*�`a2}��64:���f���݈�:�n*����u�6�J��L�J�ێ���0R����'�b�D�!�"NZئؖ�E��u�݁��֪�6�(����[�����E
΍���GSZ_�2�;-6y�5K��v��^�)�]�Ԍ����G>��f��4ZT�8>���M��ZܤX���o���	|�ohhhǎ{��������������l?�{���5#2W�4����kצDLP1��h����js�e\�����LNNf�J��+�j��d��%~����*J*,*p���j����7 ����%��ߪ;s-*��Z�߲!����0��0��Y��T�vY�D�b/�r|]r���J�+�_�HY�i�SF������R��_�5] #���5bVkDȯ�?�8Ꭰ �Mj�+A��gο�mo�ڇ1<��n
�?w�,��]��ßj���$��z���D�k�V���r��>�ڊ�7�JV;��8��3�nkd�a�ޔٽI�Ym�#	h�UDv����/�w�Ļ���B�@��Ǥ�iCif ���_�1R�I��:�&���J �	uA�W��ƞ�t��ֆ&�@�������!vAu,l���t�SV�����XjzڭѶ���v�s�-|�h��B�DB��H��I��o���a'-J���K�ių=Y�=����)���>��d0,̲�ñ�b���s��m�����Y"Ů��_�:A�{B�U͎j5��$>�X�6R��C�	���TZ[��ڰ3�=sU���1�U���i$�b ��'xMLMa�S�!�p*�G�D���^4�O��Tɡ�jeI�eK�3t�+W��C�&F��[�U����U�y���@��!��b'D�S.�K���2��Bv�@��[�N%I�'�H�4�������`�+�[�Jfm�J:	�H*+G)���@�cS��J6�4��C�9t�v��PxH?�Щي� XuM��A6���B�5 V�;��օn(Q�}?&�I"c�
�T1�&�߱�v��9�~.G�&v1>'��a����x0��*�^p����oJ�����Q�[��qu��-_���JhI � ���4M��w�:W�kG��LL�*�!���Yݲ������B7���okZ!|����&K���aZ��״�d
�㠋苙%)W��R"�8 �	4-�����ҙ�Rl�]�N���>��γ���Ν�rU|	����������㵘qho��n�\� <Ntd�7�T6W�8>7��m۶�2E�B�-[�l߾]�+�k���xn�r>������-���޽�yQ�]��9� C(�G���G��7���U<���7n�_~�e�]2�E�`���[�n�L���7����V�4�<'d̒u"���:��Q��l�،��i�p�8�/��c��ʒX��\*���$'-��'N�B�@��bH���X�Ũ��$7a�rm���y���W].8ѩY%GK�]�/��]P������{�����X�cǎa2;�E�(}���%����wb�@`���7.�}������ܼy3���*�b��M���82�n[Y>�%3��C��n[�[��
�/�\+��#�]����wI#���Of_ɥb�c��J�Ғ�h���Ț58�Z[�x��ҢzX{�С�����S�|T���5;Ί�:ZS=��Y�n���[H�C��
s�HX�gϝ��
����^޵c'vǾݻ���Ϟ:��B^�Vs���5�k�	�&��;$���9�XoҮl4����2U0a�x�g_|�ӡ<f��-kA�P�#�*4���WlHu��)S���(��A�w�>��۰�'`e�ȭDL�$�������1�����^}�UQ�-�N�C�<=��Ku%�⥗J�֠�FΤ(�ԛ~׻�57;�Ϙ@<��H �mW�8N�7'�����Dz z������	���'B�O���]�!�IC�T�?ƨ�5�t̯����i�%,.��2�v�&$���.GI&i�h� ��#L�ߡPZ��B�b֒������č�Ϡ
��CW	ɍ�s �g@
FȊ�㒢����������t��]7���x��Z�0�2��\1��Ɋ�M���M�@*�6��62�(�\�$�ܠͭЩ��*����+���1��4X,��r�0��jA�t�U�O���!$�l#��T������a!i��a�=��s���9���M?!�@Q\UbH*�Vٶ+gq��0�a@H�[�R��#@%���8�_��_�ˉM�łln�8p�?�^��+V�ŷ,.�Z�Ω�Ж�xRN
+�U:���z��Q�k�H�&죞�5cks�DE��342
��h�>1�n�������:K�Z�Xz��1�g�y��a���=���E�E$mmegv��c��c7�5�m�V_��A0�;vb1�`4`��:��BM�1{��}��R� �;�y���vn�<;��a�[n�EZK�����_%.����8�/��4[{} �Z���F�aPJ�P�7a����䯁�Μ�@��R�A�V;��O|�޶s�+�S�F+8�v�O|�>��@��%Z�v�moy�[�m�1��20����a��G���9�'��$#�I��a��wK}�����|��:�A�܋��Z��{lu�������iM��ֿI��F5�J��ܠ���@wt�1�#�e��{�)�}?����c�¾)Ўiel;/M��T-]���}�^`2�a��1J����M������Sf��0�/��a&���l�=LFA#lҘ=�C�W�.�k���UP*���Ե����2�[w�I}Yn� �����{X�,l^G��c���f��L��Z"(����v���1�t6��J5c�w`��į֪��y������[�l���^v�1U�U��S3���&���F� <�ҥKPs%9�d�|���)ʞƞ�%O>��h���gΜ�9L��B\ʩ�)���򕯼�����>��/~Om@���Y/� ��53�*�v�y���
���_״���d������W��^ӛ��`��	�y*)�s���li322�dYv9���I`��hEk�Y 䓢|���2I��ҥ��GC͢j�6�n
2
uS�F2<vO��1�S3�1�&gN���q�N�ٱT��,v
l�Z�E�F�*TT�1�1�k����⊢�0�I��D�i	l�N�U�J�AN(�$�������D6s-�rB|�[��%�[6O�kͅ�+bo�x� R_��؋.D	�/F�$Ċ����
|�up�JOlX������^b���� aLJb�lqKcpXIa��q@�b�֬YC��D����^e��d�駏=����?z��5��;�s�W�:"��U���B �=C�����`r��*H`�c�j�����L���8�<���RY�F0�ոd�&���ɩ����L���*�t��*U࿲@�>�{�����A�7�%����k�F�'�ٳg��$��򗿌y@i���1� N�`��r�c�/���/V�r|���s%�#�{�3w��u��œ'OJ�(�Y��d��r�K1<<��:`$оq���]MF��ĵ�.:�&��)��'-ʩ���wc`�5����}���~���ˢ�H ��?LPt�UWI�?n�72�Y���i�x�$���`2�q?p���&���۷�ܹS��e�x/A=*$��tۭZi���qIhp]�ƛ����"_�*�^uD$�:A�;lӧ��x��{���'G����h�NHe��a�&R)��q�b�P��[�媩����J�!>`0LS�6�C�L�M�}�y-$?
EJ��o������M�p+��-{��t�֌b����+����<.KYx��5�V�^���7�$;W�^d��.���F)`=@f��Ͳmv:�dr�Qe��D��ܤ	��v�^��Y��Zd h�$pR(�@�5�����0����8=�-��sՌD!U�@���K���?�#?��C=��SPDٍ=I�A\T��b��������@wl6U���{�#d$x��{V����*��kZ�<
�C߭�$�Ϙ��?ğ��Os�KB=�$=f@��y%M�ɜ0-65����4I�*ѪU�V��\��nF���'�g�+�ȣe5�+��UK��u !���9X�d�f!+��H8�]R?q�è?锬��8F�`a�;����z�x�{ԨKery/k������N��5��J[7��0;��Ϗ���K��Y��dӠ�L2��8N%;v:��F��Jf`�f�9h�L���E�N%s^V�=q����oXE��4��57�+�..�g���B��HG��#X)r���RX�T:���t�����M�����g.�Y��\�ƻW���j{�L&oj6 \�/ ��2�B���zJ}��)�h��	�]��*��z�r��X�j����z��Dr���ū׸y�^oւ�"�]+�$�+kӶOz�ḏ��ȇ|���/Y�Nk8��Z��K�{�� ،v�4�����$[Mw��[v�r@�Ys�k#�\�B�nP9����4�f��W�f�y�%,�ūS�xǃے�5&JC�׎���t��He0l�;
t�v*������l�5��~����'�k�J�6:�	G�^�E�zA�ުVhz�t�ۈ�]�5o�Zzuj1_RF�Tm�y�����6=�9ǻ�?s~|��O��O}��d�[�G����k��NR��W��w�ܽa��n1���N�!�8y㝚�����*&&�o� ��$Ñ�p$�z��z���8�W�	w~f~Ö-w����rCBB�Pʗ�8��Ɓ�Oז+W/]�����s�Nl��ڝ�͛]� �L���j�ҙ�����ŝ;���_W�WR��F��ɦ�
M�ޜ����J�n�8JS8��M�,�<����*a�U���4ӢH�x��Z!r|e@*K'k7,ǰ�>N�W�6���ze�����	��h��R���M�JZz3�Z��RSv2�gӽI���S3LF�8��`Bn����x��9"W�#ð��Z�񼠎�E�P��	u)�J�K_W����&m�l����i���.�ٷ���L��m�ne���d��e�Vf-��0�Ng2iv0M=�^:]O����j���w�����"�iCC�ٜ�8����oS%�J����|��Tc���͵��'6E�U	���i�ߠZS�$`��ks�����Y���+��o��:y�u�5c�f [*��<��B�P�O\�zf����f�*�c�_��ç!b���S.3��Oִ���Փiä��D��#}��)�\ҹtR�\�8U�3�)����7������S_�җ�����d��G�l�P��T!����*��
�`~�<�,�?c7�m���dZ�k�~ݺ�Z��m�J�������F��yWvR鴮��B�m�0����˗�O�%!$(y��(CJ�����K=�^�,�ށ�p]�6�O%)%�S�,L/�G�^?�P���S �.�;@ṁ�h�k�z
d�͵��r��/I�&L����l7:�So��媊@s�L($af��lQ���^���a?ձ2*H�F?�l^��t&���4{�z�P��A�K��iX���$�&"[re�]cTn680
3�u��/W����;p���y��J%��m�sg\G5E$�ϢnKtS�&��ڢ0KmE%��֑��)��p�ɥ��œa ��@�r��_���(���V_1`�/p̎K�F�D���eY4�dH#��kll��;����yF�TZ֩��%)QB�/]�4."o4Z �L�#���>(@<H<�Q.� �Zo�>$ī�f���PT+y����a���P���J�P&�]�(�ݻw���o��o۶m��.I0��x$pHݡ��>$��~�5YJqN�E��x#uF��qJ?.+��<&�\�� ����i�?=I�%Z��JzN<�&}��`w\F��X&<�J��o���sd!�###w�uב#G�����ꫯ>���=�>�"����&&&�,��jM�V����ŋ��=���x�l�����&��E�[C��$}Iqsz����<9y��q�P�vx �s
��i�6l� �A2���?04*��U��Gq���=���9IN� ����ᦣݧ�ЁP`�i���I 1��iQL���r��ߣ{t):��i�
%1J�HQ�a�#�MQvɮ�ͫ��J����� p��L�F������F����5�B_�0�V[�e�]"l=)	�R����
�������.6&�R��L�6����&J}bz�Y�:Yl���y)&b;��O��䜃q��@���%2=�r��cd�*���b�--R�țo^�JQY��*h�UJlD]IN�鐮�Q�.e�����/)M�k���U ��cx���J���㊧G�L<�c�l%(X)"U]7=|.>���kQϰU���5BW��Te�-]��-�K�lB2�/��>�V�db��܇�c�$R��.�o$�ɓ��h�aŞy]��f��k�J�p��pOI�� ��ʁx4�Y�1_*{�e�s�ǔ&��&�@�@��w��7N��ᏹLxs�&",���`IT	>�k/R*�-8�>�f�Dm�H%	Q�S �k)x�%ʁ���EIy� �Dyz��a�H��r����7�ٳ�gh�F��# �&�d���@(4�-��i�B�*�T�7��j7Ξ��O�;v+�I�Y�"��@��7��R�Ezb�2O�΍�q^�$�HH�CЈ�^��bi���==<��z5��:t���s�X��6���s�#���'�ݾu���bOI|�CEˋե2M��I|OyJ"Is�^Y�U��'�^�/���֖k����=J�>}�Y[^3:�n�E1�Jeiyy���)_7�Jx�=?7�T^|
O�}�}���%)B����zz��}=�l'Ӻ׫3�ƱcG�-`ÖJ`٠�>�@� J��e�\�x~l�7.�#N�Pm�w��d�PZO�>���,���_饗:c�n��3(ޔ�>���|��c�=�-ST��,-yQeN3쥰K���3�)/j
���H����>|8���"e���O��$�q
?*z�v?�;gM� �*��0]��!�|*g_����/����p�~r��O��hj%W&I�hR��j^����C��܊����ܡԪ�ϥS HB�>Ҩ��\��!�K��Ț��A�P�hQ���;�4ݪR���L��B�m ���?��QHE���d��V�)z��=�J$��N�H~�dG����i�{�BY����T��!�GN��>�w�T���Gw�bk��v����� ��+�)���B�B����}���ֲ�	�K�#�E�����e�9�%���i�N���e�H&�b���0�L�au
�N�΄exf�cbæ��b�����O�z梕8����a�/��yI�s0�����X��c0��T�gHp܀���gPF��Ss*�\�r0�չ_Q/Μ#Ԇ����BLD?0��J�f�.�����s�Fű|�:��a\���s:�߲�\"�R@�J==�E
�a�`���^{ٮ7�	3 �a3��`���~'��~XʍӁ���ц��=\�0�6������8�cBe��N�aOJ��<jsZf%v�`q''sUMr�:0���q�t�o�v�G=v�L���}��9���PT�
_��(�tA�m�s+<� �cΤX��-��1DQ�Ƀ Y� '�6��|?�0ލo���.L�u��Ơq���>�b�:���}|H�����y-`� t-��l3��ױO�T�D1Ţ�v�4K��9�0��
�|5��>44���%�<w=����݂{�I	��t2A'e��Ո��ׯ�h�Kyǎ���<0�{˖-�c'���gh�PcH��p`N00����DB��2Ar%(i��<�8q��70��P�`��bAL��e�d�l�)Jh����d߹�,x�~��O��n�o� ��^�
jN��,/����	�;�ks[����*�Ux
�:�{�|pd�|/0R"+P\��?��P���
�I�۷�1�|�U��ٞ����������n��vA�';�q��K��(y 2�P#gZt>��#j��\9�X�v�S�H�z+���l�o@�nIV���gQX)�<�p�6h�;��L��=�hE�wo� �H���?@q_-��V��!i�+�k�G=~)��Q��jhx-�v���XV����L2�]&��쟜�:E�PTA�ԩS�Q�T�A��b��éP��m�����)ZxTPy�͜J�B�ˤ+7Ih���� ۭ�#�[6Ԅ��D�Qŵ	I\��T�,��G�G/Ĳ� s\�q�!�R�����f��S��L.����11�I�����8��3�0�{������������<)�`J���kׁ��<�F�n�:l7l�
H�8�����Pֺ�@h)5��_NO
B|M�]�]�*�ΒP#��\N)���8�T�7���L2�/�9�R=-�f��>W]ю�dS`�0r���c�f�礩�
8�� Fd���f��C�����枑:tM��'x_E��_���lS�R���6�peL�h�m�Y�V��^��U1߻zfX��y6�gC�Z���M&S}�GB����.(4�f� ���ŢW��B��fB.��RU:i�|��B|� 8���!J%�P�둯xl|l���A�Ҟg�����Vg4J�%���_�K��X�I�:�4T�0����nT\ ����ڽ��{؂�B����@�=�@۷O@`���k7U�!��Bn�����t��%)��F�c�`�M�N=ztq~7y�߈�cBճ0�S�h~�?�A�Ө{w���O�f���f���	jw��J�HzC�p��Y̳�F��P����[܀�&�ӓǏ���;w�fMS��'�����Ivy�"�@ۦJk�p)���i5j��E�H�nwZ�N��V�Z���E���d�zv�@�D����LYP�-r�௩t��i���n�g��Z �X�$ϋ� ��U��f>�'q:w�Z��v{��8 ��P���]�#��L�e@��@�\>*���,�3I݇x�p�<���XZ{�&M�޷���$3RM邃ľ�
�7XzQ%��N���a#˂��m�lը�$$����a��F��X����L��������Hz��;	Wx.�F����4rA|'?'4kaaSPdJ�`>W�1󦮂�N�p�UY�k�w�;�ܷeb�꺭����Q���k�NiB�GG�._�JCI����CC#����f���Ԫ��yJ�L[�����ut/I�T(���#,Dy5�l�V�c#(���y"�|R.3&�D��c���@
7ZN�D��7o��6�[��Vn�w���\����shIJ��%4+��,�����@��hw�P`����l`��C㻷�6csVD�:	��L���^�_p��AޥJ��L;k
���D"�ߟkJ�G;X�ԇ��M�D�//�L�d�f$)�]��$N/U*>/���}�(�Bxlҍ ?�� ,)@��Qm�nd�N��`@n&l�B][!_</E����Mq�?K`v���b��KY75�(�Xi��2B�8�UZ]�:�YI����O�\c��@��o����/T���Y�w�9�FM��pT�n�UKmm�a�v�u�,˕#)����m}���˃$ݧ�Qe��Ѡ�y1��׸��N�*Zd�tIA����l0M����9�d˔y;F�5�Z�F$�8�g���KV'�5$"]X�B	��	��D5�e}\�����vaVZ�kG�1�T����;��ÇC�K`L
��n�
�UBe7�b:e�m_�SA'w&���T=��P"Fzo0� �|� ����D�'lذ��n=�.]"��F��P1��hQ۷o��}�0?ZP;��x5q9�ZB�N��\�22;y�&PK����[-+���=�
mI�%O\'�R�o�2�1��_yE�"(%!rg\(���4 Eq;��p�PW`���<��̍�	��/�!}�QMV#�v��xY��%��ǭ@9к����c�,
^?.:��'Ϝ�d���#]�-��P�eRB@�����С�q�u+j����n�A:���F�	�%�\��vt�N��C����p���n[�[m��D.��?��ow}#� ����޺u��{�]�~jV�����6OX������H���8��<^gN�,���E��W>�B�����J����ZF�˓B��W:5� �*��#�i��G��� jb�+�U��R�#�J*	�x
�f��~���K
P�lǋ7aH�5�UN�":�wT�c<4�lN=i��6%��{�3?��%M��H�0Rv����Q����$�35�]´sO;.yŏ�|�*�I:<?L�4�U$�EZ�TW�W�Z}�$~?�lb���)����Z��-gd��k�9�Վ�L�x�}i�k��_ey_�q�i��]�򸕒
���_4�fR��1YˠL��,��1��I�ˠy��&	�NHx��V)[���`w�I�(�l<�zxd��[o={�
������~�K)�a�D� P�DZH���O��,��cρ�"��ߋ��㿽}���cl>����r�K��t��	'Us�ڍ�(n�)�-�ƃ�HzHq^0S`���~�Ɍ4.ŏ����O=�-i���+R�T��=�,��4\�	�3�"�ѝ�:���ǀAd��q���+�v�L��(�J�(�|&>�aϴK��R_��1ȫ��Μ��9�+N]��G�E�t��~��R2�jC.�R�-[��ٳkÆu�-Q�^|�ELK�20l��m��
i�,��J��lH�crjjph(W�|�?s�f9��Ô#y�:�r��E]*��vr*D_�6E.��ݸe�exx�	c������"L���Q�������"�$��M B*���LZ�A��d�,s��=y�d_rMo&G�ן�y�Ѩ���A�$n��ĉ�3` ۶m��"�t�#���Q�2N��bw�Ғ8��ʀ:-e%�e.c�Ir�
o�}��R�L
�('[p�<��'�֢J�����H��SS��-���iS�A6B20�siR��aD�(���+M��&�h񔊏�4��MwS�8l}�H4��F�oHԊp�dj�`�R XǞ5Ug�n-�{ck��9�rv�c��	K��k�D̾����,�v��䍎����X�=ڭ�"w�$����-�~촧֨JA���%3�w�ݎ�o�J��*x�l^~!�C��t=�j�)Wb�j�W�n&Sd��/��1��z-��Y�3����L��/*ɾ�Ew}��M���eo$���F���î��0j�nwȱ�L�-#��ױ�M�������l��yཁ����޸����:��`y�1c��Z�C>)�"��g�Z_���O�KX2�������Pٰe�	M%�!�Q/Ι����o��eI��9��H'	R�^ӥ��A��Ͼtu�r8�/�y�"�F�
�i����f���k�'WHl[X�3�A�IP��ޅ�$���G�D�C�c��+�l�c[��9��{C[!����z�r���\z�s�/<<f ���� �($���~d2�^Cl8=��l����7��d�H��B�)_2��G�����Q���$R�>Ľ�e��X��!�7��$HK�:FC�T�k��7o�_ +mt�Ǽ/�eSI#���ɮՒ܊���f�f0�o������R	��iA!���ʔ��� !.q�2�~W:�lj�{�Nt*ނH���m�&YY�}C��]�9Of��a��CFIFL�1��"�*fW��K��Օ�b A2L`rNf:VuuW���9�n�A7��~���{�p���{�1�w�_�7�I.G��Bn:�LJ�|}߾}F��Uڻw/Yl� $NKC:-?�3A�¯�*<1>�s�N��+�EJ��X�&��@^-�H��_f\n�@.is�����'�k�,G�9a����+���:w=6J�*��i���}J#욠>�RW*e��9%�w�����
ඏ>�(g�x�cΜ9+W���]�x���[�H���񺭭Mv\BN���P�&�
���k��F�1@���(L
�� ��g �-,�ЁC��ccc�xb@;v�,&��iӦ��ϕڇSN9�X�c�kx�~���L�ӕ�j̓�A�s�W��m��d��-	$1V��EK&�f��{w��=����F��A�Æ��� ��8�M��'z�
A��PHY��z�Q�]�y�_�jxI�T-�6�lփ���Y���r���#��qX\������0+�/ �]^k�5N	F��X���y�H���X��B\�_��U�ʳZ��!���vW�*l��	�%�$�&En4AE�V��R�Ȗ4��e����K�`	�`����؉q?���X�`ȶ��`�t�(VE[����٨-��ýQb�$㠸Hߙ�Lw�q<A�8�ٽ#�Y�(�2j�%���x��O�⣮0����+���MeU)���SgX���$�s��<�#)e����$��%S*���V��:�~�֤�ź]tI��j�a�I8GH}iCyM7H78�g`��������31��"�mp5�a&bm�SSJ�<�"��W(P���]��ԗ��וj%�(��"����x,M�*�<��%���t�P.�˱���L�#�X�j�Zq;�G��Bm�<�0� �{ ���l������p�U��,ӢN�X��˗3�4���C�^��imgђ�5��V �H{a"��kL�����j],S�0����T�˺�%2�(4˺�d;����c����*�F�A���u8-Q�^=" �r\�6@(@���ÃX�f�EkJ�(�������r��co�K!��cV����q�F�L1�qV%1���O=��s�=�k�X�;����G�y���ҩ���:����K1�b��C���U�^��Y~�����=K4:T�g@�.��|G ��[�����qW�fn�ތM���v��Me��=�gATϟ?K��K/A܊���֭[�%:��!.\(*γ�>{���/)�*���<�H<�F<c� ��!>�7S����)�	��~,e�捛6m��`�B4�P_�m۲��v�k�U��~衇�ÒSO=u|�2I�O���O�*�|Ajo�"X� 1)זtLF���F
?Q�T�X,����C2ƚ� �N:N���8�uu�-�N��6�wg(N�ϵ�\�m8L75�tʒN��(�F�#g��{HIPbۖ[��*�.��RX�c`�
O����֖T����Pc*AR�h&����L�����̷(F�R���pԀD׬bi*(1�ƙ5�:���(	Fe��E֪�+�78����b�Sf8�G~uŰ]��_���i�*˝�8�A�(�0�	�v�A��L��c��F<��C~�M��^�k�R�fH��\6��N�}��&�"�`�+��${�� N���Hl�p��D�X�S�<\u�E�i��I��S�"�P��i���9W\qxB{�l���qJ8/��
��?�>g:g��ciU	�w� ��i�,��II�D.#�&&�On1��\�`����6�f1��_U����0n�J�u,3Y6�)�".�&7����ft�Z�%}e�r���BQ�wv�V�K�e}��tM׫�M$��f,��;��g��T-���u�v�|#X�h4�(�:lW,�`ղ(�0i`�J2��Hk�nJ���sp�������e���I�����g��*�HU������������664��M<�IKanE��e�(�!���'r�g�&J�Ұᙃ�T'K��X��P��\��_�۔G3��jI���H��*v8� ~]QN���52�W�RW�$�����>��#;��>\�BZSKD\Tp�\������
%iڋ�T�8Ǿ��j
��X�4�ZP�`fK��t#/ņ�꒱=3�.�{Q8�Ϫ�n�����IR�@�E�(����tt�R��8�jժ��7赦�
�J�[�MM3��N7�F��Ν;�Є�Ty/�	�
�h��!	.`���� �R)p��۷����q��zp{��̈���ٳ��{���tɺ��A9��UGz��c��˫=�+u<�J�%*��j�$�y���
Ck�Z2� �)��ٮ5�����x��.Av�Y��&F�Rk�W�p?�d,�w�߼�aeY��u�
���M��$m� �N�3��٠�}�fZ�@�����{��z��nn�3��?���(u6t��C�j�ߤ��q�=�S�}s��y)͸�Z��r�zw�������If�'-��Ũ�w�����q^�-��`����U�8�@���iI��J��9b5�o��W2�M�����o�>oX��8��Y{�uD������KG��I�-
"��	I�G�R����9#�Y2�"$�,ۨ�a�[7�#�u����ь�����I��=<>��k��ޤ���=I��?��B�x�E�����yR�k�����j=X_;[wp���R�����h|�L���I�GP<̙0JSP��A�#%���ٞ�f����tttd�%�n��zN9Q?3�ox�86:*�`"���`⧕%�k��.��%��o{s,��J�7(<!SOt�hM�c�w��]֡Ԑy�\�ticc�r
%QSxx��[,.,������5��n�d���,T�J��DlX��r)5ug=]�b&;U��P�����Z �HɖW(O*����*�;���\g�`lQن*�I0!igٚe4ը���)�x"�aCU���ln�X�M2�c%8�##c�D1�����ã^%g�w��R��A�����XC�eSPÆ�P!���<Ճ�[<��쩭�ϓͲ�2`��-�˜l��Fe1���H,�$$���h��Q��H�� �*j�e��A)�6���[U�˞M�8`�"e��t`m'�Q�[ K�t8�������aԨS�ElG��Z�>�R�
���}�zE��D�!�ձ<Մ�"�Y�!�[V4Ug���k��ޮ��A���gQ&��)0���X��l���8%�f���D2
M�R5�䟣�"��`���(����a�B��R��1�)� ���E����E���h���oս�Q􌖠���σ�n��oڔ��r;9��]c���+�s�
 j���dy]Y;�Z�$8E�U��T%F��~���3r,��lA�k�G��tB��c�R�:�أ��	���B%�sl�)��2�P1*%%h)j-I��揪D%LbZ���8d��Z����ÛU�j�۴�ӿ��x1!ɉ�yM�����tU��:��?H}tT(�`EUH�h̩T}�b�P�
%#����b�?}�/�R�Π*�2J 'n��Z72�ǚ
����৚_��.�,wR�
�
K�Ӱ��Z�`�:ݽ!1ӭ��
%[���;v���m?��N?�����]��/�E {}-���pĪ�C�w��y��4�p�>aC�fp2��OҌj�V����Ij�ĖD۵F�~F3�݊��Ôņ����ʄ�oZ*� ���.�466����{n���,�=%.+�l���R)�wf�^�Ōԇ�:����W��uV��z�|�,]�4� �:uw��@��!v�SPsٲe�<��̛ׅO���siG�+�p5n��)�N��'��jr�j��u�(��SnD����+&z���}�͒��k��^7w��vj��iF��$�rj�m��I���5m������.K�r����T�eLuz&����7m��V�v3:�5"��B0�#�R�V�p��5ͽ�Ns��轐?��8E��_ �s����u�0Cآvx�Uk3�/mK�A�pzo��i��W��պKQfR�ik�������}��|ƪ��c�;�a��%�_T��E���������ʥ�QhD�����Vj�:30A3�Ӻ\M���;n�ޙK�+9�Jͅ����d`j�י���Z���*]�p{���H��sF�k���pwjNg�{yގzG6��Ŏ71���7�ș��ڤ���G/�bi�r�N����T-%֓���i�o�Y#�����ǻ�R�v��䑍�g�z>oY��H�x�I�D(�RCda��	����p&W�9�g:T-�OD���yE9Q�G[fIA���:\�L+���͢����U6��*���a �j���)����F-�,���@�\+E���EK�\{�۶m��m��K}B.���a�ؑWSS�H}iAK^8�߳���0D��_Ե�8a��D��Z��� p.旜8?��̋��zuuu%���W�~��W0��\r9m�k�0��{������/b��ʥ��Tu?���5�dVH�ʆ��Vݿ����\�=*��|�L��c�M��uvv1N�����m�[�lihH͚5k`�pmq��m8��8s�[�~@U�8ʹ��%�9�h3nR�f�:5D'����H�D,.���i�Ȯ���ݻv���)_�hefPS����Ư�i��BRǫIwP-�3h�+6�T�.x�!qD�)is�ʴ�-�.e��KZ����WB��[�b��G44�DQ��'X����c)���c.��C^&��V����i�,+3�Ek��@���y���c�TLA�B&3N�P�'�T�Sr΅iy3�S�f$4_N����q6;8�.�g����qt�/�T+ᘕj	V�B2�]�d��>��Y�LQj��
8��~X5����Lr�&Ý�FE���]��	E���w<��m����'����� H��J-��Tzn���q
��[�֔�5E�gP���M�lnz��A�� �;�'j��I��ෟn��y<��[��(u�n�#��ٮSt����6Pغs��I�̘�U��K}9�K��*���Z��J�@w��v�l�5�^?���UFk�D*�W�k���q���U�LkvmTR��J2B(q���&a��b4�����ZV��DC ]ïP�	)�
��Պb�ўؠW8�����<*��l��o������k����-�0�0����W(�@/�a7�4_U	��P}�oڠ��Nn�&+k?Q�T
Ŋ��p�[�I	�ɗ���|(#��� r�yYB��eT!crOi��F>�[p�@��a��
�x&��#����@��\��c�?�DU�9.�1I:|@���˖/���۽g�r�_�z3����QJb�e����}�1��}�v<cşB��L\G�e��B����4J-k��Y���1
/�"�(�e�c�*��'��a����n�.]��~��N�T�@�H]�1�Z�re��g���U`eaO��k���0ut-Pg��H}�k�z3ƍ��|�4��c~��'�|�+s�̩���I�w׮]R��k���:Pi>qy�bs]�,�����h}�MV��vUo�x����1VÓ��B��>=����9g��0�x�1N��� ���,X�S�B�O�7KQ��,ɢ'Q�r'9���ٗh�]�t2�ݦ�4f���L�ސUj��Z��B(W������
��)���g�MS�Gޟ.)Ԙ#C��%<)7��K1��2�R�HT%�&''��o�U˔f�d*E����R;�a�� �oh���U�.ƫUk�@
����j��L/��DB�*$=[��� �1�>t>Ve�ǅ)U������=s�5M��x��$�H�|�X^�F.;�i��vx˾�^N}t_9,�_�v���ì|�} �����J����`�C�o����W�<I2Ô�w�|奪���knU�Jb�+�ͪօ���8��2�tW��~�U�����10��	+����2�/"t���Ux�щ,8|/���$��KQ�t� ���7ī�y���X���t��&#��^$�FDR�;�P�8��y�rkxz�V�����he���v��C�[6�J�)�?)��:�Ӱ��6坾�r������0��o޴	6�i���؛I}�P:4�3۱k�;suwu�Y������26u=�r��p-�1�kRj�Y95��"bz`��a9��!���waa�TL!G/���xL����[�n��������s.��O��ɬٳ�\����>p�9�|�����_�� �^ޖg��vBY�W�~Ͷ�������fv��"@m�b���ܹsŊ�_���Z�h�z-<�j��w�����Ƿ���@(B��\���Ι$<�k ���1�2m����vh�&��q���;�P���H�:����W^�bA�7.	#~:6^�Ǔ��mٺ=����sӔ�����>�3(9�Z5y��C�m*7A����R�IGb'��HĒ�a��r̤����Mwttx8�"M�?ٽw�B���Q)s�6ɱ�v-���2t��j]^g}��̸���oÑoy1�NuV8Z�X��Hs
�{W�a�a��,B�C���uئ�I�%n���?�{�pW:�`�B�"` J:':��C�]�
��Fn�D�P�M�6Gcz]b��}�,�:�m��`�2��5Yc�6I5r�޻�s��ܪݗLC��8CĽ�}��&4JNS�vԀ���~v�k�@�\�5�=����lG�Y�Kk�ө^W�FN���/e��H���ņ�j��KHo8:�ID�7#)�f>���u�������ᘗ͸�����'�)ݽ���(G^vmh����HŠ�z���Hbs���Xxxv�!;1�-�����p�r�l9!p\�����P�gNꕲ�q�!�����ن��YfRUB�Z䮌c���Š�X7��q<�^ҫ���7���u���O��C�V� �U�v��Z*�J��S�\���l�N�ר=���M���)UɷG�фRR�Bɴ���b�6���Ȩ	����`���vE�Y����א�T
k߾}nRd�*���|<�W"��$�h�גa�{�|��,�����W^'כI}�|�S��Ky^}F���?6>�Z�,ʻfs���l�˻��qk��[�Oqo�@�O(�ɘpp�1��{ZU�pQKS��ŋ���w�l�tl�p�K���.�`7��w�s�%����?�����X�L�!�xaBO껿&��Z�Y3��**v��'�\|챏>�����������g?���|��+���<���MЎ�i]>���J��ei�>��L�<_�RS��tIc1$���Oe3�9V��7o������|�{ߋG� ��q5L������jni��o;��b��@��w���U+>��\���Ĳ��*n|�ɺ��xY�jm"�[B�TnxH�����������r+2Ve{2Im���}Q5�<DU��ڊ�$0G���Q�V0Wʆrx^��9zR_���}r���9~��799�酒����қ��@�Ns��P���\��e`�6�DT�����"���d�L�٬�P9�f+�0V��m�~��	R�R,������]+̓P�t�v�|�v8�;3��7�f���%o�3�>j@��K�	������fĉmY����x��-�:;A��f����:��3��Я-��N6 �����ZԼ��C}����۟��.�cb�C��M��	T����T�t�y��*uN��E�k?���N��������-�	��4�z�}]����gq�|jo�Z������f��7H�	˯8P��ks-�JHPۙ�%�t�?l�"@�������_�$�d����_w��L�K����"�>n
yl�����_[��cJP���o�^��t:��<:���r���}�G�VՉje�dV���E��G��|�O���SX�b�`U�P(;���)f�a��b���/��=�g��7�$w�4��֓����5������4�����s��ٿ��G����j)HK��D���6M*U<C0�L#`N� K�J!���G��/Q�B��7��3o޼�~y�������kA�#�e0�;ۨ���V-\���?���SO~�|�gO8��j��������).K�A��Y�N�i��N�d����+Ӛ�Z%��Q�2)k��ۆ	�^*�6mX3>>~޹��y��O}�I2���Q�-;J$ų�,o��bs:��w��٧��o��_�*K����$,� d^i|:'՘�T�&�������*Tx�+��A�ӎ��IE�"�5�
��&lH�t��[�o�g�n�n+O?��?���'�P�G��|��l��>���_�ܧ?��O|�O<��ç�q��S+� ���\y�����`y�)�a����0{�9>��$j�����t��vQ3�^�ԝ\�9/ؾ\.��7����G֭{������⦭ۛ�iL0;ڏ5�6}k�l^�d�|�G���,W�Yڇ1�����R��l3_�gt	uQq��`ǄA����o���#P���JVnJ&2B�S�����84<��ż�V�R
�h!g4�T_8�7����I�9��)�Ӄ�p��S��d8���$�����O�sMsٶ`tZ�PX�B�1��6���j��媜�F��lpV#�M��	�˯�
�X$��z�0�L�|�ƀ��A�A6]�K�P�f�j�����J��4_N�ﵫQ�h�9P��&63��ND��,f����_(*C��	�+����-b�������8�<�"'�|����+�ղ�P�#V@ɔ
;�X+B����!���{�֭��LW_7�+B�����C�	��Q�j9��URJJ-�WsP��_%C�ᓡ�
��v�}_W��sTX0D���X��эb�ւJ՞�T�#�{��VK���F%c����5g��a(�ʕ�bV�r��X6ހ�G6�0�����M�y`�z��9�+$8(l�+��{�,7����r"�|y*n$�Ʋ��ZT�<<2�Ƈ�����A�#਱�fS�_ɔ&?��J$�".Yt�T��XSDݥ��X�q��������V�YcN�$�t"B�ѠF$V�5�o2�Q��� f�;z$0����s9[���)j�\��&(l�P�vL�/ԛ��
.����1�C�J��:U��7jNu�0=Į/_ߜ���Q�^}�����f����fR_���V�,At1��eb��H.�,^MH���&|l���x�iz\-�L���a�Uǭ����pF$ex*_���`� ҋ&��/8����M ��$6!�@�s�_y��;wn��.��mo{����o��s,�SN9C=p� ����2rp�vx��q����T�bk�X4%��J�L�z��!�ዛ�z��Ԯ�T.���(���l���mئ��Yg�������׿��������I75���*-5�2��[��K�i&����X���.ĥ�T��Ro�J�>ZĘ�.]r�w^x�y�|�X�F�cc���~6
1q�6jj����o|�o�����?��'?���#�%��$bQ�P6[��6>6�x��6ӵB��"H��P�~Ő��<H�-��b��%G/������΋b���u!'w��V(����������;_zi�� �ɶ�N��
�*NU:�G*�ӧ����y��t��I�Cu�
�j�U��-���H L�thl���?f��{�����w�����F|+5����O���o-J_��/���,ZԕJ5K�	��S�O�j)|�L���,��c<C������|LŤD����QB���l'��N�=�N�ҹ�ȷ:�S\rpF̒�����_/E�I�2b��|�p�qH"J�i�T^��lwB2��*����@��=L�&��B�8F*�R&�I���wrbB4Eܧ��_?88��,n����/�a�g9��P�t?��rY�������1�9A�Vi�^�}��1Eb)���$�d�~B�O�^�x1�u�ip&�3+Z@�X���˱	�/3�I��u-.�=XT�s�=�(X���%xTA�8c2+���"��:�mò�s�����Q: ��TJ1|g�Ǟ����!�@@GgD8����DZ���}ݍ@���01�A���p �[�Pή�>�69�Fy�Z/�C����3�Δ�Q�@��8xD��va`mmm`#��*qC��mS��?2"�B�0�:���a�>�{����Y�]�7���������� �̘$?�Wԧׁ�&���)�_���O|h�������O��a����5���߁���`"�z�L��U��B)ϻ֍�w���Tc&W^�~$��/�ओ`�����^YS�Q�K�6���n�-pn�a'T���G"!�0����}��.��o�����:�d.;tp0�W�2P����r�MHtX�i�l���ݻwp�t�UW]}��s���2-zz84��,5�x��"<�X��1�;��Hm�֭[�e?��ӯ��u�_��k��v�ڗ�.]
Ǝki�2�WTs;'HP�"ɭn����QX9u�[�bQ�!�$2uH��OSuYS[�~��\y�d���PG�Ad�ՊTs���(c	����W���y��%�-z�;�~�_���xk�]	�³1A% J��&��(�\�'vy�l�cQk��U�����7�q�k�>��E����]s�GS��zҕ.�~B�P_��96fvt���E§�8~߾�7�����.\��ɨ�Z�Q�V�J@ձ�a���hUB����'��1�em���|{"Q��Q�5�jD����=�P&���Wzzz~u�]���Y��]����e!�h�Y���c�iok�Z��S?���/}�E���~b�I'-I��###����z�d��H0�.{��h��0�"�0o�E�MU�S!�.Q����� �+Xm��n�L�XJ�1��N�$���E�n
y���*c�K��#��;v��5�(sfu�]Є��R,R��d Bܣ$u7�W�H;���$���Q��'y�jBQ��٤a]����lzr\߱sl|��M�)�
���,jQN�غ�|��$�4�jY���Lkkk4f���GƧ��JK��th�e|��W��̛3��cP� ,Q�M~�N�Q���:r7O�q��s��Uk��T����U�����S�}d�qv�F�5�)SΩ��d��\C-H���-ۡ�̝�`9�L��pr�ӫ31K� �l������'���_��5��u��?^v��<~�vZ�\�J�:T�f57�44F��]=���&G��SS'�8���k�N����c{M�M=�ɖJJ,���|��T-��I��dsd�E���7��n������J���ҁ����il��d��jKg�i�+f^�������(�@�n�rNU"S�~�<�ҹp�X&��l����ʎ8�U�6�'�v$��b��$	8�{f*F(��� !���(ea�{Ѷx�dȺt���/T���H&tc���G)0N0I�����]�00H1�$����,|f=]ʓ��>CCC'�xbKs�EX�L�KɈ��W_}v����y��iɒ%��Xc�_��7oގ�����>�����?���� �iZ0�Z������L�J�T��[���L��w��6n���佗�z��aC�C�[6�)�F\�TKԽ��-q_�H8��Db��B�?q������w�}7���-76�Ӭ��t��jbo��m���Āe����d����!9���?�\y�+W��ZC�� �O�9U����h5����G=<<�z�j���g���?��_��=����������z<g&�	��SХ���ѐ4��F�����$�b��%K_�����VH��6+U��w�@�7RCCBnʱ��PD�>0���uｿ�}���Ύ�h&���f��\���Y��,ca���"!L9�0�i'������65��/����!|^^�y|�ʙ��Dԑ�!�Yn߱��T-m7�����w�7��̓O�������[I`�{g)�Yki*��ɥq�����
�q @H�#�I���<x�c����~Z	ƿ���}���U����q�K������";{��=�ڸqKwg���K�mX�{�r�)7l�??����ݝ����pg-B�#��dƐ�) ��޸n��WR(�*�B�_,`�88/�/��6�&��Ӗ�Uʅ��Q����(N�|$�o*�!����J-�e�~J��̒dM�����3C���O����{�r6�x��R��(�tِl���tP��E8�=��k׼��8��x���l��(f_x�p��3��*`m7�tn�X�*�1ɝ$�ej(���@��?��V*KT\T#�Д)��`�8p�����\F��^��4VְJ�W�ՠ��{uj��.�"gm��R���#�v������nA����Ȩ�@�����,)�!(��+T7%ޭ�t��&��z0���G�S��W���d�;�^��"'�_sS�lݺ4��/|���/ǰ!�J�T����)&8#sp���cIUU�Du��w,��b��]���$��ӥ�D�fWr�$h�l67K�B���O�DT�Qu�ϋ��DE*�xx�Wm���T���
{�K��ugG���{��fR_œ|�O<�������<��g>���;�n��q�U7��ˌ�XZ|to?�{�����Yg��˻��K/��өģ�A�N���9 ��<h���(�����A�����_��.[���w�"i4�r̉��0a��mZ�$��w��˻��
�휷]v�e�O<��l�D˴l�,'�ڛ������yׇ?|�͸n�)��;Z���0�Q$�iqu45���ť���c�^NL�s�~��|��/�'IwZnMH;�߶�F5?]�:��;�vw)T$3��5���x��5����A ٗW����;?����سg��ٽ�nm1����]k��+RW{I��D<E8z�T�d����gu�Q�"��9���	�}�ޝgS��0��R�kSf��q@�c�����'����]5qێmX�h,LzRe��%UȒɺ���V<����@~3e�̑#���vkV?� �x;��TN5BqvrSY�T�h��s�Am�eR�H*�HFLJ^�6����B�Y0��������|�M7=��.(X�IJ���5j&)��A�n>��3]��|l(%�����Bǯ������Kɔ�Ɏ<d�J�]{�����O}����x�Fu���m-�/<:
.�T�w����N����(�L�힛��^~yt��_w�{���wo�گ~����Φ�9�cc�P�(��	A`L�p@d�`�Td��'40�P-[x.�q��T(�C��s���إxIi�?g!alX��5�ߛ�t��M�2
�!���~j}��[��s������5�N4+�	�����%S��XV,�,�hT��V2��m7M�M��t'#��<#�[U��JS�s֬�X,Z1s���OBa՟*�Z~�!B=]ݑJ)R��{�
��	���SY(.����3��g��@��0;;[�>(�BzO�d��h��H�A>2ʗ�,}���O��r\�¶
cO�.~�ZUj�����}Bg[upOͧ�t�z�P,�tT�P��d����F�p����1Ǟ�[�������<j�2b�ReÆ�b|���n ?\�&�M?������*�����Y�U<z�;I��'rh���2�T�M�0����;�:�	
kS+�%=������=��뿸a�+��D�����s�*�J*#�#�AF��R��Z�:�GS�K�e�I�SJɐ�xler��n�8
�3��R�/�/m�W��Y2���q�5O��0��̚5rsݺ�q�����K��������G�i&��H���|��N�<UK�u���©� �+A���6���;�G!#<���D�vl�M�`9rk�����������.Xz�[�ٽg75I/��XB�b�I�[�Š|8��'�j$|���) <�+���g�ټinu�ig���o&���D%���C��:�*��%"ǎP+���6�Z0POO{ �C��lo>f�1��r^�v뿁�&b�7 1����� ��"��z�-���+����ͦx��ARr�f��ڀ��.Ic��\����F����]�v͚5�|�?���z�=ܹ���O刾p(|Ԃ�`ycc����_z饟���{�Y�NA���iZ���Jf�,��Z�r%L�~��r�\nc�[qw� L�����a{i9�=�,9��;��3����4l�,��BKw�^|���Uڵgן�� 6����J&��O�ք\�rg��U!�=Is��c`�cd4
f(�L����Z;}�z{:����E$�=������)�J4�1wv�@�� >��O�~eݣ�>*��>�D5de�B������Ъ:~H �������p�I���UJ"y�_(�d"i(N6�5+U<�������)��b����8c�-ۢ��M����}�E�����}��7��2��?��fU(�j�$u�����)���%`ݪ-G;2mYX�=O<M��~��S�,��%#	]K3I�IM	��Z5����Dc<���^�����n��G?z͇>���Zا
�N���W����_�T���z�R@�����nڴ�씷{�YgŒ�fip��6J�5n �[����7�P�։byج��8lks�m��(ړ���l�H�p_Q�T=h�8�)Q���T�A���l��������uR�A��V�`p�#�6���և��nj�z�V��O�&˩�8��(6�R-
jn�4�:�S��a��#��=�����2	�Q�8�1�Lr.Ld�D�r'����` �ِ�����!|��-J��z�=/�"�u���El��)��L�|���!Y��R���b=�/૽s��}��k׿�z3l�p,L��P?(z�r�2o��#���=���z��_,~�vYW�����b��g_I�u�(�������e�e&��wM^��/��g���dI�����IV�tu&�5B�����S4~"���\���o��H��^�R��!�A��Ny��h˗/�ƉS��7�G�����)S��ˆwq����ѸY����ֆ���=�3{�W�t��fR7���� C�?��S���G/ܵk��ݻc�RV>�U�d�����*-D�\0j���ڂ�j��y��h8r�	��������?�����úJ�E0Duz��b���ig,9�����!Q���rɊ!�bW��E�)6&���?���[o�;kN�JH}�|�����SO����o��fP�$>d3���G��$@=��d"
�e�E���_��_>��Oa��Ν1�������!=�齽7�pL|i�2=��aJsL	��~�>���P����7n���lv�����| ��%�ꡃC�j��[��951��MNB�f'�b+��[�~�����MAQ�J�����{�;5A`�v�ܲ��:�:g�}���}f&&ӭ{���;;:r��/�z҄:�������7�{Ϟ�_��?aA.����\rI�\��.7(����ȶ45Bt��3�`�ܾޏ����6lhO�=��`hR��9z��U�c���%��T<9봓N;� �u+�����Pu�$���;vt��p��i�&���[��'��'F"hE�^|��O.V�]�-�%r��~e��/��Y��������D�4�B�p��� ���s��U�+�q�E_$�3�of��'�x�-��/'�s���N�X�h8��hTAB۶�`4��ݩ:�e<��Td��s%�*���A���R�HC���an۵h�O������7~s�3�� ��!284�*�a�<E�p�*����T `5�O�:��u����ƍ����\p�s�E	��j�ӭ��ohl3��\c�9	G���C�i�-b���?]5�����r���#k�Ռa���P�h�a[)sIY�38�B��E)f	{K��y�K����?�"���Lј�OՆ�v{����Hvt���d3x��D�M��{�'�m���X��s����s`ssc[*��źq`�o���m툲�ݮ�J5��1��+)�3���: s<�ę(A��.峏�/̪aܤ�����sBF�*�"t�G@u�t
jqQ0O~d$m>�^ �i2����ْ��TG�5gj���{�$ÿ��Wf����ի	5��Z�$����b,\H�mR,)��c����v��Z���:�jL��Q*��Rڪջ��5-[�����;~��}�kC#�4n�����`�u[�r녲��tJ�7TAp���'��*K��`��[D�C��cq[W�M�|8���ڡ��}�@��&Z%�Nq4d��j;-馉���C�[{�y�����뮻n��M��.mj�!���:Um䝆��VCN%5;0�Q�Rvu��!�I�5)X����cI'�M�?eP)G-�E�T�Z����:���3ϮƔ��)�Ke�}r�1���3�c�r�g�~��/���z��g _ & �[�z_#��T�C��Y�w���x@__���8QP�`�M����g��q-*���Ff�QC�D��eȃk����N>�DH�g�z��c�����зl�	w���_xᅋ-��>���D���w�757oް���u��3�8�!��@�aK��tQ��]v�e�ů���Y�fS�g��Z]����%�JiϞ=P;��|�;߹��1SNl�4/=kppK�����v>>���L\j���Q�3���:*�oڼi��c���@<��#�������pa�^gG'�� �EgGC���t~����p������;wm�Ǡ.���G�1�ԙn���s)<���E��Y�m����ڵA��XV531�����UO]�bdx���nŦ�}6��<8�59��O8�`(\)�H�b�`lP1��;Hl���N���؃����ԼJ.��)�nF�F����i�z8�S�f�I�n�+/�,�&���@%%��ݺuz�X�s�=��������W��!�����7k.t�B�*J
��u�V��s�/~�|�K��$��ֹ� �2ȳ��Q���i9�v��׆w�W(�}���U��N-c����۶m�����Y_�h	���?�	�Ls�'Ԕlhj�g�P�Sm����/p����s�����ĵ�^��K���o���?�f��9a��C����q�n��}�45���`(�;��SP��n��:��sW�Z���G]��V6;���d��!��)��#��,�L�U�:�	>�~��&,lAcʏ��}�\vSf��,�
��w�I*�T�ǠV��PV<]�˸sg�b�d`h�СC���ʗJ�8x����s_z��Fp�[&8�Y�By!##�8eP��;�����%"	�o����<�׭��G����6J�A��e����Q�]&<���lh�#����%Y�R�c=��s`���\M蠺������K��J�g6g�رc���#!���	�3`�7o���3O/]����8̞o|�3���N]W�I9#�\[����7S3����Cڴq;oJ���*>�[8B�X��ٳ1Z0���`k֬���^�ҭ�x�_���u��e�T_��"�qt$�G��$z5zGW�	/R?�	�Y��"/3���6��t���.����2�{�q��L6�M�B���655I������ǿՉO^W�T釓2ɝ�_��o(�%�\�â<�ht�������裏��o�p��?�������8�%V�(&���t�ɥ��M�0��¡��d��~���k^���{~�1p�Dc�5���Yg��CJ�������įp�Qaj�oΜ�������`p_�ַq�� ð�HFj�BY&�\ ��� _��۲�����5w�iPn�M7}��+��z����VPPpϡ!j{�M7}�K_
���k]��m_��B�9�
�z{_~��o���ǟ��r(,����f��W�8��b��S���/^|�ŸW[[��fF�k���Т��$,�??�s�=�����][�~��C� &|ƪh�I@-� U[��+�裗B�&�)z�MNL:4r�E}C�{R�HЩ�8$ʲ�!)��GX�Y=��,�'Y����vv6oۺn��M�/�ަ��p7I�~q���)v1��������۷D�`�x�79i�(�ˎ��J�\|����&�A��m(�!��$0���Nd'3Y�^vܼ�׽�����=ڶ�����|����`/J�t�z�u��͔�VR��T�fX�Y��v㶖T�g=���o~󛿻�gᲅ� �KӔo� ��錧tHҖ�o�����~�S�R�gn���C�iHZ����s��QE�R	6�	����ڧ��{vl߂�\���@gmLQw�Xc���N.����S&QHcs[GϬ�Xf�]ɖ[~���_��}�Ck^�y�9���#��(K�r`:ˆB��ZP�YU�ȶk ��90�ʺ���.��op�[V}�L��)c�͝;7�nްq��%݆�Ɍ��j���Ǡ��}�;-�4]�t�����_���i�N�=tph�ҮdCW6�5_4�Q�p��0L��1ʣQh� ��_��\�W�r$��X��d@�c�\��:0�k�>�r�qW��41<:�s�h:�kXZ~�:1>�QB��+�{�+�pIS*�Vg�|�A{��D�RV�n۹��EBv��9��5��X��ig�}ݯ���Y?��v�Z�"�J.��H-�K��_��rU��@�}������7*�Gfk�S��ѹ�FE�C��_�ȳ/*5>��յ�j��n��nܸ1Iu�v��_�uv'��,��Qj����T�!���aV5�=�jU]��L͘p]Ӷ�Z�dRmT@W�_�jJ�8�!	���>����3nS�3�p�{;��
i���d2�2wN{�0�Wc��X"����ĺM#�׿���;��q�go\��o�Ɓ�� �,��b�9J;�)��6J,���Y�̋�҃aB�S{�.j�Ѩ�9���J4���$�!��ܲeR *b[[[__/x��� }�ȅ}��y��Jƃ|۷�L���Fh���[�a�}��w�w�s��ǝw&�m�$8d�A�Wͦ�Q��
T,������K�P0���-;����65�����٥�$p��\ޘ�M&Ms��:�S0���_�:��_|q�i}�>�^���JO�����U%)��`���+ȝk�&�T�޹���X����$���R�M�����r�\�X��b��3��h���z��+��O�R@����LFa�UC.[���K�)�u��3���MK@^`��j�x�P9d�2���W��֭Y���v�i89D��D�UڹJw0H�m��ϟ?����;�}�ُ~����B9�~�[�����Քn�;�?%��|뭷B^�y�;w��0 ����ھ���u�Z<��Z��y������%K�̞3<2|ŕW���'����
�E�)�O���O(zɻ���o}�[�-��s��g��((\��8묳��^h<'�|�G>v͚�_�J[(N�O���3�XWg���?k�o6�]�����#��u�}�������{�Y����*v���&%�rђJ�Z ,�s�{kss�;�bA�<����T�L��N�� ��S,�&����"�Ϙ#�>����e+݅�}R �lGGatԘ�L1}H���M.�p0D�(J� �B��2�������E�p��LS�u*{?j��}�2������`v�W��_>��Ko�����(�Y�m�:0ƕ�A�UpS藰f_}��SO;��|Gi�^J�S����$����ܵG���bC�>+W�j�����x����z�[ߊ�?��C�����/���n�G$�DҕqK �	�
����r�/���o��9�1�O:�$I��m4�	�!_,��#������߃�~�>��kq��Q����n�y?�a1q|�y��MLI�Oll��P%�p�sOa�;��C�d�B�,���)#������$U�M� Og�Hˀ*{�|z���V�j�9�IY�F�+k�v�����P|�I�7*tEY�i>O�PPY��u_�cO{zf�>�1�n�	7.Z�h���5Ӡ���]��a�7�b�9�'o�m�ȯ��Z�b�":��	¸�N��b �V(� H��`ɰvؙ��b�tG,)c�.�/�}�vۄ�Qʱ�bî(M�ʱ��Occ���;wn��:�@�U��m��Ar ��pt��i�}��V�Ɯ܏�0%�0w�*Hu;VF�R�D���☸pr�S���[N>�2%v���\�r׮�*�R�c�pF2S��v�P���I�ⵊ�r`���y��ǩ�� �m���,N��4b&b��͝8�\�h�3<<�H��eL�����*���Ѣ��0
�#`�i��� ��}#˗/�ַn �5_ܰzu�Q˰�8aXd
n�!��J��ݚۖ��*Uk��s-�i�����@]K����94@xA8�B}�q�'P�2�<�?Ɔ�fXd�5�s�T��˨�G�^�Q#A�<���ZF\���Ty�K��HM��/>hx�1�l�h�=�od�L��|��,� ��@�R����8/�)�s�ZF�}�?�vk\��8E!�@��V��t�5��q`CW���4ðW������M��=�t0����(�Z�*�(��TuA����pv4Z�
�MDcў�[��/��r��k2�!����* J�ܹ�o����O?}Ϟ=0���ĥ��4�$��M����
�����N�������V����o��;�8PK!��BqR�X:������C����5�d�!6� �P4���ڢ���}�9o�L׬݆�Z��ľY�W�z�^0D�'m�s.����s��iUK�2n��Շ��<}5�d�SCX���:%
?��#������<�mg8��V�k�a�u?%�.Y2w��o� ?=����h$�iƺ��Ҟ�؆�V4��@2�C*`����N��|'�|�G�z��P�ΐ�aHU˅����~��EK���f{��M�6u�$%��"��j��:Z����U�V}����#~�77�� @:�SSe%�8�?�j���l����w�
O,��{�]�}�O�����W��k���=�����`k�}��7�=�ĕ�}�ۋO=���J%+�+�]�øO5��E��z;�>{��.��c����_���_�˽�O\:�pp����:!˿���\{�R)ٯdPI67�d2���Œ8����y�w���:\yͧ�s�>}�]w��6�2U͚�8#�"A��N�8Ij��͟���W]�	���Sj)���׭y	�b��°���]�i��t&74@�k����"������}s���m��NO�N�-�/ߌE)��a�^l���g��54����Kc���I��]٦�A����5�sL'7mb��b,ݼ�Ƿ?��եX��xa��`�����p�2���]�qE��i�^���t:nٙ���p��<*56��m�>��\:�yڊY�j �M$Ꟛ���i�J�t����ĖM{CAc�1�l�*U*�x�ZCWm��$:Ԩ����j~�  ��oRԊi�٦$�E���bB���d�q0���L�5Sins��^ȓlkJW���G�r�	'��J�U�e��\��?�k|����Ykkzd4whxp�tg'�yPuª�;6EOT���XX��.��2	�N���+Z�
�C1M�4);8���1EX6�a�Сɉ�C�QЮ!4u�����*�;�S[�e�)V�גɶ�;ʙ���{�@�ko�3��
4���3�����H��U����rRs�S�H�"���'J����-?TGI�r�%��r�{z���ev��Mf�M/n��R}�I#o��[�u�_.҉�Y�եMNN�-����B
V���M�
&ՠ6&1ݴ7�]��w��Ά�O����������<�u�C����sR��,��9GWP���j�Z$#���B�x��R��Œ��c�fPξ�qM/[v҉o9s��[6�m|<ߔn��r��8��@,
"�W풑
>�!|ݓӒ�왔�%��V׸Ka��CkK������(+��ñyꩧV�^N���ՋgՕ2<	���H/{��;�<	�C�9
�I�Rz��k�:�/�L�<�y�����$]��{�w�Z�U��ꫯ^�f�w�r�^>���i�	2Y$K��r4Qc�7�=�صk����?���~w�]w�}��T����2�R�	���U�X,G"�+ނ����+��A�T��~����uvvvwS`��[n���~62��hl3�.�AC2`��k��1<�	V�
�ppp�S���=��������rT���C��#���ޚ�e:������y�˗/�Ȍ]kG���e�۽G)��ڱ`��E|}����-�{}���?�p{!9C���U�w� �������.sN/,*H߳�>�p��ba/9�Z�9��~�n�/�1�Ba���}��X{�٬Ys����R�+=E@"�:��ˎ�[T�#>�?��h��1| �����d��k|,C%���Ã�����O|Z��p�R���B!��J�I,��E�6o����O/\�𼷿���Ͽ�?��;̖8����>�3g�-�ܲ��K]
(�H�ͩ&1,�f���I�yO��=�a���?���_�ey��'�8���D�jC&��Ȗ�o����{��;.~�/0�t*ݔj��`��!�op[�a�5�ݷ��ߠ�~��/?���c���_�l(�X�dc#��o~�i����Qʺ�G��2�����fBV�MW�U�Zfp�b�!�B�s�6��;w�VW[w0ٸq#Iz �Q�|0��k|bkۜ�Q���ʎ���j��P�w��ʉh'(����z���H���n���A$Rނ�$���1D��� �_�N	�:M<�lddS���
�Q(@�jo��ꫯZ��,7=�{��$�o1���UϷ�Zu�b�r���
w��jC��H�/'���A�8w'�{ǎ��c<��`��#a��J�js����=�$��s���T���g�{r�H1	��`���͵� x|`'�	�d��m�d!�����(L�=��9Vw�:U'��U]������J�U���g�W^�2D��2�A�[��v�ؙ/�/�_ mؕ��7�Y0��v����,]���:tM(����?0l/�0RY ��$c0�d�{��y�j���h��=�R �EM��l����Օ[���U;��p���;�NWՌ�b�*� Č���;��|{a�0�L|[�N�9�&G��%��U� $�ĳ�f�$
^�!kP)�n�vKA��Z!����2��_�`ނa�.x�)g�~��L�+��F�z꩕����]���˓X�M�{10�0;o���W��e���g��O_�W�y��^��k�`#28?�4���J@ɺD	te� [�N��j�,����M7�t�-��b��jj;6B�lp�e�9�r*v6�6Oٻ�y��ד�B��I�?�J�g�/5!sƇL\�<C�(��O	t ��f֌)>x� Ƈ����p6g�`��ɟ�Sg�#O<s����7��ŷ�b���
�*�ǤP�V�IЁH�,�"�%4r��..�c�F6A�����=�20�{��[G7�,� ��XE��,Q�z��K�\���"�UM����E�1ƹ�Z�-g��p6ہ����^�{��{���x:k`�F$՛}z
5E�����b~Q��&��_��0����;��7��uX�'N�n�0\�T=�fXS��v3K4Y�D=!�l�[^Z�E)ѯ���#�]Z\���/���������z���M@y�H8�I
e"�hr`��s�
AA��O.��T�p�#�����TW6~AR���̅Kg�����ݔ_���>m֫[6aq��_��#1#�+����-*�T�}�F~����k�]N�x���go���[�ɐ,�Bd��4�p,�E�FH�8��,�6mٸaDd~A�["�s)��h{����ّN&;N�z������@��5Ls��O��x�e��pU]�A3������������'?�ɑ�4�b$�Ftrjު�#��@_���١�����.�/�{��{?�?^��?������>ϴ�?u�[�O'�M� ۭT�Z�+��93f(A~~�az��wl=,��x��O�[�y��+�G���9V#b��g,�24r�艢��x��7���7����}�{w�D�:'����-��V�ڹe�27���_�]�����~��/�ӟ��|��dS���m߻��o}��፲���.�Sk�L[�p].al}m�
x�pEk��Q��ƅ��
�!ݒ�3\��f��z}�0b�x$��Vs''&Nwf�<�m�"c�����S��P����ڻ.O@��::R��x,�U.����@&	{Et^��$ߩV:�z���n�x.���z�t�?�ݧYz�5�3��jo_�M#�����#�cx9B���*��6�]�3�tqz�RG��d,	u�~S!�C'�U���Y�������\�\�?�c��6�Z�&�6) �@R%�;�7�hӢ�~D���F�R��Z�bp��&���Xrݫ�Wv�=[�z��&����IX`�=v:�!��~�n~����?�n{MVT�a�HW.*ss�|.��ۦ���4�F��M�fG�� z�E��_��"!UN˒��1�+�F+
K==�=}�J�>66��CEմd����m�r������ơ��6|��ع'������m��VY�tQe�O> )kI飧���	7�82�V��>�Q�AT+�Wr�\e~%�*�u����Av�ށ���NML�-Ne2��D h�����M_�����;�S��R��ӏ=�������G�Ϋ���t���K��$��(VWf�ʄ�v�٣�Z�@�������ð�~�����=b����'��|)����2�t �	���1\�֐T-���yKOw/x�ŋc�K%��"��K�H�^o
X�Xʢ���t��	f&��zRxsB!�M��`��<����p��5\��Wࢺȁ�����_��� ��)7��0|u��|�Fv�����h����l�B��v��W��ɿ�����w���L�RP$�R^�c��k�m�"	�.��w��FD۾}{:��5�
����!a`T�GX	b��,Qw���i�m���pl�@}����_����������wf��� �<�맛�ҭ�n��;z+�k�n���������'�xc 	�V���I��$'B�4;^'�X�S�N���P��^������_������;�|�������!pץ�F��V�U���p�C�t�9��P�rr�U�*���`��[�>[=|�a<�w��;�O>sm�ΝXDaH��j��bH7���n��9����/&\k]c���=���'O_|�+^��=?e��F(oE`���D�ss>#L@�kH`�D�T,�'��m��?��ٳgQ��Q5~��H�n.�^�����r�*��gn���J�v�-��ƛ��}���C��J�P��#��x٬����Vz衇ڒ���}����꒢W�
*yz�_]��X̓��3ԏ�;�e`��c{��{�?|��?~�A)0�GG}��Y]
U��jz���/a��%L~Z��z��'���w��Ϳ�k����$�D,��&3aS[�H[ru%s����L�����n�����c?��u��~{��f��J�"�f5���M��T�|��<��E"�Y�J�����2�G��9b��N	���M�*�^:ٖN���["��[^�ad��R�ĂZ	z��� �/Lj�@墾����dzm
Y@���脦S�Ȱ��d�� �v�c�X�ݓ-���`\;�
��'1o�t�F���MU^�T�\,���3m�؎o�s9��!#ҝ�~�����`�Mؒ�����p8B�I�z]t�! �j�r��$z�E ���I=�n�H��JB}� �ȍ���Y�<*rɓ��j*�=a�|���n�JJX&קn Ǐ�g��S)�
\�@��ɕLF��Ԩ��yMN�94���G@�2]��0���Xh���n`�0!x��Dv��zIr�T�W@��(u��i�ϟ����ag��s[OUVv���dCwvv�"7�VD$�`_�yW����',5�p�(j�4j���]u-�a�M�x�� J!�ŝP ������;6�i+(\���b�����-�-4��%�=���{�?����7n�o�|�1B�fT>�v�:om;����#O��vn���'��巟���?����_��ײХ�[����n�*8~ .Z�����zp�K��.LPL�k�2$j�w�ɣ34<@C�Ɛ˭`}� d�	�H?�C�]X^p��o��C�&D��?������ޥ��6�����9����6#�0;�ɥfX~Ξ���X]�f�;66v�����v���O?~���}��_�@b<���5f�	*P��+_�����ծ�~,�zau)��9q����B�V���9��ȶ���m������f�g1Ÿ�Jn5���r�R�F_��_����Ї>��o~������$�&,29q�%=�P���004��ø��O=�7�7�8����7��H�	�TZ���dR�{rr��BI�#̯Ba�k���f,�.Ze��3єz���ſ�����ƛ�z�K_���{:r�k%�ɚi���ή.E����ȉ*R⩣1$7U�۔��H�x�j���w����r��7�pp7>_X��W)��Q#����*18�;X)�v����$����~�Ў��7����������7ݶ{�n�<ҵ��x��e<�t}϶�w G��	��.�)����g�6�l��3��Ppd|��"����zQ��Lò�a��K�jn����1<{���
Պ�e�m;��>|�wn��_��?��׼�M�b$�d"��8�Z$��M0��L�FgW�󙙅�r�?Ӗ[ͯ�EbK�ؖ�[$���V�/��QX��^y�"�}���~�[�=�XIJl߽�"Q�
��3�8)�(�V4kr�^��T��0��Wg���z0�}��y�����o���]�� $Oԙ�E��dX�u��j����������o����$M��KH���
%�5t�,�++��T��馛��W-&����%�t�]B�S�BoH��N��2���7`b�v�ё�w��c'����������^�Lu`E���B�R����r�h~ C�u�S�������(a��.T@{��=�\1	w�ض�w��&O��T���`���ɍ��J�2��1�y�)�`V�t��X ٥r��Ի:;u=~���������p_�Xmnyձ����t�w�w��������!:���~�N�d��8�:d| М�J	S7"�xL���.�\c�'�����Q�,��S؏��L�O�
����R	��q�U�I�Ȩ��0;11�h�ՙ�l�Jݢj������^W�C�j�%�y���)(
)�\)�����|,S]�7mw
�5�������#]�Gɏro��YZ�_:[�"g{�Ҝ�,��PP*����2���:v�O��+_��}7��d-�ڳ�R*�*�Ƒ���\��..�[�n�.������tvkP�n�x��y�Ӫ��:��]�U�,��TꍘJ��Z�J�X,�����/��ٽg�@O�0�2�UE����RY]>68pk�]������?��_���?�я���2{y��/VX��!�,i�����I�HۺΞ=29�������������~����;|�pn��ث�	�ҳ��"Œn���������)�IO��N��ON/B�ݼeg�V ��
�j�Ԡ��t�ЭF�Kf||�J��V/A�B�hYV�JIN���ޒ�,�q���x�GΜ>KI���w�qG�Zb��>g���n��jk;{�$ԨD��QJ�I�	�TqC��b�j:�R�B{�����W�O��뮻��F�S��ݭ��h�ǘV�HG�)�u桇~ł�jfp�d��2b���2	��T�}����]��n���c`c�Fa~�3ա�bQM�F��F�܃�C�}G������#�Ȟ�۹j��;V�8�$�u6��n��������w��_��W��Ȯ]�DНrb	�\t3�4r=%c(rG�$�TW�t��Z��)� #�_w a��{�����~������{z��q���	�-���1�[,%3��f�:M+�
���tbtt�=�<~�����70�R�oqZ�O�Z2#V��u����	�ccp:�DA8
��O)T��O=�Թs�\w$6�C(�\3�9d�x�a4�>U��v�֭[a�>��cB"<�J�$ꎈ�d��%��% �)�����C<���=�a2:)Jޗ������\��y�(� "��s����JvES��#0��+���l&c{���������
o��_�z�hWX0U��J����	(�y�79��j�L��J&)�
�s8�s'��ӟ��#�<�[������/�
�u�H�X��)� �������%L$F�J�	`iB�f�;�& &�L8@�t�7�}=2x���Sե�JҡQmE�y�
2�x�Gہ����=[0?0��փ�m�v|�P#��-���:�H���3.R|�p�Q&?y��!���M�1|��^EEm��z�ҥS��:"u��n�T���'��'0���1pgݡmڴ�jf��qG���P/�>7��|ףuL`����C"��3�㘓��8��7V�c��H(.��=D{���w"�����gR*tۦ��>W�gQ�8#�b�(J]p!Li�\�%c�ޞ�Ryu�Xu��y�/����ɤa�\�x�v�J��R������:���j��q(��ё��cc'N��+eL�Y�\0�$V-�;�J�V��^][lˬT&�iJ�T�	L&�2��)A3.�_��:�{|/��&�#E�^\�����5�Url�Bo��_}⚕�4k�SK++s3+X-��1{�Q��,�5����,�n�e�ȳG([la!!'pwQQ�
�yK(�����>�{���w��-������*�pu5ǡt�-W["���v�ԩԦ�mo{���G?z����J�������)�-���w�	�qfzr>W`f�n��F$����g��CF[.��	&L-�!1'gf9��䦢2:��~Ի��	��0��/_:Ӛ-��4ZΒ;vaהK����7��i~���,���c���o���;@��Qm{��333�=
�ԓI�Ϟ>ӨԂx����83W�,5E��Cj4N˞v��|6?�gזC��x�kg�}�\w��O����>����w]�֋c���j����b�"�����}��󣾼2��(��Qm����{7�"���_�rl����g��t���a׮��9�+�	�N����6������;w���������iq�%������ª�[==���>��[���7�a��I��x�b�2�Z�������lO6b�c��ƥY(��V���tOR-׫C�+�ɝ�{ш�*Zy�֝�k}�_��|���~��DVԞ�Dae��l�ǭUɾ��	Uޓju�nV�vn�����Z�@�3k����G�7-Gu!�ˍH���}��s��SU���F�Q�U^�SM�{�QZ��k�@�\TSv�d��/��©����n��ae��,װN�>Hjr��OR�\!��=m�z�;sdzfg�lH�kU�]��)��/r0]��14љV]�aQ�i|�6�`9�Q����r��C�U�v&ɝs����w��5�}�k�����h8R�\�u
�j>OvI'Mvu��"zd���ĸ�[��<�dxtxhp�X(|�3���}nSOW���h�l+�z�u��E�ݫx	T���B�Н�|�Ũ�a�2�^L��n��T���D2�=���g�������7��w���T�7�T$��oa~��-m���u�l�����-��t�ı�Аm"�F���)Q���ss���;�6n
�����_@��-��կn4�5��aIuԄ"�V]J�! �h�Ү�=�նPL ���a!���0���زu���7�o�;�Vk���P�lw�s`,,�=)����m��;13�-��2Mu�����Jh�wmc�`ﲺ�{�CoŦ��م�l�����8�~�7ʴ�����|�'�n=f4\�s�
�Z�qe]D�JW{�q�bqa�Ң �܄�ec��ŋӢ����VV"�.�o��ǎ�!�00@�$l���܆�}�(�8��� �v]Ҫ�mT]� �i�,�R+�v��Ut�0���7�2�.�^%�w&��D�z3��RI�fz��b���H&^Z,�/�M�%�5'ӑ]*̶���B;;�_\JBf�����FȨ7�^QUB`*R�����gσ��pG�s��4���ɮ�p"=#�+�guw`�� pCap�,�>Y�!��I#�W�b�ذW|��,�4������W_�?��d���=��e�!-E�Í���eW��\wq�,�=�.���d����lz �@�/�5*���چ�]��qū�0ֈ��P/h;�����[;:A�3��c���$�?�\�Y+�S�fWGG�R�U����~;��w�{�׿��?��׼�5��o��r��!:�q8�WNy�T$hd�{ꥋ��٩��v�����~���3���8�̩h��B���׽��ߋ�+�n�\Y��zP��55fDҊl���
�}h{f�h�[��T�@ ��@e>�� ���a�3��s�t)PYTt�.����O����y��=���0��I_	��s���ԗ��-�V�%�]��8�j��zyV>f�n�ࠤ`|x�>�D�����UZ���n������;�+UY"���8��P6�H@垶Nñ�/�ŹM!(������I5��7���2�'��Ha깿�0b=�	�i|j�o��o_�K�xͫ_#QR1�"<����Ξ:
s���gY1
�`e[�L��D��lbM-���v��8K�������z\ԧP�&�F�"TP�hVxV������?��{��72٬��=�pll���b��K�\O��L�{�b?�7A�H��Z<$^�4<H.�`0��ȅ:r����t���T�4A�͊R\�k_�ځ�_�_R�C{8ݲ3�pԥK�xơ��O=u�������r�\O侉JB�7�]Sw�j��;�*m��.��N$����,��ѫ���J�8��?��~���~�~�͝]�7x�W.爴R�@�0�V����J,=��J�q�!Q ��/~����g��J�@�#�f������iY��RBm/�0����\���A�{�\\؀�����|��sw�u�m���� �K�me�ڱ��j�a/,����E/QǼ����/�y��%/�}��|�+]��]��^Z+
r~!b��5��R�t�]qΜ85���HEi�%�d<�ٳrf����*H.��?���6ʅ�4j,�GGQ�-���"�d���.}�[�D�7տH��(/�T�~���	�9L^����d9�j��0��\.�,�sM���`!@Q����n�:���zmٲŴ�D1�*��|[X�����oP��������`	��7�	c�xs(BŹt4�Y�0v�r2RQ��Az���œj���cP�Ν�a�.�|(��HsZk�x����p������$j���3�����������RJ���I������T���r����-��.\�D�gYB���2m�0A�UԽ�K������ 62Bh�S3ǨZr�q�$�z���Q�;wNNN~�#y��~㵿�◾�-�Y+���� n�94�`�L[r߾}%�x��ɑ��;�����|��_����̝w�9�a�D&���Ą⑓́X����36e*F�`<]�'$�|���8M��XG�R풄��g��qd�������9s&���_�����=�:���O?]Ģ�k4��С
��Ņ����ё-S���*L�fN�ͯK���ve�o�o49�m_�p�M����aP&A#	��w����m���A"i��Q������_:!�<��F3"�v	kf���Rww[<*X�ղ�Nd@�B#JFS��H��;ںQ\-K)r�+�Z)R����`<�v�m�x�-�A�46v�s��AX�eG7����b���p��z�˵�hX������v���V�]�!�"�����aK7LǪ��8��f����@_eb;~�������쉏}�c]��F�\11��݀��N'��fWWs���}��G�������k���)A�&�O6¤�bV[R��^���E��^����O���Ӻ���U7o�x�¥3�w�ޱ���Ӡ	�P(�2�詓'w������_~����.���D1E�&�/!��<��+릞K>��Jiu9���K�]F�l�DGѸ�5&V�'�؝�H�JOW�7o�����|�џ��]�z�ͷ��j��QJq���v�aAԺ]�ًc�._�馛FF�B�����O|⡇O&��>�JYW4Kd��kX���`=C�SJϵa�ۚȕ����U�d��"�����԰	d�\����ށD{j!����~���'ƹo����Fvl��(opx����C7P&C���"���3CS��_z��d�<���'�9I�{
a�tw�ޙACS]Y�r�Kjx]/�+-�֤�z��Ÿr��5hf�p$�c�n� O��'�����U,�rH���l+Acd�z�F6��T�rH'T��"�R<_/�����6�2�8��b��J�ֱ�zu���]h��FS�u�WEwE4zw%���bP��e�\*WM��vt���ח�ՙ���3F�H����4-$�u�<ҞGZ���d��'/f���qG�>�i.����0K��O8ԭ^?��2����A������ިK�m:�r��n��oV���۝��>^3�;��Cg���YYY{�T7m̌Yk�C!Y���8EE���K���W���F����˗I�Q[�����
y]Q\Y��D59.:)�*lt)�ğŬW{����c�/���{~��_����|����M)C�ΌB�NMS1��4B�G�S�@gx������'GFA�s�y��v�b�C�z�Oy����k�(�G�j�k�x��_h��h �z�}pK����p��J���/:<&{"Qw)���{~���;����׼n׎��ha�r��3�J_!�UWn�ᆙ�ׂT�>E�(���?��/�$���%2�h�?hcP#�,xpn�Ơ�xC _B���q�@9 �/a��`H.��\0�>�]~.V�z��y�GѨ=�n>��������Htfu��Sê�t<!��J��^pIl]���IQ�ތ��D�'���[��|PFe��3�J�j33Q�"�BiP��H�e�Z~�߈�#G����z��8X�b /�3N�%l*�
x6��~�.(�h�F˃I?��A����	�7{(�8�����XZ�"FD&�ܐ.��K��a'�4R׎�"���I�������S�P�,t!�D{t�h�&A#}`19T��~b0����/�����2?������O?�λ�����3π���3~"-�@#f H�Oˬ_/��}$[����0�uGK���؟�l�N��O�r��U(�SӋ�N�������ï��W1򭣣�DK.��(��J�u\��Y�j�fs�|b�.��cq��U�ɶ�:=� :�Jۋ�)�sjB�g;������?N�k��{��E/zVdyi�7�������<̚t&s��������߆�����QE��qM��4U���}��W��T��u��/��f�a홚jZ�Nwt��f²>��c����������K=1��"�5&s�|{����c�p�������������9ޡ"#A����8I�Fmn|i]���ZGyu%	�2s0M�Ye4��
y~|~�r�k+L��Uʳ+U)��H`6�h�j
x�cC�>~,e���D��?���`a�$l��Au��"�_��Z��"�O�Z�z�8��<D�E��:�G(�>f#�J���R�
�!�`���%ĝVV��L���5���{��B.�)kǅP-ץ���	�ӺT5`�������'	��C:�/�M���f h5bh�6�)J;3��g�1�x"�y����D,�\�|�n�k�̣]�~�e�s"3E���a�W�"�PS���������o���L/�%����ؖ�4]ʕ�-m���^�2�&���߼w?.�[,b��*�T��a�O�w{�.^��EN$'�d�	Z�F-K��t7IZ3�T�=F�S�|�Ա�/~��s��{�F�z�yX�d������|~)��L�N@Y-p�cj��.��� T�n����;w�6�#�a@�p�6Fc7*�9yb�3��_ؼ߹X�!��_ب��(c�8�H ����W�H��$2��,:]����Yl��q�hndd���X�Ph9��lr���d5�x.�LK<x��GЪW�+t�&��E�Vˮ3=:8�����.Q�k�U�U#w�67�P�#!-�Jdے�dT�<��Q�*�kKП�4%$��ꇄƃp���b	D?+��B� ��sʏ��l�͑���[�<� ~4i�&<�^(S鸶���dM��Q�g`ӿ� �6��ա�;ш���F8���_�*��<
��{������j��)���A�U؍���8;ՈƏ}�\)&ɚIZK{Z��y���m�G)_>p�m۲�0��`Q�`�������N��\}&��dy�
R�|�k2߀g@�����T?P�Z7"
�n�Y`���t1��[+��gϞ�Q�m�Fũ����Dp��+Ҧ�DInb��$�O:��*#J�X(	���QÏ���i��ҿHX�}� $���Ņ��̤Ӱ1'/>L����TK+�{�|�[��)��������X��9;=�{��XD��w����U�m��7�F�IP�� D�\RBb���!=S
�&&#���S�A)g�0a=�4��+IM����v����y�p����s���~��}����/{�+�x�<j�C'O������b�RJ�]s�����=� ������-!X�v���Гz}��yġ�Pԣ^s>��$������쏾�	Oo
zCr-D�5�[S%[�n5�;_YyFT�SW�Ź�-[��c���y��07�ў]΍/��_v�h__6]y����?�3w�fS�IEOx�g{VI��R:�9����w��֕�
\A������'z�i�d�P&p@]���4������J��{C2J��G�z���rr|���l[����(�����<w��Iׯ`�����T�z�S�)��O�vUI#[�9UK<m~k�֎��jRKڅ��UE"�Jk0vgf�$���r��caidpx� �$����81�ʹA$�Xwp�s|�L,�o�֝�wt�%�0;s��C��+&("�gR�^lv�Z�1E�T?�h������|R�R|hz�P�߳;5;[jX�W��!��������o������>�rs���O��MB^:u��ΰ���������H�g�=�uk��/#����x��$�vO��I�ڌ�)��NhW�m���p�f�;{Qc������<՗�Ѯ��T���x���}'��/y�K^���{�����b�:п�kbi�JD1Z]ۖ�N�%���rB
|��Z��<�������=@=�D@uwSA��7��UjY��h�q��9h��c=�L>�l9��\N�9�hxK6�~�#���V������������"�3�9Elet��88	 �t�֭u���NKrp ��A�_�(�IȹĐs�`�r� ���D����0������-�n�\�"q�x��V;d�������c1��U��i�aw4>g�DH}�rK��$�AEk��'Dbb�r����H�5��bM�F�S�[�^�bn9 D~a�Ѥ�
C�c9���K�m�h��5E���JP��p]�Sb�w�&0�t����( onf
�$WW�J�3D8�ї[z=���P�+Q�+N�V����VrC���(bP�Q i ��<���E���$��^t��
`���S�{Od�˄��	"��hI}
!Q��|?�Iy$����;սh1*��M�GKz�
=,F�pב����G�1��t2��1�����	�K&ϝ>�	��pg
j�s�_��?|��߽��1ϡ�*
p�(C#�:䯓հ�~��$S�'�z���d���>,��B-��O؟6��J�0H���{��,�U�M����������������ki���]�v��.]�d��o��G�W�ۆ1�j�L�c��4�#x>�	�IV���>����[��z$�@��8��82�"0
?_�pj����f�h3&S��L;�=a��U�ʦ�˦a*B�
Nc6��Aܧ��jX��@��y|Lz+k�1U0@W<,>Մ;�M�3�Xtx��)l����7�ppn>��U�x������>J�
wy�F%'��E6�}�Wrzx����!�(18h�P�Z��<�?�"G�2)��U溜��O�P�j*�b$�"�6`�j�U*�e��"�St�g�=X�Fp'�`��y%�Z��kX��19RR�,����.���o��2�gN$b}���{p�s��E���Y�2<������+��%9WX]Z^>��g�Q���e�N� XP�d�-���K-�ϬL���nQU�LH�3��#GpǇ���ַ����7f2[�����[.I�ѡ�R��6o�|�ܹ@!�L0��8���U���@H���� /���uF�����L��!�-8!޳�g1��]�<�LB.l'��"��0�	\�����>�o��~���G�`o9��aL��H�"�hwwo4�(Wk`��TZV���	<�𦑕Յr�Y4�P����{_[������iWo�����"f�Z+�~��{��qR�Vs+F8�N�`7,�j���#���J�Z
|�
������8�o�]��K����Y��f�l5*��?w
\�:777>>��r�E�`���I�ݮ�8���ԗ��5���g��O�F����IBY�)�$	�iᔲp1���)�
^�G��bѰp�z�r]`����j�$Z�S�Q��9��*0�<��ǢQ#��k����+@���Q)���1N��ӝ]g��:Ғ�l�ϿwU���4��<�����>r.}[)� K�@�T
Ţ�L��;!�I�����zq�cc�B�Z)-�����jly��\)C3�Uy�";u��w��Ba]�x�'}n�C����s��7C�G��L�Pq��Mt����8q��������QCc"i�5jD��M�g���/�r:-*���_�b(at��l��Z�c=O[�S��h�װ���Y��{2�)�XU�[*c�� �-�
U��>����=���(�����8:OD�!}���z�j�޽�U���j�f��x�#�/a��=[!B���P�@DZ�����)L��h�ާ,8�ݓ��MbO Z�:����Z�T����v����N�|d�V��'U(����jLՕz�j�n:���#2?�D*�B��D�P��5�8ٮt�"�5�y�]�����A<k�l��`.��dRA	�Q��O�x���qS��Y�Z	���������Y\<?80�J�EJ��r�[Y�n�w]G2����A$
��n��(aAӯ�Gͤu�l��}r��r;��Z�qr�v�J���'%ɚ��NBC�`�<%nZ�>���P�7�~�+�o��vE�T��nu>��^�ֲ,���VRa�K��I삍���T%f�r��r�ʔuB߅��{�^Z.�R��4>�ؼ�m��ݥb~`ح���XێTeq>7y9�{C:9���J����۱�V���ՙqsf���^�3���,?Q.���thH�[�%�"s9��V�
�NZdߓ|XH^	4Z��.A	d�a�B�W��]�9�F�.A�����s�?����=����eߦ�m��Ǟ^ΕsU����8,���l>y~���/6����f�P~��R^�i�oP��A�&�qݵh4�ؖ�_U���0�d���/��u�k砀"���K��Cٔ����C=�����}�|�������<_�V¡0�-	���G�eq��'u�4�N?���Q$�zG��ص��Vk�i�E.	G�D�.etcք�D]��KK�rb�	*����V������Ir&����@㖻�_��QԄO�E/G[	�wesM����R�Pg1�l�jnצ[��)����Lk9�������-�~�+� ���&:B6/�
��+B
�����.�Ʉ�L��A7C#c�q����>b�=?��çO��KT����w��C�7,A|�����-��U> ^5��7�U+r��nK�X�r
w�c�
=�0;�������p#& =|���������HXK!I,�>�`	U��GrXhH1ʚId�r�;�2���#:�~�d0��Ou�g�ج|�!vHC�6A�T��	X�#�[6�V�ĿI���:���䕘����]>�ߪGPC	2�\OT�k��$�׫�����2M��
E'�5'�j�[�H}lRۡٸx�"����=��#�H�UwMqw��)��/
��?D��Tc��1�?�g�0襐�:�b�j�����$S����6mڄ���FX��Ry�B��g�K��˗�e�8�)�!�eO��P�!�D:�U����>&���fb
dQ�L����(9K۸�]U��M�U��D|���u��K�	����z�"�1�#���T��-U���B4��kH�iu��o�S^	U�0���X���&n��������_�H0|��ZH��Gm����E�^���KV����bF��k4��D�{6��c?^+aB~�¯1F� �v����.�Jd;��9ѳn�����BW�0�����F8���_���gNc���ӄ��J���'���X�I2K5Z��`b�r�5�@drJk~��b!ڳ&�����g� ��PH9y��>��׾�Eo~�n>t��G�勅���g�yF�6�}��A��#��/��pN?5�=s+�yrr�ҥK���"�W��.@V����`��-�-7IanI��t´U��뮻tq��D��k/����vi͟�q�Ύ�z�Ny�zC',!�樍[�cO<�Q:|�M���\�A�y.l^�a�q������*ήCl�L��Ju�!� �2�uz(�	��pc�,ThBT_��,P�������"w����d"]��1�l�M��z��K�34���z&D��T��!���d(���`;�T:�6�r��N�)�2un3�8丘x�V�J��u��J�R� u��8��獊'e�$q%D��__�a(�LT��]��u�Ų��������V�Z��"��:�/���aKQX6�\Lj"���'&�A�i|�V����������dCh*�H�@"�p|P��`��,��$��=iL�B-��4@ډ��^�!hGE#����<QPG�m��j�{��@Mn�N=Dբ+H&�6;R�SPF�f}Y�=!酪�ED2,�̺槒�XT��Dö؃E2� �5L�����P���W
=p����eQ���5�ȉT��io�h����I���NDQ}A �f5��mO8ujB��x�ʩy�U��2e��x��J�/0B�|�2��r"�u��f�!}²��+"�՛�笛&vx`ȳ3So�8$��t��=ힷc$�A����j��Dm�L�@��k��[]�vw�3��FC���]V�PclY&E�Hd�S�QVEu���}����:�n���#�[�=��á��d�A��#��k5�b�::�˹)��o�D%����R,,u�(�_�D3��\KR�h�I�Tgv2۶�!��rE�n�,�йIbRv���c�bL>S�ۗ]���)���tjD-(W"�D�����T�h T&/O`\�<��=J����WPT��Fi�W��3����&BoϷ���Ȯ�VV�R�#YB��
����ɛ���?�<�Ŀ�?��o}�[����z�����#G�o�a���X*��SK
������2\�k�ۦ�����ϻ�@I�\����9�k�@ꪦS\��>qi	K�{ϾŅ�b�����G�r��j��;5���T�����n�={���P��;;3?q��c��:>t��e�Т�riyY�49Oep �A�3)�<�Ƶ���`3j���a�����x�p�"AN����N�V�l(l�j�ƪ{z&�Q�Q��ۅ����������m�����Wڳ�'z�{���4��ڠ�n��y~������� c�C�q�t6���)#�+�-[�pX:68��q~�S����&(;Sm���-�8_�}	-m���k��-��&]K=a��қ8&���y�	s� b�b��=x�M�94�Cg��U�w���:� Zi��%�p5��Ň�Q�0B� \�RA@=(LI@@8y���
 s�w=��M�Fp#�Nit���UU�ۊιt�|�eIx#xZ8�����5���r���f�S[k��N!]w�f'������q#:����U��s�����0�.4�(*�^�(TD�ݚA����)wϪ3z���zMS�N�H,�Z&>�Ξ==���B�k>����ij�w<����d����z����e2��l���G:k�"�(fh���4�[�i�xji�M�C�Zi
rH�cT�+�[[^	L(k�-Be�Zx0��ҬPC-(����4$��
���f�U��)@�C.�B�zT�I.�|`���Wt��k91�T!����'��چ�w���q�ǃ�U��[����$��iXH�,XY���rP��	�W��e�3�"Vm��=�k�A��� pH�+�v풴0��')�_j���W�&lZ��bJ)�Cw���5CH}&N�*���婸2��2���	�`�ė-����zu�����J3���7�d3B�dJ&ooo8�W��U'������.��O

bmm_	����3�\bO��=�0�}��7s#W ��i���X�cmS?�i�F�iH�x���<���=��`]�2���:i3�@��L�e��E}����STD2/h�x"s���vU�
%?�h�2���0�x���'���i��hc��4J���-�<8�eH�Q*����͛O�:��,mݺ?d�7N����V��"h�U�\�ǉh-��U|bN��}���dZ��e/��N�����ϣ������>$�L��!#By¶��m�d/P��~�j���vv��ǌ����C2�JM�QM�ܒ��̏c�-��J>s[n2�����X��\�~�j��a��'>�Z(���QǕ
�ja��j�	z�qe�~�;�RoP:��o�%Mw�X��j$3�:)"U��ժ!��R `�XEQa�m��G��Q�����소��AS��(C�!
@Iͼ��mFuV��D4G�TA�D��
.N`r)L�&���V��QlOd��
�mCl�T�f�#n6۱6�"qؗa[�d����]�4�Uʾ�늦X�E)r��i�_-�k�b��#,�]"�!z��PR(��d�m!H��!f�V$[r-��EB����&u5���W<�w`��=�f]I��UvG�5�T��U�߈�  ��IDATQ�j5UU��N�ᐡC���Bx�U�߅�,�+"�Ac��h�\q5U��	9�|)�p���P(B����XP<� �q�Q/V�a�/l�������J!�@k�&�wÊ��/���|�ر�
�b�b���6|�#Q#z������Iѳ��T��D�p@ǆH���B{��V�nޘ-l��&�-��T"N��SIS�(�\+5b	������Z�a�^��Z�TL#%e4�����ѐ�.��{[�Q�L5������(ߎV���i���������?�e}����=M�Lp�'ރ�k:V�*-��nJJ�^@�g_!� V��?�c&�����Ӎu��rk�l1�[��ӭ�R2�=�Iwe�Jh¥����� ��3�ʎ-Qȼ�ڞ�k������r�y�r���Z���yJ����"E�q��G�<;eD�������P4{{:�ѐTi{�e��jB���r�u?.b���m��$���(��u�!�tl�D:�(�����i�b!�5IZ���\K�I�LZ�u��Qll>]�S��Z ;���=��&\h9W�J������b��di�{���xN��	��y4N̋KPv]�k�}{φ��eSb�)\�l>�LP"�-τ*�'��O@
Ԩ�S"�x�O�;6fӱ���>��gO�߹c�����G.Z��_Ŝ�a]KĢ��Gca-�����W�B�OOO�unn�T_m��ZN����9{t����)��s����`j=}�����4;5����]h'C��[�����-M�M�5�C� U R��TL���:t����D�5kl,�)S���<W=	���)�3�;MX=.w+"��B��b�@��h�Kˋ� z{{GŁ��Tl�3��l�0Z�2��"��I�K����
'9�,:���͉f~+S���c��M�S(�ܭ��Pe]�~+�� $�H3PH�0[�\�NI�1�ժ��P�H��F����Y`��h8�Ym$�#�ba+"�TS�9��i�Tg[�D1ݖ�u)N�fÑ!���㤈\ByM�K"f�T��(�+	���cP\E�-W����l���	�Z]-�s8�������ֿr�O!���"&�ԗD�Gy=�����G���� ��eQԪkM/wX�ِ@P�@�Gu���WW)����x>�ܻoΫ9�j�D��0�q	0+���:e��-��a���ԉ�����<T�ugEM�)aK$��$�-��aq�'�J��}}�l���!B������z1�c��4��Z�����-���6�x`tu�TZqn<Z+�f��4�XH�?�.��W��Al��s��q��W�>���k�)4����Em�����*h^W�(JF�W��R������,�j��M+���0�M���NX��K��|Q�Æi�J��<sfUTR�n?#�
�~�W����D�OO������f~(���d/�J`�qEn4U�՞ �
d���y����`���ҿ��#�\�k�y�6A^CXi�,�� �l6���
!�N���^ۤ�Z���a��Tn����K�FFF._��x�344��08����gl^lvHON�k%6��Q�w����@��'�CCozӛ�Ƅ����u������.����!gƊ�����5NbT^��5�0���*$+l/>�vJ<NŁ���h�Y䰼��;��g�nC��7�l�|��%�r������ף�2��>�fƦ�YSn` `}5Ξ��!J*���q�b����g��,0�G��%a?i��Q��4���E��9!��/,Qe U�'�h*��*:b���uS ��L[�Zh��!�����A��a)_l�L���ؕ!1zr��,>�3{^���,�Y��q����+*ߨ�'����2�	� �kوk~u:�~]n����L�c�a�(BƓ�";��V>V����(�a��<��At�HQ�(�i�m�jGB�ݠR��i	_b�_�W��`*��tU�""-A~1 :�K��
9�d��65U��������XeKd��Be�-E)�m,~,�4Y�@9�l��L��L�B��q\�$�N���I��@�y6V+�a�S"�BO+�Z��˫�FE��]� N�x��^�9lC�6���CZwdRB���z�f�ڠ����}��z҅�F\�\�|᝕I%�m٬9Dc�A�եBg�3�8���df���
)��-���� J&{y%��f�^��W��m��0�|D|n�7��R���a�H��\�������v)нz-M'R^)�ؓ�o��d?�r}��p,F'EDӱB~����W��18�[2'�+����y��.��~��L ؂��ca�
5�B�Ԡ���yv|N+^ �����91�����辯�E�=ЛOM2�#V!I!�e�8�2'�M�����������5J��M��K�rA��(c�r��Wp7a6@6�"S��e�峚o�Nq�|���\���m�\2m/_ɛ��(vÕ:�R��V�����dW
�]� :�2ż5��6���1m���M�b�u��r 	�e��buźʞ*���u������TFE��Z���*�9�T���C��m�P�-ۯ�6^#�\�UC�zT8(!�-�rM�Brת��<G�p}E)�`򓓓{��9�|�@��>���}�v�����`�����4��[��B�ef�|��(O-��b�b����g�}v����;u���_/�y�Һ0�ZPP��1�1Nt�c���)�,�;����&��X��v- 6�y{�"�K}�"����l6J��7n<v��'Nh��Ъ쒩�E3D���ܗ�:�&ɰ�f7b���TP^�'tA�����Z¦d0X-�㻢��Y�����a݅�Z�_�TZ��V�<?>)�RՎ�����c�RC/��9��l:G��7e��+l,��aH� �\	|����f�}�&��H;$eY�j^S)B

	_:�oG���+_�� �!��'L�D�Ӌy��+�*ɫR~M����g� wY4`Ѕ�D�VE�EL����h,��jm'I�-IkQ]���]*Fk���N�׌{�I�"~�s�IJi)|5�U��>:U������h^b#��e��Bԁ�H
ϓ�ƶB��CL�7�m��>%���dU�&Iv�Ʋ�oi���Rm�l��ϤJ�j�3��KL?�5�RKE�
}N�k$!����~�
�����SIE�<DW���x�$��3O��o�uD�(Y�J�Aq�U�����I���uk�x��Ц�����X?Ζ���0�V����5����G�����-
l�����P��}��oU������Q�h_o�����j���z�[�}��J���Yk*\gT��K��R%�̆]��(��-uv�ccc��q��[|�\����>*�d��XHk�.����z#�S�Q�nDɊ���qofIYݍ�~�{{g�af�D@p��[��B%E�h41Q?5QQ㖸E1&���D�5,��:������������s��[������4���V����=���ˆZTU$[9\x���Kgb�܂�X&k�;V���>!.A��
���A�&M:��{����^c
���G�4����:�,�`t�W�ӥq.�NY�|��_%� FC1���pg�s��%�U��K�����Ә��)҅=�����L�cC�[r�U����$Ӧ��i��(�3J���n��bk�H��R��In�||5�}�\-���\����V��Ŏ�wx��������
-�3o4!�(��L�3Ak� =?]e6����N�Byv"`��h�a�i��s^�T<B�xL�a�$�<l6+��A�<�L`̸pK��u[I&�-�� �\��_$��\�l�DB�5��oPb+��Q�0�B\bA���ti��i�Enu� w4��djb�uy��$�WK�F(-atdR�W\q�x�Q��e!zx��z�tH��Pf~�'�[P��A�vvn���TfF�<����=i$���]�5	jAhb�[)n��B
j;������!�&?�
�'�}��B�~g���9��e/e�0&��O�@�h l�1��NH&�����24R}2�#��L���P ���\�)�*d��]����!�ל���#�:�s��VH��lAӛ�4����)a�����Ws��J;)hE~e�Nl����`�����_��So.(���Z����F0c�W���@s1��4��^���l�Z�ZTe�1d[ܓ"��8���	�����;^�Zi�6������Dձ��Tnvf~��z-HQ�H�������rkT���|�&Ӭ��q��G��Dp�lObU��1�֢�~/W٦���c�G�s�T�Mܒ %H�bO7��-�s���.�<���PP�EI���Ks�Yni\��Kx�~A��.#�5L�Nq�>�z!팂���2z|�����EB���f�2�x��H<HL�D�#� S��TP4�x��ꍚ�
�To��a[�Rb4*�M9�ئ����]053Vi<�v�F�U�B��\ۖ�攤���P;M�ʐC8�ƤC���ż�Ě(��Hsd��J�3L�9�Ϥ�H�k�OO�|���5[����Es������н�j���9!>X鬓�c�2�v|r���|�����N:�%Ў�zd6������=��r"?v(�K�����G��u�]���0����ګ ��o�6���/C1˩8;6<B�a��O��S��Wƫ	�
�i�#��*̝��[�C6D��m	��$-�8�i��]��_5�
�D�$]@"�Ĺ=_��������7�	�.q,S�XQ&D!���"��rO|瓆H�cS\C��ܨ���}�VT�Ք�!���`�{���)�Xc`,>3g��"�_�u�����}�<R���4�i!���蜇rt\�\ʶS�9V�o�Z�LN.UdҤ��Qe���V~خח#釐��N��q��C���'wN��^��'l�E��ֺ���!�)��=���f�pTP~��4E��Q$vZ��[(g����� �B!N����;�y��rh(��,9v�'3i��Ѣ�|��rg�khD(��0e�a3`��m�s?�/B~����"7�}�K�~��XiR)c._��dlK�z
�RV���Q�IQִc���+7��?*_}��ao�ј�mDL��4�;Nꥒ���X�-�OЪ�����6m�D�?1����*���͢x�J%�ueGP��N�m[ļ���TY�@�bLd�n�,�/����	k'�?My�%9�-7>Bn�6��G�����#�V�8�Itv��V�Ze�i�<908�i�u��D�2����h����/�.�(�(ԢY�7ˁIe�otw��Z��L^/R�p/�%�|�q���^=��3IK������}�@%%��Q�H\Ў�KB�ï)��O%,��K����!\]�m.$���c�j=s��!6����q�9gx�Dx;vL��
x��n]�wX�z5N�۷O2 p���ئM��+�JDS���ͳh����^*�C� ,�c>=J����-��<���X9��+���3�r�M�PqBg�t"�s;�e:��7u�Cqu��ngL/�fS��fr+�3�a�2�2a�O��[�P��+Y���W���}n�Z�4��ᑺM��������?��z��u��lQ�2�lO�ӶAy�=�?���W��@D�t=�뒯��� �j5|+S���l�RkBg(4+�)�a*W�9EB��<�5L��Py�lT�NQ|N7�JI�G���?��J�& IԢ=/�=�@H��u��^5tHgS�&8�zK?|lc7(��Z���`|6����i/d�� �6Y=�\��"6�4|���s����L{-�8<�e��R��ٽ.V�� !�������qoŊ�V����N�5 j��r����8�ѻ��l!���<��e��?Y� ��xIR�#�
�efɍ�K�)�#<"�"aY�P����t��7���=?]��cTg��q��Sfʴ�!�|1�i�A�����	�и�$F�냫Vئ>:>>?OIy#���r�+������e��Ml�v��|Y��C�М��y髯 uP��^`f�\g�|c���}����+z�X��K�4Ҕ9�$8Wg��t�tۡ�ʥrQƬ=��6�]�a�uHk�y�ks�D�Ģ/���ޜ:�2����y�3�V=�o�<[��Lޢ�����3�,��U���Y,Q�1��l`U,fV*��e�������q٦�ʀ"֚1Ϣ�[T9-�"�6����VD�U�2@&��{������� �J{�8����-j�Q�PsB���v��N�X��9����|g���_#m�I.���[TIe���ź��J���hL2.3���xt�PZ�h��W�Z��}�	 u�VN�g��hy���&d|�i
�I���dX��* ]�%�|q�9�[CUNz�ON-�"'�-�t�zF���Z�ٛv���p˩,�(�k��T.M���h�M�=�s�'OyEY��ܡ�0�j2�do�G�#��L��t1R۟�����p��[n������g=����X�w8������verj�M��:�m���g�͹J~����$e�t@nڡ��Z~wI3�jE�z�)�l桇��9J�֙��؉BQ��1=����?������DW �8������smi�#hc;�2���m�ޤ�Q� ��
�f�X�dǮ6ق���=<�J>-�k�U%Ő���S`�P�泺�	�;�ȁ���B�i��:`ԏ\Γ����]Fփ��w��C��1M��y"]��].�΢c��!yFy���@��,T����k�o|�����A��VV�R�Dſ�Ń���r�$�4v���L����o����w� �&c�<<��$g�ʥ�+(F��)r�lj�5`�<�h� ��ǭ]�I��6a��H�06%}5�JG�V�@
5E=N��E�����Q��;D(��P��:�>6uC�
�f�
���v�����W�K�r��-+�	__[�S���  ���B[�e+I?j�t$+u�E����^����\�\�bE5Ml�F���(���+l�Ey����������j~G=���0��F;�/��5��3�)�M��ITn���98|�Rǈ6�
�ǽ��C�?���6U�3�	E�
�wmJ<ڰLh?�8i���҈��0�W�m�׏=
�"�?�n3�S9�Yj�+��uЕ�F��aQ5��r�\��QK��$�Ǧ΂[��O�c��<v˓���zAW�l-����%G�E�c$�Ö�@�I6Z��Z�C�Z����`J�K�0��²�y�f͚���C��Z=��S�,�La�=n&���}�w�������b�:SP9�͍vv��I��}���� ��0��(Gu�����L]�"a����}�`S�ו3�O�ß�����Q��[f4;"q��ꁑ���VOOWw��^g�|�E��'�ɕ�|���y���f�	��U�U8��,�i|r��y��G��|))�M�Zz��,sY;����KD"i�8�n��.��(R�m�ć�ԟ��C��4�9�/���hW*Z����n�Qmyh��0����W��0N_����ԏ�Xd�����Xuz��<�NG�/a�S9e���ŕ��a*��c�op���)�˱;��R_5�B����wT,V��B�,lA��v!I��7���ܬm·0F��-3ޙ���)�7�b4,C$�B�C'�*X��B���]�;[����a�;0�-��H_�~?a�\��	u���z͔e
�6`�V���dSپ<� ��95���v�\6�\�5�bL�Ý��N!��cd~�R�s���q'��Q��O���9�Z`���T��N�� !D�/�u���w�*���l���Q�>+�!ES4�6�%%	�F��쿍w�_"W6�00�	�2M���0���ɉЬ��f��',�-01a�JR��"_t�gAc���ט�uG��4h��p/��ˍ�U�'c��@�3�55+�"I�U0��j��Z6��&.>H���I��t��03^J�� �'�|e���m�(��g�� B�"�#�K/Z��B���Sҙ�jy��i3�_�i�D�MS9z�_����PBa�����	���S�Z�.ҭ�9^l2�[�>���9u�]A�\�3�D�Y������#�+W���^lH�|>�c���	~>��#���_�LLA�_~��w�q�ƍgff�#� �����*yP~��_C���/�B��,�F=�K�����{�uA�߶m[���͗|��q�+��T9up�K�`1#Q�������OQ�]L�3�ySS��k��q7<�u�0���o��`K�tg���𮓲<�Y^+)��/�0p��,���Դ�[/�\�(�-T+I�K��ߏ�<%q�H�ދ�-pC"z%6/������[Y�<��(����J�ë?����ǞgUD��J+�3
{/���q��G�$�+9����)�\t�w��W��e[���]��-?�"#JXG�~儖&_W��ӱ��:��|3m��X'��fܠ��k"tN�N��9Cj��-	�GO���D����K>���M�,��lie/���S��Ep?�H}��h�+s�ej��*$�;�~�.��IE*:�%3T=[�u����`�򛜤:م�}8���)�#�/�̌F3�)�Z�١�^���Ko>�M�x���֔29 �B�|�~��Ƅ�".6��v�;:*�&����9< <"�d=�=��t_�:����a�e��7�J
�����S$5y��*O-�Ҹ~�觚�衚,�b-�i���J�Y������%�ʲ�	vE9�a��j�!ΖK�V�����S��Ӷ��;9q�.��顛Lj���p�>n�|F<����1_�={��d�V{��'!���� ,x�JZi�����S�)� (��~��P#\I��&G����&��@s'�ܹi�f<���_jS���q��7�E��@ٚjy��(A���&�|��W=
cG�m���)kݦ�˖���X�ett��n�Z�7��A��ժ�b>�j,$<�.|��t�������H�۲r`��x���K�]�PE��S�2)wuΎ�㊔��^�Qe`�|Q�u5Tq3��@�f��"��↼ێZ[r�ZLy5�$�U���K�՘c�D�d�Ȧ�:�1�)h*�j�m�Hi�;��4�YE��������B�ͥ�YH��I�jQ�2��q�dFG���ߪm��".e�?m�ZB�b�GmӠ[�z����o��X G�nZ�˝"}��+�P�&���G�טu|�([�4����D�Z�t���:R;I#C�2(
�����S��cpɲ� �I6�Υ�a����&��1�'�FjTMc�bΐftȦB�� ت39b�8��[[���U�m��g�*�1�[��q)���Qa�G�h���xV�"���2	ۏ��3�W6��$x��$`IjT��j���a#�����>�Z	n����=�B-�@����ysͺ��?
m�L�ު��.�����^�h[GzLx��&!�x%Ze��	%S�:z)���Q�xМ��K�Ζ7�Zi��V�'4)�t�%m+�d��*�A��$�皥.'���}J��d��c�[�����|^�ߦ:vY�!�~�%݊r���������?��D#L���M�`<7����X�m,.sPJ�b�ǐ}���.�JGG��R�
�V�2�����G���(�L��fꄯ[,�>��~�}IN)�0���'��L�];x���X�`���6l8r�ȹ瞻o�>(p$�����:.�R�jRi	֤���#�������4����/=�^�+����R�j��%��~A��⋥��
'��S6��(�{'�PHg��)&�n��
�h�]+��3�҉tO5;K�/���Oj��y�5
wO,<�o��V2[�F��&��=�81�Å� �`/�x��
�z���!����"a2S���i(o�o��8_@pz�ۯ%��0�9b�h��,:J�X��
��M�E<�P["A�;K��ixz�$�ʌe��`�䇱Š�b/��.�"\,-����]W��;J��`4�������+��A�K���[�疂A���]#�fl��(3r���0${���+N�j�	�j	�q�[v� �-R�x�B	���]�ϑTU5�x$`,#ǁ�J�6�EE-��?&��c�"�k�tͷ���qJ��3�aL�$�ͤ&mr�vc�:�:�c�!����C���
��������ЭM�M�K	��w7|w�'�4(����F�Y\�®����V�E�dr�#1%�Qp�ի�h���`�_mg��W���4����$
k�,iz��~���?�*��ȧ[��3��ꍒ#��k��=��0Z;�(l9�/	/���W]5��P�@�]�O�`�b�Q�)�hjrN��+��F�m۶e��Y8�֭[�I�e�����v��q��q|� @?d����(���[�ȇ ��±mN�\*�e��]����#Ɠ�f������IC����1�N�B�"��O���j>�*}��m����N�h�ͨ3��)&�.��մm�|n�4﹁c�,�#��4����/��+"���<_��p�$D�BX35O,f�9�݌$�6H ީ;$��bӪtb��o�#��iz�����ib������d��%��Ajq� CAL����c�L�슉!*G���{.��2�\#����?)��!Zע>T^|H9$R�/�#�6�1�I*=���E1�~cn�ǻ(~���V�5��[�g<�z���{�p&��0�[��!�&J�&X��&v�&��V���e�C/T*]��Fʣ�7�!��v�+9�Fͣ�↭��J��sG�Ig���T&��@�yj0�ӎ�Mۅ\:�IS�{�4!�#K�ؗl�+���A��+&w�,`�g�/��"�7^w!�슭�����������=.�O�ěۡ�1�{~��TZ���b1�!_I�'`����L$B(t�o�q!(3,h�-������Hl��E���Y���o�ފ��%ّ�Z��l����K:'�Z�`�ACkUa��Ʋ-�^�=
!+���Gem���خ�\o;��R��e��#�j[�*�xpR��9n#����},�ǔFT������u��.{����-�;`,P���4�o�}<?eA�ޔ&�с<ň�L�i �¿�5�dkX\�R�J�3�(8�+�܆��B��:55�z��\5��8�]ͧve�-�����_�r ���fc��~P�t�,7Hn)�/p�<d?~��/¦ȓ]�v�&�V��8��<��+K��8�U�8)�&ml>�3������y�ƽ���|*����.��V_��{��2X��M=B��V��=sɻ����K��mKm47^�
���練���_�|[)N�I^���$�b`E�Hfz�a�x��Y�.g
AB���Pc�/�e����9����xR�[䌑�H]�ө\V���`�xI[_��F���V�|?��@��+q2+j�*���G�\�H�sg�/��J	l1x�A	��Yu=�t�����[��Ǡn��$�֖�`&"DI;U�h#����h5�I9ӥ��f�9�;���[�V*j�Ц� u�QZ@,�����%*�'�^Qp%~��LJ�-ހ���@i�Zj^/Z=�c�Б�äX���va��s:�2���\[����,s	��1,?��Q���h1А��F��Խ224}������!�EEA!��bl-'�ߖ���g_�U��yR��}����_��`�7������w��o�4_����2V�LDg0�T�����ǧ��gܗ�`P+[�ʭH�dA��/�1�RᰆQ&l�	������`F�!W�P���j�yd�rG��sq�
#u�wU�E�.�'bFr�j>��s�� �I[n���3-�O����sM�9�������������^ǎ�P���"����+V��0@�>)��������X(@^`��K*)�R�y�x��)�f��^�~�`��HQ8�ԗ���������Q�
ӱ�\�F�%.e�og��7)��ܐ�i�k���j5�����:;:g�3H]�\!��'�fZ�
ŧq�jz�fkzf��i���mn���Z�B�*���cS�&��p��ŌX�8$�"���0Z��|�Y��6-FE�|,�Ie1a��n���V|��&a�����x���J�X���oC�@<��'I���L3��.5;;��5�-���(�4q��`D����0��ʭ��$0�[:ŭ{qC���
��$^��Y��|�A
!+�4uM�לt��_Ö!'6�Vt�WA�W����>a��P�:�Xi"�T�Vi4m�");ش��M����@���*�'+[m�+yࢾH~(�^�J�zj[v�V����tO�j��q�,�F]H�N�[�n����������CH�@i�� So�iA�yS����Q�pe��qm'5��P"���J�sdjr�!PJoR�mnn�t�M�===Y,滻�M����0�凩�i���3J4�;[儨'��.�PN����D��{?R��f�n���&>��C�FgSF�
��)tΘ3�h�Bn��-3c��k�ͺ["���b���I>�!xP��@=٨�<�`Kx�F�\���g;�G�~Fk9,�M�I��#�j�E�==r�5��t�1��|�g?�����`�/��7=��|������֯�O?����edzE���\Z5����g39�s[>����=zdhhf��ه��ckz:�RlH9��k���U҃�XJG�ȓ�.�(ÿ̍Ȝ�����%�Qu��PӢV�R���H~$�uR�us��/u�:��8���4��Pe��a�^�@�7��hSOa�HƱ'��Ym�|��Ngu˄��� c�?�3�u����6���T&��Ė���AƷ�F__������RW�ڵk1�ÇK�<Y{pf(�w�޺u�ʕ+�Xr<���&� g{�* [[6�07�=������S��-.k{a���
���/=N(���,�A�w���2�Äڥ���"V�y"S�O)�*����dm�O��(\?W�2�1�CK��t�z���GA���r�;GĤ,��w0P�th	3|`0T)!-K�|*===�)(RA��Ku�I[
�0ھ2�x�"%-��EE�k��n�h�hNt� n�J�@�Ҥ9��۷oO��c��ot�Xcх���$�-�e�>���*J��cò�a"��jU9/z��V���2��Xn%�����C! �����6��ʽa,�3P�� B���L��
Y/mI�?�vKм��I�(�I��ta2�lJ=����4���#Hx��T�@%B
͇~4W��kCrJ/fu�OΰǛ/9�I#^��B֑W`�nHi�,�Ā:Kk\1��eA�v�u�D��P	iw�(u��wc�[�����Е��Oa���Ɵ�9�Lh�GGǏ?���eiVݭ;"�~�Q�,|��7��G�̴�޽���?����:�w�w�_~�u�]�y�����_����>|���}XC��H�e[_RH�� wڴiv=�$��&��u����pR�Ӵ�|g��9̂'�͉� nO9��&����%N*v�X��+G��RuF�$*(#���c�aE$�NZsEn.Y�'�C�яW�e�����;(��<��9眣R��8�Lt�EJ�bbF���TC��P)����IUJ�'/P#KJ�$K���%g|�� �:�&+���H�Q�5�����?;3��Q�|=r�ܲe�)����X9�G|���`��'�<n�B�N]���$Ԧ��J�\�زo�5Õ >�7���+j5ἧ�DnTb� -�#RT��اM�#@(�/��*��X�b�kqꍚ[����!:�������A)R#���+��<x���� �,�\���2ʽJS��\9Y�yU7���Y�Ե�R_~m�["�$)!PF#�$9��g�`ک��A�Qӭ��� ���M�;�􏊐�(�R*B��f@8�5�Ӛ-�x6"��šn�Z�0�h�8�(�MW-��^ƦE ȝ���|#��GuR��5�3��������(�E㧍�[ԫ���8��t�9��*�+J�"v֕� ���1}�(=N4y�mi��Q�e������ެT���A#DȘ �{�s�al|Q�qB��(�����_�i1��w���'�.����������6ɘA"}d��t���F!���k�D��������L�L��z��Ei�z����z��d�l�q�8�:c�| 4cp�=[�	����������ӟ�z���4:R���.|�_\u�=��ٟ��/�޲o����x�o֯[��6�/6Za$�XN�\s	=�/;G��R3>>Yo�\*l��Q� =�{�B�ZT"??���Y���y�!)�#�G��4��w�.U�qwk�;��*��$�,��`G���TܣIe�tHj��h�A;�]1n��0_��J٥j-߳���,����\�Dj�Fx)�\~p�����	w�Zi��x̂�^�ԥ
_�m��?���BJ����a����v?5.b�����_��W�x�3$LcSP��K���v�$�F���ȑ#J�Yz<�ԗ�PS��ƚ�"�o$��C�ꃚ��F3�_\Ǔ�U��Un � d����~C�TL_q�G>A��%\�ۿ�9:-	<����g��jF���l]�I>�ɪ�O�H�,�к��1�%���:t�W�ژAi�V h��50��z���%1㒎)�R��~���B���AԎ(���ga6Ħ7�6�>�$fw3���
�Fr7�6C<J�X�>p��z�o�$RQ�x�kM��e0�?�Z��G��(��������4H��@�fk5	4��W^S�r/��O����~�����&�#���:��U�0�9�ߎ�im������U�)��-(���_e�F�D馵Z]�J�ͭ�I�������:�i����j�`ڕ �~վ�v	��f$@#���81���1eJ�^A��0�Hw��?�f�`H�Y�����	e�=���9�c�CBK��w��Ps�Dǲ�~��H��\hP*�7�v<H.���KY��3��̡�!L~G���N�����`j�~�����?�����n�:����l���f�8��?e������kl����v7�?��M��g���[����R4wSv��#މ�J+YB�r�yuE�����i�I+�S�^MGأ26� {Z�L�+���R8�w����-t�B��6��V���'��S�<j@ra����#2����+E)�PI���t�nu�"i.Yb�����*��D�z�4�[�"�x��ѯ9�kUFRo/u#|kv�V��w�\���c.�S#�<[�V(�222f�O�ރ�U"arj��H�vjj*X��$���,u��D��Z�Xl��������kxb�#]�$�1)r]�؜���D�&I�~jjf��ݓ��۷o�@�N;[8I�2�ʔq�0U�4۩^1�c'�L�ԷH�@D��m|%z���`���hŃ���tY%H-�c�;��0ä_Aѐ�H�TR���t[��
cG���^�U���SOO_�.)�+�d�R+��qqV��W�i��\�ʑ#D�	��E͓Z��*v��f�Ha#�6�3lD+�!45�o��rKQK��-+��&5a�>�
�&pj�	��mT��*к��|��f�������-F7p�吚6�B���t����A��"� �p�Y;$�M��r^��|���5N���p[MX,'���Z���&�:�#�e�B��ւ�'��0��0��iޢd���(LW�}tV<c���?�U/��-���y�����ʱcǶm\ռV�r��/��ʁQ�xuƠi�8�!�/�o��>X�·��3���1Ȥ��+�N�LO��b���V������y�gaB]�]�)��|��޸v��L�X�z�\���է�Fplt��;�����z�����I�g �L��\�L���Ѭ:$��C�nR��$�fppp�͗���x����^�4}�Ԅ��ſ��^z�>�nq`WP�C�׷~O�A,ʱ�4J�s�������B����t��He�8�����[8�#�Ce����u�y���?���RN\��at�'0��1�l،D��H~g� ;A)�hd�8�lټ���g|�p�`�I��0=�X�B!@�ʤ��ڵk���Ea���f͚���7�ׯ��?�̅x�K�se'���{�豨Q��ң%$�ؚ���������b�"�0:&�1���kEf˖-;�mڹs'Dx���Τ\N��������� ����[Bf-d0_��vAu��������=~�I�[��f��c���˸ؗO���U���fX�_���͛7_q�K��՚��`0��O>�d6�c�(zV��,�45��o2���T���9�A�G�[��a�C��@d�>�(NA3R[�J�>22"'%a$�ʨ^�1�%�Uk�QUy�z�H��"_ͳ�W��S@�.�~�c�0�!�@O�b��\E�ۏ?m  ���H!6���pl�lNh��D�	�b�;��Q ^�E3J(����-�=t�D�d}���ə�i�g�9���\��pMG�@��W��|_��8�ORr�&�8à�ɐ���o�3�����JNMr��
��^oD��D��tt�!p�$�j����Z�0Ο`$��eD���z�/G�BkR��'��'�|,+�G�[����zvy����zl_��P�.iw�~�mqM�ӧ�wK%��}>���X�>�{�/:C���>�ԗ�t�ĝw�	����{�L\���bQk��~j,<�)8�N`�������L8v��K��ԛp�$s�`i��K}]�Od�'O����t3d賄�$E���ͷ���#ϔL)A��ch�WO9UT�����j>z�h6G}x;�0�YHw)ɓD.|KB���H�֭í4Na��8����(m���'Q/ [�8�5k�b$z\(��x��� H05�ё#G�n<b=�� �$�j����i���9rlxtR��w�u�Y�7��.��pJ���;��׾�u������C����3P�Ri;ղ+5���F�U����j9�x;�w��>�b�%�.�}����������~�k^��>��<��}j���.�W]u�)��ر!Ŷ��S(�K�0�R�)&��EH~Wg��H��ӛ%_\rll_?���;�<�ڪΉ�-�A__���x�\�R�J�`��$"2<5�~Q4<1��Y��Rog�����W�:g0��@�i�%%�sE�\2���,b���Ta�c�h�I�S�	%[;)�L�f�����J�J�q��X��~i��Ds&��Q��m��@+�Ή��<i�L�C� ���J��v:�z.כ��t��_L�Q�2ݎ�(����IE7��N0�hT�@����`�i��Uo0�Iidb�+�/��X0X��f�tʱ���|�#W,�\�,��b��
�%�T;��-Ѡ�m_ �9�W7��E$�,L��'�n�b[��L4�M�7�����V�2�"�$7���<�H�a�����z�r�m�3�%T���2 ���ޔvI�KG�T�O��o41F�J�A��0Q>'��ς��%����Ǵ�|�K����k_t�����/��?~f���7�|��_����_�rgt����;y�%�W�qE���,w9Q+H$(Ds�U0��.���W�Dʈp�S���a˥|����d?(�E�j�A*�?�]f���$���h;��P��&�E�$����|��L�HB9�|:w�ƣ5��������m9�ק��F���rr1�)Q7Hn���SU��xXq��tqV¤/�T2KZ�đa����\&���?.�bq�Es�(E6�ή.|)�G��x�9���y��СER_�i�h��_��;<�9Ϲ���_r�V:�/S��=�^<�b�07�x�	L4�_�ݞ=���J�
BK#�� Sy�}��{'[��ļ�8�QI���N�$̌�$�F���o���w���k���ǏkN��i��9,�i�����ndd����?7�x�g����)�����-��IUL)4�jb��J^�c����������7�u��߇%��&&�zzzp1&s�֭o{�����?���6h�'��ag2���L�.�ǅ�A���|)������-���z�@R�(#�'� �@j��us���043��۟c�G,v3��l�T�Cic-(B0�[E��DlR>���	
R�R4��������=�f_�2~���X�E��>ww�zѢ��s��jl�}��I�Ag6r$r���ȣ�tE1%���Ӂ;>*Q�V�%�P���YTң$�.Ig)�!�aJ9ŰZ��%�K �U:�H�:�Y��7H&� ���9��]j�뿃�K^=��J���bn��`�$л��,8�G6��G���$NVĢ}�i!�\=��r�L�{��'&�r�WN��g����������|b׮�]�]����������m�{�w���ݻw?�Ėիכ����tpp�*��pŊt[��r`�(�&�q�1!�����tQ.Cg��YG�]�N�@z�����o��Z� �-�K  ��	m��,��W��BbB*�\�$=22"@�����T*IT�a xp�\v9�� �ΪU�p[�k�+(��|�N��,�k�3�l��1<<"��z��������-������h,�@�������g�X��e�)\�5��|�� A~6�=�O/<m��+�
Yim
D�˃йO��{A�}F!�Km�F�&�N:k�����_>��ؙg�X��h3�n��[��dL�c�.�0>�|6M�3ۢ�ض�T����W�5�J�I�R�-�Ʋ	�O޷�q���
�Ν;B�q��klZ�=��Ӯެ�S����`b}�?���o��W]�j,!�F:Ӽ���4��](�j�:֣�3*��D;`���O7��SYR	A�$Hq`�U�gJy��C��x�-��z������j��J�:3C����o;����k��o|�7�p��'c����.�Y�B�<A�0!��4
d.���A6�X����H� �@��LG�|�2Em׮]_��.��$���{z��UrD_��_��W?��ϯ���Q�N� L�9r�{�Cx0�*��[M��t�R�X�Z��k-i�i��8˞2�͔��5k���ɤSVN����\]Qk�;S���?z�Uo4����r�R=:4�z�����o�t�oo?�s�]�ǟ};gdJ=}����D�H��e�I'��t�XA�Tޞ�~�9��2���	<���/�/mY_�9��u�4������XS<�;� �=��I�����������\�Ѩٝ���XvW�z�}�?���{3�ۛ�"�V��U�q,�<=uk�t+~ӁA�k��ms!_hA��-������]���	���o|V���_���	)N/N��u� ��h��{��i��� h�#G�׮ۚ͐+qv�ɍ��ۙ�.dɭ�9����mӰLz;ۯ2�����Z>�Yp�<�B�Xd������`����$M�-
��ZT�I�m$�&��Z��
5�e��"���n���a`���ww�ds���<�zl �P)�:��:5	�h��WX��:��]QugAW7}s�����������m?��7~c��^���Q�x�E���֙ӷ��聡s��r���Ǉ������_gf�\�53����1��P3����^�p �<m[G��Q�&Á�l���,���r��O�=��E�Q���E�V�fY!N�{��rܿ��_����Bi5f���v���ͩ�I���5�k 
�z+4	����))Xk�2F�JIp.w.�8
���ߖ�I��6YTC�}Ν5s�7kff͖@y
��6d�h��8Y߶f&B#H����Ә���u�P�O��V��]�m��|��aH��R���q���۷����v����cW�Z���1K����ċ�� ����=�S��E5�_��lL��2c�C!��x�f�'�Y�p�F���*�up7x�d�f�s�<���q<5`�z�~��^tх� ��+߯x���PA���M�'^@�M�N ������a:����]�+Ӧ��W��U33S�?�8�_�{��@���ڌ8�%ǞZ/$I�������q�n%�j�F��������ϓ��36T��(zILK��1C�>_�r�����z�s��\����G>��Obg�y6���of���Dɥ��(~��jK$�	��M"����!����G~x�M��G_�Wtv�`��Β҈�0��N��.q���B�_�ܕW^��w���;�ܶm� BH�f�Rx�����H_��,U�.��3̻%{��s{o5?��#���Ї���:!���MJ�56��������������<�p>���̎�O��%�:E��4��P���Ĉ�K�ߍQk��a�R>-;�p`�rDn@�MVUM*'3����Wn{�߼�6y1u�b/�N���&����g?��xׇ/��d�Ѽ%�B6���Ӕ�,��)RM����I��=z#l_�?_��dS����6�. ���P�{�ړ�t��elX�p�B�O���K����C���(��洤q6��
�1���X��m�]b8	�R�r�J���f@�?����T�,堆�B>[+���#ࡥ�������G��_4v6��J��f�@�Q���H��N3/MsB���u��0�V+��l�uI�a��E
��f	�.�6ǑQB������tL��޾�j����{�t�Ղ<���U��R�Pd�+A��9�������{�gݺu �{�s�Ǯߺy�Oo�9��⳯z�k>4U�/���b���������kA��U�H�QG9.�����C=v���@gG'����I[#M]���g,;4H��[1ҳ�|�N����~�i���
𛒙��BhaJ���֙���Ȳ�"!�?��+VW۸_��M¾�vWӴT~�p6K�l�z��3����̸U�2�#_Lcwp�/"<�Iu�n�H$f_�����\�%l���*M
��^ �1�����F��)��ϡ����AX�� b׃0���R�/����\a.=pg�*3������|3�Զ��}�5��FFF0�O��u��A�h��!g`���Z�*]r��г��~�e��u��`$��2#j�|��/�� @	�k��<iY�n�̗���%1��������\��`<X\������w�u�K^�k������l-�t:�\�H���h����\�P̤3-�����}�n0������������������>|��ԅAzud����N�_t�q(]��1���4����c{��^��ա����E�a<�.Ǐ_�f��m�N�w���g�}�/~q�g?��~����ƍ��]	s��X�ԪI�i�8%�A��dfɕx5���	�����z�_��O\��btg�O�Y��s�.�:��==����|䃣��֯�Tgߚ.��х�N��ҹ|'��\>�h��j�&�{��0��F�
�R2v�!��]��2��5���|��d���������]�2^���p��'�n�����kc�K����7�^��?��u�/~}�%��L�ˣ�7<�Ⱦ����<�McG�y�-�|���f3���`��kh�U(D��FZh	CG�:i��p�yn��-�ְ@��Q��g_|��-[�X�eA�r[���\:��#��z�~�5����n�Vv���7���a�\8�k6�Z�79�]����(J�N�0���t~�|Tt&���Q�k����a�ö(u�znkx��j�����v��pYrQ/���;�㜳wB/�+�*�� Z�R�;����Cg�]��2VYD����2SLJ�'�uԎ=�;���@�ݹsg��@�:GZ̀�y������s�W�%܄2C#Í
k����Do� �l�~Oo?X9x]&�o�����ÇO=�4�k�)��P�ׯ߈Q}�e��u��P)ff�!�Ŀ��u��z�9������Ѩ���=>��jt�<e��o���C?88|pǦKn�ѿ��N�
���~V�y��c�H���M�>k��2�E���mb|
K������'��t'֜�rԹ��6I���6����7� {�����.�
���-�딽���#�G�~�=(4��n�'���l��}#�wlzt`e��U����Z�U�S4�f��d�^#H�xB��}ҩX��j@���:C.^͠�s=�r��Ӧ>ٜ�`�V�������]�M�5tUgg�O�3#�B����X.h���/��)�:��f�J���׭W?|��	���O>��y衇�W� �^O�z�Il� �Bg�ʕ������eP#p�h�=�%V�N�E	f9bY�=X;�F�t�BW.�z�X2��ο�x*�/�+�۠�`�$�\�O$FG'���+��l6�����V�`��9]���b��fY�J��jI�5�W�>p`��]������\&�y�f�)F¬�+�uA�q=����E��0��e�������j��n�	��Di�?�8���_ԑ���]��eN9�����?v|�7����������k5=��d$g;�hV�� �!U��ů >s�&�Z���W_}�[��֓N��:%lK��@̳�&�k/S�5��} ���_���7��Z��~�K_���Q3��� ��%!.�����O4<��rI��dp����.��·��-_|�bҢ��Ͷ���w_0��T�4::���y�;�y�UW�����wn���&� �k5�w�55�P��+.2�d��1��R���yQ��|����ѳº������W������Ż ��Ci��`��~����[7�~�m]t��~��������ׯ[�iӦG}�4˃i����q΍��ȘH9�rf�&֭W)�L�t�`��xD�Pq]���Q�y���/~�K_��cn[��¬��������PJ�}�߇�������[n�뗷�uz�,����h�jq�u|f��h2
.����T�Q'�V�m�
�gDD�A��F���p������>���<GRI���/^�ַɪ�n]��˱;�D�NK|{�����$��'?����vqꩧ��E�Q���~��x(�4�5"�"��Z�b�$�BRV����(Q�9t�{��zn��ܰa#xF����Oo���?�����ԧ�l9IH��/�0S���?o��G^���+������33��Jki,�+_���;�sx�1�l6_F��.�o����SD$�È+�A*���,4�d��5�xL�L�5y>::�����Y�VD��mA�AfЇLF���U�2�Γ�r,�I[���6�boxl�������&��TpS�(��U�̰��r#�\<��y�Z�rGb�U�}�>eյxx����ir���xe�B��i�~���f2�3�<�k5��F�a�p�"��B�?���6��СC��b2	#�҉��9��4����7� ��I ?�2��>��1���\߻h�IM}�<�k_�8<��vPꉵ
�SI}A#d:��Jy����qa��� ����yl�\6-��0�9��f��I�Ȅ[�������ā��c�c�,WBtr[n��%�G�6Q�ȡ����W=�y��Ї>����z�	�
-�T�7���&m�)��iP��<�L?�B
�����]�B�TOL��*ɀ}_6%��͊�ϦS��{`����w||�uꩻĞ� �F������ꂰ@P8����ɧH�FBA ��=�u�i��O�t��'���������LjhhB_�1�ߋ�se�.Ô`��ۡcG
023�_�}7h��������������v��>���\*Y�d��r��������O�'�u��Fů�����������߾�e/�Hƃ�,h�\�Ȍ�# S'���{fwg��������Svm���}�]��hQ��z��ս}���]�CCi��\�ٹJ6��< �8]�\�B�I3Hu�;vJ\���kU/���)-����dg��o۶�y��hY�R_`>t(Ԍ�k�Ζ�{�Ѿ�=����Mk��_�~��S��R�Or8���^�����:��];��Tz[��w����U3����b?$��T^l���M�݋{�6����6??<>6�󶷿�/|�-�� ����*�щ�1(���\o__�^#�u����{�_��K.x������g?�	�y�svn����5O@7<�a+<3t�G�|��yT J��x�e��ʮ�+.T���K���ju��R���y���)O�j5�V�a�e��ї��r����|��ꬳ_���w��@Q�]���ZT�;�\��w�"�������(O�0Y	�!��އ�ćg=�Y؃��?��Ͼ����k*�*?vtdr��۳�qr�F0U);�i�R/���=�cc0�a�!fF7m���ڶ����^�z�s���zڿ�/���P���w��'�m���믿&q1�<&�6�j���*�eGg�?���HX,���"7jh�.�r�.�o�{�i��n�������@�ئj���[~����;NJ�oK>�CG��V�\�P��W��T�w�����'��nq�R�7��4z�{���.�؀Y䌕Z��$"�Z�Ӑ�>�#���B�[n����b?!�Lg:�.ΙP�<t�Y�f����:N^Y�螞+O�{{�_��܌�����]@]���N*�� ��a���f�͹Y�ӝӥ�_Kk�:xw>Ex��ϺM�.�6�}�]d��g��:;�9������}�OT�_,��Ra=�X�%jI���|��f���\���O� ��7Wc�a���)EUX��g�ux&��"���5����D�Ġ���@�CÐ&~'>z*�/�' �PH!!�HB��Œ��D��b�E����8RND�e���۰av�m��v�]����U�/�˯��+!'֮Y'Q�E���b���>@I���~���]v�(od�����2Y�'��=f���^�LM߲(~��T²{�|R�W_��2Ҏ���M(�?C >Pc���7\q��α�c��XAb[s���ħA^��	�
�%�\���ח\��!��``x)|ft��AY2�mC��[�BÐ,n�%$��	��qs��_��W?��O_�W��să�Kජ��ܗriY$�-�z˭���s����U�JSo���)#�?�x��X�ɲ���<����0/K]�"�gv������r�|�]�z׃���+PN|�(����]U��xG� F���q�F3e���J��O~�K_�~�V�Sb���1?$m�<W�j֠M2�u�̗@��J���a
�g�n��7|�+��_�<sr��Y3�]�����$l��6c]h�`"S�{����%oRۡ��@��ٱ�#8󲗽�5D��M��3�W(x�t�ئgg:j�t�tc����}���k�p�_�'�x�;��.�ً���^b�E[&a�D���b���7�t���#M	Sss�SY3R�'��� ��U����G?�>~�ʈa��c��L�A���Q5�	l}+��wB?P����z�����Mo¯7����w����?��׾��!Y�6�2��bG�3_�C뀡�O�'U,B%���N;ĳw�ގR#��������^z�]�]۷m_�zl	l�뮻n��u3�3��T��۷�2[�w�a����/�J�ǟ�ɟ�
�1��"��{��~�Ɨ�+o����o�Dn�B�h�ʹ��V!�Ra�H;+C�J8Y2]�\lv�ن	788(hq�5�4ْ�<UꭴO�4�$"$�kЃp�ᑚ����V�\�^�y�v0�(���M����	���Z�Oo�� YM]��}��7٢���N��b�&�a��sx���\p�i�Gǎ�����N�:�4&��P�@*�!=��'��yj�����͛�(�ƃ�B
��O�5�EJ'P��y��H�W�:v���g���J��Tz��O%�}F���7�J@x<����a��V0hIGE{>>�W��w�ѬrBx��jlݱ��=���՝8�ݕ�fV����F�}�~ׅ^����)�P��k�*<׷lS�������u�!���E/|QoO�����{�W�B���ѲBU9�<z�$��_�rc�6-�FP�9�&���xSHS\��������=��!��o|�Ҧ͑�]0�3���n����t��g�[=z[������_��_�x?���Ȍ1õ�$�W�+VRq��n߾���������RA��$c�P�n\G���8��za�����l�;v�[��� d->jq�cx��BA��g��]~��~�_�t@�XS(:�Vs�	��:L�����d��O~�E/zѦMT=,�vl������zr߄L6���Ӧ��bX�V�vR�9�w�j������굯ǿ7\s��~��G�/��R6O)ֺ�-ӈJu5R׼z�d�d29P6��"����}�q[֞G?�S�z�K�8�l�K�Z�E��SA�1-���G��v��������W�5�=��5`Z�e�ϰo�{!���w����t��|�+���7��N�I��_�AU|�B��$FF�mZ�k�5(�"�N�����J�O�⤊��]C#�X�sϻ���/_�v#�����:3�?��LO����EY�n������(�t��v�86:�kC[7����{~����C+eRI���e��<O���S�<f�j-�g �Q�-ν��m��a��4�|ӥ�~;�m�ag�Z��\�2a�;�|j�z�����ry���T�{Y�r;��o:<~|x
����3sձ����>�(t-R�C��Z�u���=Ƃ�5�3�n��fH�+��R����.�^�����~��?b�;������ӟ��##Gq��-���/�W��`�Q�k�Ƹȧ�N������jͪ�R����GG������p}W'��W^���}�Y[����g>s�-��,����N�q��]il���I�䋭Uk3����Ղ�ޜI
����<���v��Ҳ�VÝ��K�MpW翾��b!�^�q�4jӘ7L��3�J�����j8�|"���<��/}�+]��D�~�}���'�)��l�q6��2C�3G-���U�9�:~iY/��%�OjHt��w��d�΅^���P��Tuݺ�ή�X5>���d2�}�Ml�<�j��#�����#�z3d��N.��U�6f��}�ʹ8��٘	�S�5�5�A���\o��_E��5�ڦT]��5]eRȯ<{�2\;��]/y�e�W������N�u�Lέ�(J��17	�� ��z��SN;��G��\w��C��-[n���}X(�����?Ae�2Đt�S��
��䥝HL/J{��_�����Q���l}�;#��0h�*�x�3����BHU �2�	��
���*���BΎ��>��<|���s������} �1������ܽ{$�W���ۣ���:�~���Tg�*۶m�N����:x�0n�MƕܒQ�Q_��/�����psu7	ϋ�*L�C�8p��3va^�_��� ��K/�7��޶mǇ?�AXKd��R�� R��ׇ��>d�P��+����~���ħ��`gT%��B�e*nr�wbl�}�{���7���5P���!Wš��b`ă԰��ͧ>��O|�o|�A70nv�ܩqsB��*+VZ�N��p��o�����}����裏�zpCL����1�1�N=��_��W��_�r@]�Nsݔ�y��&w7��P�?&����n]]}�Ւ*�I�Ų$�X*�t^�\��W��=�o7�p�С�}��o|�33��R��l�}/i�Z������Dɳ�P�.0�6m�Կb��|��.�n��ؼy���G���]J��=���W��R����t���GWR}7�˳�_x:4��"��s�u��'�܏͌� R�RI�4أ#;��^�� ҅��g����N��kv��;0d��b$m��]ď�,�+���)�0I�j�
�s�����<�s`�%��P~Q$#��K��( ��p�JT��e��yfv��α����|g�Y���~��g��������$�U��_A
Xu��i��2��8� �!�������_�"�����X�8�`T��m�4��/+��*&0Y������ �N
�,+�t�ߡ�Q���fpRRi��*����-�O��I�!��>�l�ߟ�����q����/6nܸr������7�p �e��88�W#�#Խ��El6����_��x�.��*�H;�۹s���U�X�C�0�q4@8�O=�Tww���5����~Pբ�m��c�=k�2�z"����$�-�|�s�"�;�PR�Jɒ/�_x���6��p��a?n=2��⾃���<��O�IX!�be��H\�?5jA?H��e�]H�Ǘ��i�zI�� 4Y;�?��T���	�����g�h�rȳ�ϔ�|��?�����DQ=-��=Ŗ�8e�O+7�׹Gl � <s��ո��=;����^,dĶB��L��,V.پ}{p�@Xp��Š���o\k�)I4Ã+`14�;�G�dqpl�A�������|J�wj��]��ls
�KH"D��By�/������A�Q�&.�Z�nf�`?����6���aUi*�e�Pj����D�w����͛W�ZN��c����t"�K'sYJ	���.XlQ��J��#WE������-7�Ch\���]^�Ϡ8D�CO� Jz�!�����z�������s�s?v����gѢE�\
��#�<�����A�ݻ����oڴ�o�闿|즛n��*
n�"+�������j��I0�.����N;��k�}饗��X0�J��D�7����F����_}�gM�X�X�1p�����v��g�u>��c��w�}�:I���X��ʘ�$Q��q$���QpA�)x{�x��?|��W^��{�6(.��a-�c����+�.Dh�p�|�fJn����U�e�D
����7~�P����~�aM+<���s6����Z����V"�P�������ڹ�4�����飏���s���s�vΟ;�-ev��ʢAY�J9̀I@A�\�j�	}?-�o}�K_��@��r:]����2
z�n�"�%�h��^�f������M�Gy4��@C�$Uku������J]��'S���
��K�ٱs�>HG}����f7�ԝ�+���k.;����C"Id��#�)�S�t.�	_<�cX�J�ɛ�%$YOg5�
�LL��1�.��n��߳e���:ɠ�9{���@��Њ�,Y C*�T���;��ZZV��rQHS*��1_��]K�<�
c�^�-4 ��	K�JUK��)�1=cѨ�z��p��gʥm�><2

���AkΚݪ'���UUւ8�
9j��DM]-I��N��Pw����f�6�j\<<З2Z�ݒ�@��n� jT�Z,���++o��h�#�:��$F�9s�BÂ���/ZzءGlڴ���o?���ce�r��8�����iA_ptx$�����f)�3>>:��k�4�'�M���t�q��عܾi�:��>��T2�-� �|؟��V��}��׍� �����?��k��ɝw����~ࡇ�[��ʾ�!�j���-Y'F���߫Uq�*qf����;n���˯5�8V�yݺm����/��eh���ڈ��h�pQk�N�}�������f��ϻ=��7����
;��;2�Ք�9X��0�����^jz�1�l�멧c��
OĒ�Gl!�b��9ZC���r����ဵ:R3�f3�m��Z[ZV�j���7��
P3��MQݫQ��]�L��d��7	q��򔗄��O���Y}�]r��#��Foc����sZޥ�A�.�8���۽mŬ�k����i�<�h�	�5O�[0�M�&`������qxw�؁�����V��y�.�v-����up��N��7	�;����1ܸ��#�`W�ާ쒀0�@� ��cO8�S��Qt�U�&�B�����Z_��E{t%�c~<��R[��+�e�1�s�zϾ=�;\�����ii��җ�T,�<��$٬Ne+h�T�#����'�|r�i_"�R�� E��d{���].H	=�$Ժa���s��_�z=�KW�^�3�%vk��"��?�E�?�L���!����ʕW^�cv饗B)�r0M@7��^c<�n������o��C�
�80�!J��{<�.]�����I[mК��0��D��QX38�0w�$Xc��8�pM�͛Gͩ9*��>}:H�_���_��K��Ǫ�D�_l�}�@4HC(K��ڵ`O>y�q������?+3�C�bNh���չ��9cMu'�i�:�����J-[�\��x�N�Q����'����?8���w^N?�s4����6e�ƍv���U����o��~�Ӈ�OÓ��p�>w�����=	�l�����������=���Y��4)�L��Qj�r�C�1:������b|��{�W�uᥝ�܃�Md�P�%�41d��>,x���?~�����5k<^;��C����
բ�A�nJ?�/l�'�9��r���8�<���lF�Pq��b�|߽���\1�ߋ+L��f���:e
g̞�q{����D�`��T�xlk�9�_��m�_,F�����w�%�%��IViʧǛ<��O|Tchز<;.V����
���
(Z^W��1L�΄V&��ð�+��t8%���ǴRF<$�ڵkk*�T{a?н/�#�2��,� +�pK<��� !
OT7������PPdB��F'��J�����8Y�t�Yz���zDCM�g�}�m���˗ϝ;{ǎ]�� ���q���t�n����n���p��q =u��U5K�?/���+����k.��ZsS;����0ˋTT����v�a-�0q)V���i�y睑h?��d\�	�B����x����9c��?�	�}��íz���I��r��_z�śo�����d.��w���K�$��K�I��u4J%_0�ݱm��@
������BѓF�j�|�a�XQ����@.E"p^��j��M+�*����e�=J��:�$�KmbL��EZ6J�;��k/ᚵar�q#
�2�-4 f���b�\sM�H�n߶-11�&��驭��%��a���^��B>���"݀k�\۝��qY��`��ǵ�����y��J<�r�ڸ,>SF"��Pj�w�/^G�*z8������O�>�����`�0�W�ZŠ� O"	����� �ɐ���϶?������?��%Ktu�T�M�d��>�[�e�E���'-�c���>�pEmI����������u�p� |}�mRs��	
B��j��?���[aa�r�)UUa��K<���0���n.~�$�_��_>��T��a�qY�%���5y�6;���#}�'_|��K.��~ ��L�}�n��Q���w�����Z�d	ۃ>���ޓD��1���o~󬳾4�����E�jbGb�q� �/Xɂp2�7�g�D�R��(¹6P�1\䢋.£�8�5����42
���������/���w!M��x��q5 ��W_�?��O����Ie�R0���ª#Q��~�͝�X�w�z��[o���u�~kk�����r���0��<��/~�o�~�;��$��v:��}���ڦ�^|���v���~׽W^u�����,Y���q଒��!��iw��v�n?���q�U5�����b��q�"��ڵ+�&|���
-O8�p���~7${SSݬi�f1�v:�Z��|��G(����]_�C��y=6'V�RWC����
D[��� �ig���=���������5���d��f8�������j�21)�O�\n;��[ۦ&���u�M�`)KF<5����Ţ{v��_y��l,��7��jgw6E_K&^y�uk#�W�njkW�v�+��6�'���04RU[esX���n�[5�x���d�d��Ӛ�i**Κ�J�r!��*ɠB�a�6�"e{�dE�iڋu�dsIаd��T)� ��������}���h}C�E̜R�ؐZ���ld`C{��������Ȣ���v�lu�m5Nw;Ut������9w����C��1 )b+R� #���BU�QT����J��H�\6��"��������,V+T>t�,-[�pE�r�	X*UU|x��Y����Ǳё��>�����Ӱ[%=?W��J%`���&�����Ï"���bx���~O�Y���6:}��߬>Y �k	U����
���{�}�/��r��p�N�Qrɦ����qd(i���D��e��
����:�,���c�:,~Ϟ]�X��|RH$�uƌiw;�+>� l��˯�\���QG�&��o�u��_�={:>�kB&� ��n�M�~�A����f��`�{<��7���Ѹow��pRUm��ӡ,z�Cktx?#��=4�Y��x[b�ѱ��l�\�h�:0�#::��^�1�Z�H=�z�t.!+(�)[%#S+��@M��-Y4W��갻2XC��:�O�P�����R�)��|�f͝+�j_w��{h���120X��B�����"�}���(�KU���b��mv7u�>����]��ŨG�4Y3rj\�9q��]�Q����&���,sjɿ���<��x<n�'j��Z��Ag�?��˵��(��!�I\C�E��#��	� /�����xI�5ᨀ,*���f�b�Ƶ�I�	Z���{o��=���'�xb�G@�����r!GX��BA��'͂T*�%0Ł���+�w��x:��{�W��1c��n���'�Y̿�V����ut�a�7�|��|������׾Ψ���F1��Y|x��ݸ�5�\�_aW��9餓���/�L������6��z<#xn
.�#b�[�]w�]w��\�	��X�#���x� q�<a���%����g�BI$��̙���>�]@���}��{��w��(@[�n����;/��R�
�2�;��D��+q/�����ꫯ~��� =X68��v
�7��ڊM����_���~xc(H��wNvX����g�u.Z�(:4�m3�<�e͚�����;�Κ��V��sg��믿>k�qV�?8�T!S��n%;	�$�zZg��ۯ��oUUp�L�j'K�Ny
aw��5�7~��\t�aO��g��Q簭c�0�`��1_啅�B_~�9P��6.�MDA���*�&��%2 �g���9��kE��L&c�	��� # ����7�~�5�
��%+&i���������CaB�R�:�x�
\G�r h"9��D���>F,j�B!out�1��b�aN���ёd6�;w�u�)F���".bwx@Z,ރ���4��I��4���}dx����2k�3[�;rB̔'O#��4�<H)�͛7�s4�����Y�`��UD"�T�L�M 0�ђ���/
�Ա/���z�Ikb�Xd*��v.��y���h?��OW�\�}|衇����F��L�m\X�]��ໃ���(H�u���v�ʾ��]���ޕ+�8�䓅�4
�dEB����v�W\��?�°�I"�PߝN�[2��u������u�G}4Ũ`�s�=w��j�.4e��z� ۷o�ށI��7]�|yA($��wa�vvv�����Y���1>�R>����M����h���Y�ѻ���r��ᨮ!H�SB�}����EQ�Ku�\xĘ�{�ص��Ƚ��H�q��X���j����L�eXmAj�%���\=o��+;ϗ���+,Ne��uO%c���<��b������������	��d���b��!fB��C�r0��N����s�'����g_ߜ�c,B~�� �v]Q�����Z��ox(��u� DT��t�S��5�Y��^jgg܏��C���z9Cqlt�Ҋ��>�lu�aSi�64�����X� ��.��������w�}���nx�����V�X��Ie(�'�sZ��;vƤ�gk<����n����(�I��.��w�\�v͓O>���2 <Xd`�/_Ըŋ�����+a�D9<KRG�"��x?��Shʍ7~�+_9��#�����\� ����Q*��t>��=�hN�#@J�	xM�T����d||,:���H��[o����XY�^7�����K�l�(�����f*(���{�|�O�s�v��*\Ǭ���q8
�Y��o߱D��5W�}�97�p0��SO=ߒ�e\"����)���q8�>��_꥗^��׻���6�JDA
�>��$��\WW�r;^y�����׾~���b1�`����Ig#�Z��6�����|����p�1�7m9	����s�Cen���~}�J6��y�LN!���eP��68�E�����C����k
���y���\�h��Z�͍���7�-4�T�/�����k�w^u};��ihցD���'�9�3PS[�����;v���(߻��w�yg���F�|k~�X��5 i{��h���O����L4�42�7��T�](d�̪�m�h͚5v���\m�uUNsY�Á/�Į���|���cO�����'�p�#DюbV�*��˸�!���`�����N�B��j]FF��laDӝá��q/�xj�l��A�;>/٩��7�,�3#<�HQ\=�	W#\m2J猚�F��y����l�B>���t%{Ӧ�+��Xl���s�Z�jټ��y�C/z��L2S�ԁ������o��}H�3;4]��T>4?d:�tS�txd@V��{tt��2����7�}�JƱ�Xj6�9�t���vo-�	���9�C�9���3Ϝ��0Js�����-��μ�+p|*+�j�����fI$�����D��Qb;�oim���K>ټJ焓Ί��7���ˡ&�����Z-nIu�"��^q������/����w`�T������ڠ]�GH��ݷR����z5u玽� ����J��6}:���|֙7�xݭ�ܾx�B�YM�A����GU���m݊�C��<�s��9�c����Fn��Dí�wP'A�H<�ր���)���%�P�'FI�9:�0tk \�;b�1YN�O�v��N{�X���a���Ag���SeL.S-�f�� 3g�iw���x8��l�֏������n~��ɉY��S*�C��w��pJ���Y*���1�R4���m�u�ᇻ�x:sx(��AA�:���Y*�	3G�wLoY�|	N�믾j�+0�"u!��\��?НN�|>���8$���q@��d/����/�����l�6N �+~I8���l����up�%C�r���<i���b����w{<b&�d�g��+��`�e�ʶm���}��Gu����={v�܉7!�gϞ��@�G*)�[�����4]n��[���|��Ƞ�Y�T^|����_{�W��^����~�b<��b��Td<f��GZQ>O�/qM��#)Ũ������xX*0��yP,`Uh�(�G`g燇�c����u==���o���E}�������}v|��S�2�,�;�lW��+ $���C��>N8�S���W_�V{㍷$jd���:��E�1Pt9+}6:pD����_����裏��o��z����ĳ�q�\�˓�xj�;��{�_1v�ŢP�Wq���8��pߴp�����ׁ9���Se�7�����"����H��)�����Nٯ��@*m�t��O<Y�ad��h���e��ܹs��pǷ�|sΜ9w�y'N���5N5�2u�l��M�)+f�Q�������q"��-kkk��ÿ\~�w�*j+9��+C���/�mvN�U�4��d��K.9�'^|�e���L�>=:2�Gþs�Ĥ�(fp�bz�q�~�!ຑ�>|��������
I
�M���!(��;�Mó\�������/��Bb�f=T��3���8b��ķr�H1�
��5�}��V~����m Wl��K�x�! �B;�����d݈
 z�[$����s�J&���:�ںFP2�Lx|�D[ @9�H����Ā�G@����ۅ{MVi����@ԣ+j�S�J�ngh߾}8wX��76L÷��$'�����C�s�	oY�|��SN9����mm��ip` ��f��(���T��f*pV�-�8#W]u�Yg�A��J�B|��O\~�����}�y���=݌k	��q�-_���~������v�}�����]w���L
*?�N�Z����zhEM�UW\�J�1�*��.*���5�c��>�qٲe���u�����?L* ���#�<餓�ɀDؑ��^м��������\e�N_?�g��E�z��---�\��tz)Ț?�ߗ�)e*�-JK1����d�4k]]�D-y�r�`�`N����ƶq. '��U~T��(]�ׇDmVb��ݝuئ��P"���(��o�Ǻl��y=W��cm� 8��15��|��>up{B'�|rc�|e��-�������`��&���{�>`@�ھ��?{� uݺu��x�w_�0<�O�s�*�|<�@���� GqK�:&2�*U#Z,\m#�{�2�A�b����y޼$
 ���������<���m���R��8*D3OtO?���W�>���qDc�d}�~��ǈ�fiI݀�Ze-O9�VTP��R6��Y��֣�k� %����t:N>����n���k�|�-���˗K(���v�b\ S�s�{��;�*���׽�����e}����
iF	��PT��Z�n��+����(�$�]^���r��Db|L��
�+��C�_�_���SW\q%|���bN�_��k!�
4fT��qp	d��<�Lm�S���[o<��#������@�|J���� ׋b��c:rI�P���.�X3<c���__}���{n��Ɯ�%��".�loo�� �jk#��}6��TbEh����� d�̙�q��^{������ߨp����eu�+T�,*�2�uB&�Ʀ��7��p8mp�M��M�\6��O�=�����'��#�`�REE|~�/��t588 �����K,��rꩧ�v*b"^D �@�"\�W�������ٹ��%�d��Lj���ټi�3Jyj���5KzA/bi�MIǇe�C�fIJ%(��}�k��Ά�=��~��\�b�d���t8<��"Ljg�Pʓ�'�y�o�͵G�:q��Ϡ��͙�h�
]&+V����T*#�m�dF�FG�\ctlt|���v����T��?�g�_ �;��s���K)���\��@ǀ�b*�YL��t��&��`���s�'��� a���*���ptH�i�@�����j2lu0CUd�[���LS������o[2���cc�L�m���`�c��TsZ,H.�c�⥹�e��A��qY���m3q��������L��ڼ���7���{SwW��dA�k1���30��9Bu8&P,4pQ.m�l{}C{QY&�%���v�ʕ+��=�<�9sf���Q_�*�4�$��&�S\�>�?wvsc=�j�6G�*S����[�>H�����ٳ,�󨽣�s�]�;�777A
%�4n
�rF�^��~���m�s/��ܶ�Ec��{ݞ��޺��Ԑ?��ǣE=%���㾰�r��� \:�5d��q�"5l�מL��%�����t�ҏ���[o���vQ�M		�T�y����	ǟM���f۶-℮ز�ӵkמx≐ɸ8|3�����,Y`Jp����#������p��Bmq;"p�;g������T��$�X6����N]��T[�D�^y����)Օ�k���5����u`d�ohD�0 U�ݵ/Q��E"�U���e�(;V�B�R�-6�͞+���S�J�5�����Gsn��Yf��wOUr(���։�x^+����$��ջ/�s�Ѳ�rz῟��oc/=o"9v͵W��+���ֲ�k<�'a���B�
 �'��0�M�aF@9�ω$���q���.b)�2����/�1�Mi�޽4��cO�R���j}�|[^9�V��'+��:pZ8m��[B�@�g;v������p��b�22�?6�t�Fi�b�P]Y�KV�E��^<TU�L9;+�EAhk8=0 ��W\q��_���r����'�$M�$�׭� V�nXC=�<�={�A]aa�6.g��x\�=��d����4����<
N#�� �B�}��o���_C�?����&��+�����|:^镲��7q`�fL\p����5)�
���x��(��+M9�bv�ϖ!}l��S	�oJ��������կ���o_r�0��aҋ� � `�fj4����qn���r��{
 5�맟~���V�D�U4���&�ȴ׋�8���iª�d]T��rY���W!Sln��٩&��{������Ki®2���i��%1@��Y��5k6lv���O0�57��c�)H�|��"h� ���O�٧kA�<iNO3ڏ�d�
%���4#�"'�DGb
��ܹs��/�&�ͷޥ�l>���y��⢶����QJ!ð �o�kޜ�.4u���M��ei��$��ibU��P/3GvD��|�W�~�E�E5M�V+����TD��B�QuU&C�!�l|��w��ؓ��PO �v���,y!����V?G���=?��
f�)x̚���5��iMF�%���<8�����%�m���¡�M;EA�Ѫ�gQH�=�	))T�����l�b�����ۇݜ�d�slj��ښ\Vf��V(
yE5����v��񊊰�`M���\47���v\y
����*11Q@����Eԓ�m��أ�}�(���P��7�v�)���������<��4�!D�=�ּ(��ynpݴa/t�o���L)�o��y-X�@�R���޿�P���L2��h�K���4Y������5�=T�$�<l8�o���k�[��������n.G�`pB!<qB�<A��@&���9�[�n�M�����n��O~b�'8�xAڳ��jb�E�ғ��� 4���Z>�5�>�S ���$�N�¹S��	nii����Ld��-��V��Im*��S��9}FeI/�$�+w�1ؚi� 4�S�կ��ןq�y�D1��>F�ƅ�A���Y�R	�dP-M��Ra�k@Á��#�<2:���/Pҳ���裏6}���c�]��жֶ�>�I�~�&�hhh`��@�g=6_���qL�����W���q��_:���U��j�0��s>qX<SM�����j�g͚}�2��	*��&�Dc�'�v��k�uΞ={dl��������.�yFG��<���ɬV�@���Sb�|.�LR�D:G���QcOR��M�f�&�jh0d����$s�a����'uYv6�v������7�|��K/�.�4�A�7D5���E��N��e+��?��_����t㧕������B�eU%y��W�U&t��"T]�r�ZY��t:]b|K��rCD��VXU�@ .����Bx�$��K�l�;t�M7��BA���V�Ќ���!ʒ�r��A�;�|��w�u%}$%syQ_��hB����|2��%yE%!R*A�[\Ŵ���OQ(�7�������h�KƎ}]���_w�{�k���d���o����c'$Z��\�	u�v�u1F2�[hhNј9s.��=��s_}��,u�E@"-�lp*����&s�|.I����x��`�Z*�
Ve���VٝK��l�i�t�P����o��������P*^o��_%�f'l�b)�T�t2��V�J.)˅*k�i�ߎ}[��OK燺���p�k�T�w_z��7��"�VQ�m6	|����f���L��jqP�	�/�q����Y3�+��1
�Y���g�~��'���w�Y��{�o}��紌��e�=᪊TJ��+������/�f ����tڮd;��� 3� �q��p�g���{�c���\,i9+5ե��T%�V�M	�1� ��p۵",
���j9��N$��L�f�{����g�%.?��r��f\flT�J��~l,�6m15)dT�����8�M)UC�f�T��hU�����|��[�k=��V{29�q*�M�Q@	8%E�Lm�1�S�ZC���n}�f�ZI�L�*��V�����Ї�>ٳ�ÚHCE}C[���Ą�8$���Pr�E��}���m[���aH�O�m�����?S}hG~;����9��(�mZ笾���u���滝$�&�=�M��5SY��L.]����q��?{���!���@+,^y�.�E�[���kW�Z�ۧ�����t��d�jjk��G�h��f�ry]�a�DԜ�h}�nM8"�ng�w��90�#TQ�7�}�Q�x8T):�v@ p�v�o�����m�?|������t�|�yݐ��/���?��E���|�-w���a+mo�F�(�{�W^y�e���F4�#O&/]-��jHf(\���B�{��@�Џ;��c�;V+шaY��$�I}
�'�n�-�X5@͌G�����F�A�j����[U�⦢��VQL7�F^r�
���e�6Ś/�*R}�
���G������?6��d�Lڢx}������J2c&��#ovc{ �ܿ.= ]6���Gݽ�{�V��תӱ�lz�����a1Ub�x6k �����i��M�X���ښ5kѥ�&�a�\�\"���n�͓��²9ձ��Wׯyf܂�3R���������K�3��ν��*��c��654�FGa�B��)03�'2p2���t� ����ve%��ɒj�9������V�xbFF]}D4\�_����m��<hA������o�	��UR�D{���`S/�}�'���kK%���E��AK�e�EG�!�BQGW�[�T�>���]a�P9��$Fy.]����Ǘ\rə_:m��%ё��0Vd�G�.8<0�}��7�x,�|�����.��!���q�`�͛7C=r�4qcc#ϑ�9�?q	:���g���Ǎ`��*�/���Q@�01��O~.ڝw�y�Yg3�����pNb�� �>�F�x *���^�{�4��T�k�xS�
��d
���T+�`n �pn�l'r���eq_x���v���qQD��E��7sΉg�9E��!(�3�AG^��p"���{ؘ�&�R�E��[��Olܸ���Q�K�㖁Ճ ��K�ʴ�2}��o������`�<�Id���S����4�|�̉��?�����_�?��~p���q��s�-�< t�46vEnL��H������s4�?�@�W���
�7��C�w�>�+g_z�+�����@(>A"�M	���ƣYnȦ]��hx#����·˃�B���n}��g�����`��Z�F�T�oy��!j:��K�6��uC`Wh���\+���PE8�Ǘbq��һ����v��+]>B1KR�@uU��p���>��J��F����b{�<�u�Ľ�UV���$�/��݋J�r9C'0��6/u%s{�lnn��������m����r,��ڴ�*Po�������s�?�iӦ��Qd�F���]P0���'䐦�\�J�\cZ��7���Ï�_����~��j!�Y��V�ǻ��?�����_}��/��2+�T�-��P�V1Gx�~�p|M�?1>�� ���%p;��&޶m[m��Pn"��nkk�����a����Z��~�=w}��_�9�� ���+V��:�{���V�^]EuBdPC�z�,�/>�Z����>��#4i��� ���0g�n����d�cr�E
bV2�_�LB�������ۛDȧ ���x��_9n�bMU� ���H'%fB԰`�M�z�\*d�Ν���M�Ys�峄ᯕ��F�VW�;7XU[tt� Icԧ��R�KE8���l��>�`���xƙ�Z��u�-/����P/�Eb"O�'8I�q��� lJPLԛk��
y�g�	�#���w�V6�O�o�l�m�[!�H؎���m�ڛ٣�ii�f����S�˕[\��}s��3*���L8��S�Be�\�
�+����Z�g�HARd�J�E�h��_�e9�*[�rNzxdp|b4�Jj��jэ����h!g��x��zl(�������ap�"F�R��ũ�O�Q\H+P�,��:;;E����?��S ���e�L2.����?����㎓D\t!ĥ`��6��v���E� �p�x��SN9�����'����뱼w�}��9���An��я~���C͚I������������D�\_ۀ�\�������ַ���4eZ��q��ǹ}��Go��v����/�����INd�?D�
D��q��!��z�>F{���D#���}d�`��&8��]�˖.�jz�����[oŭ�������Ʀ������IK0�)*X��v�~�w�uH�0�\XP���_܂�N�a�-�������9��)B��B�ޥ
B�&�Nw[S�n���_������P�E�洈�͊��׈��es�U�dׯ�������%,�{��ug���3�N���m6�R3'���dOH"��h�X���4Y����
֎'b����"��Cy���ޙ1� PY�l�2�ԨK������E�F�C��2�?h����X<F��s;A�_<t�V�fϚ��!8x~c*YK�!ї.36>�i�����P{�	�\@n�P�T=W�x}�UG/�T���נ-:����!���:�BZ2e�͗�Q��*SMVOw��®��%�`�h��Ɔ:O||_���U5\��8EJ��>OC�7�{�e��=](fJ�
��tV��]/�
��n	V<t@"
�ϰ�����[5dkQ�G�c��X��Q]�ǣé��֣�ӦG�+D�k_*�GB5�]�#Δ4]V�h ��[eU����.����t�
3T�Ec�xp$
�J�|�{}�]#�=9���B�����*i�+�Jd��DvK�����eUx*�l������#Ql���X��uUE�E�E����z饗>��ֶY_��X}eu�nB��I]�l��|ݭ����۵h������R)�/P���9��y��K�v�I�766AWutN'��h4��NL��z�T�04D�&E�.X�c���v���p�Д��E�J+� �1o&�i���d���5��`��\��B�%�"�$��E�Ud����Y$bފE�i�\�Y%E&�Pȏ
�d2.��7B����MҠd��#G�$e�Fw���P���ui_�n���}����։x��g�i�5�TY5���8<�H5)Š��z�̠i�#с����;vl�<�߻u�.�J`Ұl�������8��O�٬�SO;ipp��W|��.�.?�+a��?`�x'�Cټ#��Z�2�$|������ol�a�ׄ�����*gl��V�P.�MK�����Ҡ�����o��=��R��]�������I;@��rQ4.n�
 ��x�F��ͥ�6"���V�4"L���!�i��z���TIݻ9+��\'�h��ϥ�~7?���כ��9�X|�K���C܅�S�d���~\
��kb��Ha��5�����?�`��&[���s�=`]���r�- .փ�t�MX<6얛o�n���'�x��{5�̚5kÆ�0��@�>��c ũ��\�B�Q� q� �]^/�7a򃞜�c�0�<��z�B
R�L��:�M�'"�]!��7=s�)���r�<�R���pH���x
���ښZ�lҊ�ST]U�H&��`��N��O>�k��0`a�xda˝[�z�ᴊE�+]W�Z���¾y�7A�RQ�t�ŋ����RN��}3g6��K/��7O?s�UW����2�b��IP߰(EE� l�9s�c>���o�][����~N��$ˠ�A��%pEi{&��,�X	�mL�㹸���f�d�i����];��;�9����{���?�ν}�*�ƜNg����������F����.���/��/��!�дY� {ZUJb^T��G,>�������lRv��&�F�2q>SY�R�g�����5﯁)�X?�*\U�&�ْN� bF�[��.�Mтl․��ŋWV�a�߳�*�]V��A�`g��5!M>�YS��-vx�$\�?K����`I��) �Uu(\���������!gp��W?�c���>�R��PF��Q�ol�?>c�e2�lB���I���d�iJ�RS�\H����fG	��w�jX毈̔��x|�f"F�OUu5`������8�0������`k�}�p�sy���ǆ�x'��[���U�%�Uw�2��j0�r��9_9�
�V�4����H�>x����O>�,N��p�e@x�hr	����k��lW�ڵ�z�U?��S<#F���Ǳ�Y���$�A;��X��}&�{�﷟�)Ѵ;�����x���� d���s������ӝD���(����H$6|<0DՂ�a{�7 ���Q<�f��y#���>����*n��V/���o�E�=�0,�<*�A��bc����>�3��A�s��y�混���CC�.��#lٲE�Źņ"��ª��]d�����6��Ǖm^-� >�<vDp�}��Z�];��-���������t��MY�Xl���\�X,�x�Hm=\L����u�\��x.�dg��,�'�Ƅ�%��h��X�b�$���2HX7����<��e��4vR{���˖-kii£�عs�a���چ� uuuK�.ѱ��Q\�7�1G�241(����2�ZP���j׎#CC�t��g�1��J��_����|ߞ=������o��+7�7A�TU�y�R�uΨW�!�bkK;v���˯�z��  ����H�m$ꁍ���\ ��x��6+���I�~�ָ@��:�x�J�?L
�r�^2g�/�XL;������Ϝ9��_ �2������bM��"L-�����`����{��1�.Y|nM&j��u���ν^2���h�����VQ�O<��9s���w��AR��)��) I0� �7���"�%��R�j`��Z˗̎O�_]���뮻�e��M�6���e�ĩ������=�����ׄ�-��"�c#�MP���*MI�Yah��
��t�ϭ^ዀE~� ��b�	W�N����LQ��<��`��pb.%ڿ���zVGî]�����Uǝz���3:������j"��]�/h��h��H���������1}Z����9�ۑ�Sz���u�K�L�4�{4�x[��gR)�ns�*���G��,�r<��z��wx����]��3{�Uj������	�dg+
̀�o�I��s�aa�Ͳە���	w�Oxd��$��E�.;���&-4���HȊ⤌����������Rݟ�!���r�!���!71,#^(TUG��Bs����9�!V3�B��+�����D|���&PGj*�/���{�aw<9Q��uJN�ݢj%3�T5fӼ*MB�ir�0ٚ�Lһ����	-��4�.�h �Y��r��L%���:_����@/A]��jo�-�:�d��i�⣤h��i��L2M��l��	Q�PS[%�, �ea@�*cOI/2Ԍ�� �0NtՂ}�U�;-b�4��fW
���� _�!*�*N!C9���9CD`�����Ï�Nڸq�i�r�����f	z(q��1cV0���B���Pb��m]]0\�7�&ȥ3=��
�Un��2X6�/�%��G{�P,�y`��Zt�	�%�[��I6�b(�"9�9VG.��w����C���١�:��@Ld��!I�6P��m��5�b�J�A�@]M��e�L&3M���])x^�1_�6�sQl��ݷ^|��o�ګ�r0I��4{E�FV�v��L��r8b!���$Lg�펊i���OM�>���Nkk�
�<��c�1�K���ω��Mh������P0ex�~���(7`�c���~������}��@�p{�TYY�������or�����`h�膍���8	Pu[�}e��	���mYWY��K��01A^r>/�EQ;�I6+�~ٜ�IY*�u�-A} UT{~���]���)�AZ��cq�]�v����>Z����eM1w�"
"M�jXЎ�tpw�Wq�m�0��f(bծ[��W^a�g����.�u�ϸ��M��|�P��u�<}��4xXgyq��Nظx�9�'�ޱ	L����$�h5���(��&=Lĸ�d�R����ߏ���T��$����3k֬SN9����_�h��'�����h��r�׾z>��cc�ŕe(�c���*�@#�Wc#��=��#\pt��䬳΂)!�n+��%r9w�>�S�.D�z�7�5�;�zy�$��V��/ep�N8�/�pb�w���Y�����4ʰ���`+M��aԁrϛi�l+��Œ�P�x�N"�3/�'p}jEų�6> ��T�n���k׮������E���r������Qϑ���*��U�&ƇI��a��T�Ũ���vR�1o�x�!�3ʩ}�q@�}IIzWDPE��b�Un�$�&��������i������6�G�u5Կ����y�,�֭[q/�(�2l߾]�fE��nf'��2�D!;��$OEx�틃Od���W%>z�rb�l�d@U��FO�����V�X�~�D�M8�4j������x�6�Lp�'�`7��.�l��ī��ʸd�lS�SX&�`h�,�:,��� �d�N���E-�٦�D�h���+������Ll����4<�ρLZTvG �55�675�Sb��9� �d�k����m
�+��ZU�,�5��ոa�HUfv1��U�3珹��	Χ	�į===8k��E��� �@6�V�y��G�����2�+�B>m�~;��(aV�`�c,�����A�p�i	������_]�XU]�UF�Gi؇BK0A�Cc�봨�Ig��u�	�&&
<s���|!�i��u��fɒ%��b�����0yS�pД�2
�B�]qc��)b�yAB��m�	�����͝;��է��9U�<��v��Ig�J����*�;_x�	���,U��������'�|�J'����I�\N�?s�E�-�Z�fwfҸ���]ؙ��8���H��T�=�|0)]M�&���%��O���,�
VFv�	�p��$�[��FG(� &�1���B�>*�H�^�¸��B�y� �f�n�P�A���\���ә��J͉`��v��dT
n�ۨ����A���析l&M-CE
cNd�k��0!��|X�d	'	�v��O�*�lB���B�@�&���o� �R�8*n
�$��1�T>��ȻԤ��
_Oʦ�YX��TKm�;���m�#�`��\6[ZZ�k�$���"A@X���^��x\��7��y��3�9c�B*�B��@ (�y% Ipp�E(>����D�p̰/۶m�>^�b��4Y�A�R%a	��*�j�8
C9I�$�Ů��N�v��D!��+��=ӧM/�ÐK�B�2��`�4�̗r�����8��
�V*p��$�`F4�2���W��1IC��پV�{��\_ ��[���4��>�U9OS���	y�b���z�ŗ\���c�0�T*aU-%�\�pVbb��/:���顾�]�!g1�25��t��TJ�tk2����"w&�H�&n�ý$����
��,�]���	%B1���b�s	��`����к�P}}E��ACr˒#�(�M��_�{�&�`(�G���t��9>���,lf
�Zer1��m*��n1��ipY��3�$�ZR��-B���+�U�'�)�J5�f���w���騣V�Y�fd,J;�����%5�?�#^'��#O�C�?�Ǟz<NY�kf�$�6�j*n��F�
/�$DZ�d��R�:���t��٨����.�˰�H;,6I5��l�u����ծ�N�\=�X{3��N�Ҡ'�xݐ��G���QUU��>k��c�(�zB��K6�&f����حv��I(H�v�eS�eRZ�R%({}
����B� U�֚n�4'����xx�F���41��v\�b%bs%�y������͍�%}\/���XQKtL��ŷ�sѮs��i��*�U(���,�"D�N.�����Y�t*�(�j!��d��cw9��Ll|4�M;Ñ��� �=����9#�-�|�J�Փ�g�Ο�M?��=�߽�F9vmY��;4x������N��������p���#:J�V)S�g��ŋ-w�Ue�ݦ���H"$�<>6^��b�l��oMu%�ۏ��|�g�rQo��A�%���w6�gW�1q�`ǰI��y)]/�pQ؟����9��y���>��׿.���~.1��� ��U��8<��ϓFYa���,�C��rE���F
ۡ��zټ��`q���T3hz:�\� q����g��8��T`{�G����̙39� $�)0��0���G�F�{��$�]7^<�4lkh��l:P�Ч���%P�X.��TZ<0P�E����$���0	5���܂uI�09̞K[ib���s�:[c<��k6$a�����o�Ju1ŋ��p�Aմx-[��)OP�Q�4adKBP�0�#L..P�_! �t��5TAc�r<A�������p/��ysg�}�� ?���&;W�LQ���mQ���~���l��������R�R��|"�����։h~�F�555<J�`����xY����i�iY��Ƣ8/�_=b"�aѼN�����I*�Ô�Pct9]+-�2�c�W,��y��c�=���(��%�R<�Z�spL�X�"�JJa:��>/���6{y#ʒB���H��V�䕩��K�
\����*��-1�nl1�o'��E�[�@�bB O��D�=qW��(��?�\����_�xn�>}�'��5��&��Q�J!��	˾}=m���O"�P���R�nŊ㰐��>:����|��}ht8,����TU��3&+!�) hV�p�
��3P��|�Xpڜ��\ �Z6�]�n
WTe��}m�q�x��,iw�=8�t�L������e����[�"e���ꐬx��*PS;U�+(�
o��-��]m�?���-4e�d�枞ލ7��`�˗/߿'U�h�cH�-;�0r�L��r��ץs����6w����l�1�K��ف1$�hV��"�G��R+%Q \��E�޸b?䯙?w~߁�(MyV��6o�H���7-\��Ԟ7o^kcMt`�W�����I�"���7�K0U+u�TЈ�T��,pr��ZTu���Vj�D��"��:0D�����i��g�}����ܯ|��-�O7����fP����~�sD�(�2G��S� �ev��_�r��wXY���}����g��z����p�qY�TE"�D�U�y=�xL���L�`��W&�c��5�\#���L���"D���$�&���~^�h��n%��383~����,��$�̙SU]�Mh쫕���ŀʨ|��%cԤ!`����^J�n��p��<�T����+X6dM(PE�w���BwC�
g������*��I�,j2m�f��jE�S��$��ڠ�֚(KI��p0#'�$؆`�c�����r;���]�%S��eW	����|���R*�-9/�3i�F�b#��Ջ�,�i�E�i]���B�g��f�bIy�I�U9�>�a��w,����R<`e8�8<ܰb�Y`~q�
�Yg��ԓ�eDG5(oTZ><1�2�!H֋�:�_��âsy�t�^�C�-�'�PAΔt�G�P�gQ$�ߧR�]Q�u�ǑN�T�*�*�ҍ�g�r�z�,u�PQ1��2��v�ԑH�/r�-K�������ܛ Y�^eb����^K��U�wIj$,��H�#1�M�8� � #	#CL�`��k0�D���1 �q(�E2<[CkW��ޫ��֬��|�����wν���T�Z0�"�������/g��w4ͳ�dk#�;Y�LsrC��I����Q��%>�c�(��BO������߫���5]&���K���B��Rd�)IT���p�u��Mٱ�U���]�)��<\)���b��O���^�=����d2��U����!�:���4*Nk�w�=�fz�V���b~nq=�|˛ϔ�4�7�+a9��$�7=��&&S4�� �9-�J��c�����ðأ�x/h F��]O0��;���"b��x�	�����1�|��=|�����7�V����[��VZ�4���� "�A��ouI���.�OQ�%:D�B�WN�E�����;Z´�<Wn���GΟ����f&6͟J���i�R�l<9l//.�1����=tF�����[k�֖WΞA*��*i�T���4�30v�
C��k�S �h\?��zUP�Dwv��0F�N�8c�f�BdQ���2�r]YY��������4'	��3<v��d0���|�[�Ο/�,'��n��^��E�x�.V�"ۃy˴!���j�/��@�x^~	U�8s]�!|�+��|�����avk�����d��=���/<X%2�'�-�ئ�x�h���?���sg;�N��5�$-?g�8!0����ӤCg��=����Pۗ/���`/&�&���z��C�uRE�D�γq��Y:6�iv���7�?%����������=O�?��+����W�r�=��>����IQ{�8:Dh�%V����7�>X��^gΞ��~ꧾ�����9|����gΦ���I˴_�t	�ݮ�=������XJ�N|1�9N(Rx��f��>ȡ��4�4��&Ma{�z�B-G_M�/T��{�7^�~�_�����c˨l���={18l�X^�o�C��%��q�P��x���pѠ�q�e[=)+Lr���̸�n��E-A��Y�
����ҟP��$U/��;;{l�d	5##�枮+�lBZ�7�}_��>�<��D�דˍ���B)'%�-�=2�dn��(\F�y�]��)h��Ɋ\>�3ҟӦ��g>CK�����N�2�u`�ٴ��c쨙�w�ֳ�˟7-T�a`?�}Iz{7u�#"s"��6 �iA����O�,�l�[{��ɪ"d.���\�d,S�<�����u���*��y�N�)���rĔɫ�Kעjo��ɞ�0�@�%T#O�[6V�p	FF���<�'3H\Ob�Y'���5����;]���$���Jݹ�_:��m[�=a���Xnd��-w�\���(?�+ׯ�<a��w�vS�L�N���Kԙ*N�K��ƨW�@�U.o-����%	H�����oP�c��C#G\"a߬�/t�pw�DHw���%'�N�@͛L����v.���/�"��1����<8�`qC�u�Q�Q贺�����{�[���'9�a�-%�MUs�	b�B:���g�#fr��1���Q}}OJK�������_"������^~y��^���3� D`��Z�&U�Ԩ�}U��7��������,�^|�N�y�Z_�]��V�-4��\��[���$�Ԓ�F��(u�)����C/%�?��}K��A��^��z�I�_�|y}}u�s+V�,yi�-��7HZmn"�p�̙���_��Wh�؎���mAh+ �4��+�؈�({$�JX�o�1]��� 3�A9F(�E�B�2��mN���9ќU�HI���H/���O���	�[� Ӓ]��\�^Py�5�x�_�2y&dY�!���h>�r���4��H~��2�\�X�����VFH~?�x�N]�;���ʢ ���b�GO�鉓����~��ŋ�B�����<��S��+�B��\�NX�Z��ڜ�y1�x8�ݜc�E�z�J�K��ޘ\��%�>辭I�zP���^"������N��h�Ҏ��K�>��&�ɠ<?�lJC�Ñ�����#�Yr9[)R��0�*��"B���ne�E�7<��\��+����;s4���W��Γq���>�mP컳7�*M�.��x`L4 8P-�Cf��`��^�{(�|��"�͸$��Enw:���-p�֗�n*ϧ����z'ǝU��-����v=g�^'iq9~�[�k]�*�6w�7�
:�Zz��u���`�����aB��-��6	Ǥ��`���ɸp��ށ���Q��o��R�}yA]�GbA�D���S�����\������gq*��v��I�@�>�Ϗ�7o�[^^t01Z1�q}m櫁8 ������G� ���}1��]�;]�vhu�?�ҥK$5۝���h~���ic8�0M�!�I�אK���L�����x�x�K��Cf�����< (�\��)�h���{��N���f�"�x��MY�o�{��}���ȏ�o���_�G Qv��r���~B�?'�����G�Q_�0�66L�e:`:�R�cE�پp��h,��*y�*T���r.�hkk���' �̿��>���>��O��$j�.U #�B�xk���j�Y���"�Q�wZ�׭��)U{*�m.��Eω;K�׿V6���=�Z�3�Zn�R��|�Rx&R�NR^@�g�֚ԉ�|�b�rZYY�����2��>����󣪶	l C�TI(�ǲɮ̬��|�2'KJ^��
ʉ�:T��L! ]�E�Ұi��U��l(,>}Zr�!e��2ZF)��jc揳"@�̝�y��
���V@�t1hlAJ���q�ćz�
x���H�D��3.\���QZ�_��_���gy����>�+Ș������;�d���Պ3C�u��zљN���[uܙd9�ب��l��M�����\&��?�������"�)a����q�RH�Ġ���ں���T���$�Q��;�0�e��W�V�Dbl�>�4�| K� �*��B|ex��m���#�� �
.s���.�W�_nEUgK-�\53�z^�׷ᇦ�o��qڿ��}������_l�����I�p)
É�I�U�Q=��H�)A�)V4�5\_g(q��0��9z�q��aW�
���[�sj�rZh�P��c������]g6����^�-dO...Jd��U`#Μ9)��˔�`���_i���y��Y`��&x��{"�UhOژ�h���~�:u*I�/|�B�j�( rq̧���~��Y%�YG�9;6��������G��+��
�^Ғg{{���|M���+t7i�Gf�9TDW�޴x~7�e���@3�O�{����K}�;b�94�����K(g�Ū3G� ���a���r������n�l�����V�R�$f��0�gsy
�wcz�L�
2�o���W�uD����QtT��[��t�90`��b_-#��Fz�A���Y��M�����}4���Օj�P��;�:��� �~�d�2�I)Sׁ�J��x�3��"m��fK �)/?/�גY�EC�^i�B;.��-M��p�s@g�t++�{6�Q�'y�,Gf?�g�����"�� ���ӎZK��4F��9����)iE����/�7�裏>��{��������mE��;%��_��_%�L���K�K���԰���X�o�!t�12�Z��xA[���?��'=�4��msn���]ބh�ξ��m��d�e:!�{�����\O�KxK�ݝm@ǈ���d�q�|�����p�Y��n�M>��%y���q;�YV��#�B�$��Jz_�������^{�Ϫ�f3�"1׋�dƖ H}��9SҤ�҄C�͙h��#�4��ƭ� ���Ћ�X�ke�7OX�Ƽ�d��4_�R,I�/t=N�ҡ��x$'G<I#��Rr�sv��j.`%��}A��
��x�XV��aq �xJ?Om.+W~�:�N@F�J�R��T-�TN��q>��O'�R_G>-_��ԏr136��!�ې����8jx:㔜:���9w19g��ݒ�����{�O'�#+���_�:y.?y�ڗn�Å�hq	1�N��1f��q�<�}��9�s��n�ըDT�k�6��Ѯ��}����b�"���>w@'���,��),#(_ɒ�׺�qc$G��削z��}z�%��¤n��H�
�7fq���j��µ�S��f,\�뫮�`��y��o�`p{-ON�8��VH�!��s0&ŕ����\p��{`��ȹ�J��(@-4?���S�J�<Aѵ�*���{����Q�d��Ih}��O9&}���=�r{pK��J��f�|�n^M_���ׯ�S�z�{�H����3������\��G*�Y�z�᳓��b�.ݸy��C�DɘJ�D2q���� >s������?���M�Dw�:B_ Xh�2{���Zܙ���մ��O#o�;�5�ȧ�,Vgm$�y�8��5/L[bx6����~}	 ���V����JW~_������JH��r��,p"ʾ�iKC]w��������6us'��ɛ97�T���1�J�^zC)����EF��%0E͐+����|�#��ַ�y�f�.A�R���Ơ/a苆��T��h�_�v� Ѱ�|�L�w�*ΫĐĦ)i-]gk�� E�$�s70l{P�� 4DY��8�P�!?`w�my!���Gxay�i+�n�@ݺh�siE�&�����R8
9N����e5���ƨh;K�������{0g�E��!�%'�I�Ǿ�PV�:Z2<�3q���f�.Z,K	n�_��m�yG�~�4W��J^�ǔ�y�D���'g�X+�4�M�[�FE₴8��y������_eM�x��J�r��R��T(5! wH&���(3��tN]UT��MP?�J�`L��g����ѽ����r�/�2�O$ߨo�7Q����W�R��T5:��>��	�h'|l0���Ѧ"Q ���n����k���,̣���^MϾQ�0�m8�
�L[IU����ܹsR���|�� �����
��hP����_l��r���p�p�ЇG#��&ܝv0��G�s{.P�C��W��<I��lI�7��Jά��mͶ ��{��i�N�:%������uk}+�z_��JZ�&����z��������E�rT�8���D�b���K�rQr&ު.Ji�X�D4q<�uqS�!�%hm4�L�[���T��x`����	h��D�y%s���(�fzAU@���D��Y
�@É2Y�^A����jU
�ϓӟ��������c���H,�b�dlؓƓ$�.�&���eY#ceU�zht)I��a�>r!��X�sBLc��jw:�lA�Zg�*p� ��/.�Q�P z�(>�.�aW����x���hσգ+Y�� ���7H��[��8�[_�^IA�qy[Y���|4:=Q��K ���Ev�r�3'\~l�q,����%���S�	��:�O�:M���FØ3m9l�4�͆�Ս!�	�n+� K��V)#
!<W�:���;m�#�ǥ��X�����S۶a������Pp�� 4��-I)�:G�� ���V���h�㉞$�J
lqy=�_I��o��O�f�y��~{�GO0;2��q���t���Y�e�>�]�3�ZE|9�~�r]L!Q��X+���v�O0�����*���w<V�����z\��k__2��֌��O{�l>4�[�na�#��Û�:���U�d81E��P�Hh���*�"��V�>��ru-��%�F�U�j�9bt�a��Vy�F��`�c�7��]0����"E��Y�H>��w=kS�*��=����|ɀ��VY>�t�V�+JXZ�4���d��E�CUͫg1���{�F-��߼�oCI�c�����1Ti?�9�/r��ܯ��p�����,��SW�p��v�o����#G�=�r��M���x��V�Z�=D�Ґ�I$8n�f/S�������x��w:JTn�q��m���୸h��1إ�*'톓܋[�Ə�H��t�{ k�N+
�Q9̒4��v�Bh
�F�b�m�{��2V��^�ϷhW*�D>&���`�D�˪�|��T�߰(��d����������W�dy�Z�۷G��Z�FR��e�_\jU�%Ew
�N�i��W��(+dR}��M�hN�ϨW���g?�Yŭ�Μ9u������5.���P���ss�PL9ix�D�[uO��্af�~.Q��S�P�<p#�Ľ��Ѓx�����Z�b��PŠ���&���2�SF���2���I;u^�o��������l=����t��\�[)���pM%ْ08��(u�a� Їi��zccC��]��=�O�LS���&�;	v�SK��qx�������l@�*igG��UՃ���T5�R4.:c..s]	x��]d�Ҝ�%*�>�7�1Q���lTl�t�Q`g�)t�bW��
��~:юT���v�bH��/	�Y(B�w�4'UVO<��Jy�`�'����U��o�o�No]�v�m���1���x�p��
�"m)�o�f.]|����S�A��T3�l���r��w�MW��������O�=��T�x����`�1��%����
n9�=D� ��]��(9(��4�MSm8r�y�a%{{���W&�!6��T�x;*R ���:^h�<4�\5� PQ6|��萔�r`�"��D4�g���@�j�Ҥ����M���3Ͽ�y�G��)������Dr���/��	��>8�_����Hv���rN�� �EZ�$O�m�P%]KKK�?���/���d�i�s�,�D��+�*�3�׍I�tׁq�P�	�UD�<o��GH�Gՠ(Q�$$�+�K��	[�ь��[h׽z�����j}�h>��6�L�����x*$�8%S�U�CU��uE��%K�rc/Nu(B�L����2,&�~w��dgh����~���w�Cᑇ�3��)94Ÿ$�n�ۢ�r=������4��lG��on\�ycL.��v��5���A�5��@�7��OJ'��s�Α������3��M����ۣa�?�����G.QP1�AE���uzg}�s��\��Zj�ہN��������x�7e$W�Q������"��C��6�p��M��萛��.0xm�о,թ���Ϥ�SY�F�d�/g�#��Z�K��x ��K �hZ9>G�����ڰ �v&*+=�ߢ�_lw{$f�$&'��םo����y�d�,/���`\U��h�w���G�x}}���s����\��W.>�`�%�g�K�J3;�Cl@�`Q���:,��3 %$��y�|����$Y�w�B!��L���kʑV�|Ğ�i�����8*�%7r���1aH�,��w��d��ݶ?��G{dշ|�E贵��:�X|��C��^��tU�������έ�q��N�a���t�ȝ�}A��e6S�}/�y���=R~O��Ok�~k�ԅ���ʥ$�#-F""IѸRE'uۋS���rB��G��G �1��a�k��N+O��΋%$��:���x4ͧ�-�_{fQ�ڥK����ן:s��4��# >��z勴[�<T4%-72흭Յ%z���h�聛�c�+�M���JG��c���Tr���fnN倦S{�>���u�̒ݠ:nl��|u~	������Ϋ��\��h<,�<�ڋKgVo��[�Ψ��b�Z�z��Nf�S�wE���I�(#�T���9�"�ߐ^z*E����ջ�!�:e���ݪ?�[����*��|Lv]���0�O��XlPх�FY�i�L�$mzˋ�"�Z����2���p&�y�P��D�#��+$�`Vĺ�O��}Ff��g2Ss6�/�v�/�|ie�����cK���w���Lw�D~�-Z���v��\xn\�q)#\�Y�r�*0$�F�M����Xc^�V��������6}���4��$�t�p��s�N��.H)���xD9A��/~�����cǎ�F��˽�4��@���Jg���F�qћO�����t4j;�p���)����d8̓4O:s<�{$��nYE^�pU&Qqh�w��Jr��Iaܰ�[S2I]�w��乗�v'KKh�zs-��dH��������#XYY� -�5�i����҄`_����qh����vi����/o@����oQw���s�'����涕���Jߊ���|�[OH0��?g�� �I�#�e�Z���6�n�2dC�d�	�ssS�"�V�.]B��X��jM�7RP���Y��L��.��f�0�և�Ye΀u�A�� ��+`?��ފ�Bc�N�@���������A��q��w�Rll�۾�!����!gރ"y�98��+����Q9�?��ЪD��1V�k~����C*��eEl��X$[[[��_�T�5ʁ�snnq�VVV����=���跴�w�-���Vnh�ʷ��������:��beu �e�-U�.W{���(�B|���J�C�k�c RE��G �,I%��{w�v�q*&#* �������*�=�*\�
�>�K�j�%�"����l~��
�H�6�u�7��b����}���J
W�t���rFB��9����.p q�3����.PU��^�����r4#�w�+�w4|��m�_�f���lT]�y�m  �¢*���,����_AA�� 	��@c���z�E��Ȫ�>G��;0�al^HMR��T;q�y�����o��>%��a)>b�����)���S�@J4��K7�����1����U�tIR�бB.N�T��d�ѧ#��,���3���%Q�x��/S�j��m�\p	B��&%���c�ďD�������$��M���`p�
����x^��g���8���F��h�+�%�,�%#��Լ�cr����(�L��F���?�I���6G�������t���Y&�Kz������VMi}��dUG�0�@������m����d���22f���>��מe)�je�!� ;G������<%1%&q>I:��Uq˝����"AP�����:�*_�Q|I�wZ�tY�9�R��B�	�����y��i4��zI��@���lR4��s&�-�KU��a�*ry�>��?�������/hV���d�)p��e�Ǩ�S�l��D�蹢�c*��q*b�:�\�4
�~�"���n�}������|嶲-|o;9YC��dB�Ҥ�^�ES]�06�0o<s}|*L�����z��M�3�16��aI4�tR"�,M��<��i����6��o�u�DS�ȃh���tBd28-�YB󽸜7����-rC�g+��a������|hqU2����\O�sc�K���0;;S��o��{�w��ձgh�^Bx���o!�Z΋��3��{v&yX��5Ye�Xe��H��t����LoU�8v5�j��m+n�͛/do0e��q/H*�;��lX8Rc����yIG�>A�����U�?�%I����{vcUu歩��|� ~���I�xC�>����n\�X%�A��Z*
�����Y��n�Z�Xfyjr�
�`����m���uXy�[>��3G������~3�v\+Z@��p(UN�� ]S����%I��p�����,��y]�:���9���X� �X����T��&R��>T�g�T�ͧ@5��Ǐg���J�|K����IS�̾쁜~�����#����h����a���`�4ꁔ*�������pGqH�|�)���D2:Kg���>"^ S&�dX�a"�-���1�jb�N��<y��ŋUXf����$YL�E:b.����q���о�Z��?Uݹܕ}�2PB&�m��fQ�O]�\��,-��@|M�pz��x���˰ݚe{��kǫ��<*�X�+�0 �<��� O�ܡ!#�f�%����4�2<�&���sbu*e���s�4��5���N����������~߻���o~�)Z��0#;L��UQ�-���4R�b�ajO��I�3���(wVS~�� U�x�;�q�b��T���QQEe@U��q�H�Or�jqD��i�B�F��O���
�dJ�"M%��/ng��j9b"���+V��XE?��=>5\j���&ۆ��B��i`:j�DJGه����P���[�T�ʺ*Ĕ,}��5��7��1�;߁%�����D��0�O~�s�vj��f�Ft$pp�el~���d��pG��@G'�I����_n�c#N������5v��u����zȕ0Y'���*^Mlo�����w�8��=p`W�����������9u��=����J��κ�N��f��#6��3J4p�#��[Ni%R��_����QB6���P�H�P]����%_��[�::~�[��Tǐ���!
�ia� �]�������U��l��C	N����[��kfwI_�^��V��/K���H쒽�AS�Y���������� d1�_rxvt��k뷻���v�e�x�$�h�|F���F:�nE�yZ"ڬ��!S�5"��x�,��)��2�h�E�������v���@o_=k�+,�)4��m�Z��YGZ��3���]��b����R�Ƕr<��2���6@���t��&a�2],�d�n�# 	 0ap��S[(�|t|�+^H��^�J*���Y|�������A+Z���n�`����T�U�[QqlJ�B,B��ׄB
'$�'=N�L�@�s~p2���kE�	au���	,�,�lU�"�k��܊S���(Dg�5���X��[��*�S'h�7�Nk��
�7ۥ�;9k�-�J��\��x4N'~;(���H���ݼ�՛;�x4�!z�:~�zP�1VP�?
��8��
�#�7�}k���wT�p�&�]���y�+���3?Z���).�g��R�d��RP���. �NU �{Q�q�a1�j���M])�� j���qg�3~���m^�|F�pʹ.}p8H��&�io�^3��a��aI��<]���Z�=���+��B:B}�ւ�<����>z��1`	���D�U*�s���x�����ߵK�$�>���4!��IGZ0jydm�ȡk�̀�񺠧��}}�[��nS��Z���:kC�H�޾S�|b�{,$j�2��^(<�ZR袡�X��,���^�����$w�ȩ{�D�2M�s�Bhb� =f��c@;Q���o꯵9)#�{(QjI�Z�C�d��6��;�����cJս�H��v;�g�{3Oam���v�رcgϞ��j��SkM�_��VM6b�:��Ha�'�/i��ycX���(!e�qp���ᖳ-uw��}��r�ؔ3�"���W_}�ԩS��9s�&�>#�zq��%QT��n�6�;��x���+u�Ue%�~��^���z���忛��L���
?A^���$�m��K6(�Ңn �+N�J�a��e�+ǙU_�M����FY�x�J���F �/{#�Ui���Yp�(1�U����!�Z��������?��U�7���3bW95���wO�G�]��cB��k�21y�L�H塪����{�A���C%w�����x��݈�O%��Ԭ{����Sx؜U�WW���,���h�����f�Iڑu���έ��h~VWW��s�.&Gʡ�� �D��$)��I�$K%�%�S����@寬����l��YY�m���Lyd��]Gb���~7�����7]y�^�����)��Hc�˪�veL�6MM�%�Ϣ�&��Jv����v���b�̏���#�=�5)֑7gwӗ�x�"��Z���ݭ�6�&t���M#Y^PE�9�T8Z}���6"��Ph��#��hY=��p�#��l�h#�Q��W~Vl�N�JR��пj���8�J����\wy�;=&g*�������(
X&������?+U|����/���=a�$�@�pn�ȷ���}`{�ԁY�ð�9�Y��P�Jf�B"ì8��ۊ���4��\�Åu�0NǪRQ�b���~�:��O<����/�|��� �1E����ʿ򁘳"�̤;�bK��?����7�B�9����&Ƽ�e���R��n>z�ʱ0��Fx�~��������X��*6��@4�ĠK+P�̤�!�������P7�[�g$�(/�V;
�KXb4������y�}oꀶ<��B$�H�սp�~Z��/��K��O'dumnn�]V\:Y��ma1hi���>�e���5��*����1�t�q�%S��<�п2�B>���*3�$�2'Lu:V]��Q��x�����y=A"c/�~��;n�E耊�ݫ-Ԓ��B ��/���b���ZGGO4Z�J�Y���G"��o&irss�]�{�~?��V�9#@�=x���x:��
�,�3�ڕ����a���
^x�pGs����������b�4��yv/*G��t�}�ӂ�\����qk� H��Sl�i�yK*�W���}�&g��7�����mÿ��뿭�:i�[��d<�)T�\!�a�7�)��[Q�6��s����J�r�d��J�jT�8��������>��D^��@y�M+�'�x<?�-��߫��0r9�N'$��߈�A_��@���ŉ�Q:�͆M\�Vf',%N�*�D����u���h�ϱY# �Z	b>἗Jn�aP�A��4(�EgA�,YE�5%w�H�mR��o�+���Kd�i�Do��hԣui�m��Pm���j'юx�����տ���J���wu����(Gr���M<���7]f���f���SO=�����::�������²�$s`dw�!r��I��{����$�ZULQ����4';(��*��M����A+h;�ؤ�g>�׷Z_�͏Y�I�䡇ZXX�����~��t�˗/߼ySj�Q�77�U*���8������c+B(��@��L El �b^�"��C����H#�X�tK SB,��Vh �]g�+��}���U���&*�_�1����/�/���&r@8���)F�ʷ��N���Pe��>O6���+?�?�����>�ֈ}�Pt]�*g(���?϶ؿ�����>Z��+�N{ib�+�
�ψ����_95�]q]��ri!����g�����M�rӮ2\<υDt4��M[Mv��}��v�h���Ŷ`#~��0��`����;}���6ˊ%3�z�"��T�;��4��0]gǛ�\;�Ƈg/�>lJ��n���uɣ�0 L��Xז8�&���ҹ��6k̬�)�C"_#���5bC[�ޅPai�F)��?�B���W,w�)��]� H�䦖���g�Jf��c�����=����?�u�O�a�������jP�k}�R��j��#�?���3	P[KW����vV��w�!E��'jww����'i�H�n�M#�׌{��g�z�Ο?��+W�\9vl���{�Q�k�6�s(�";@l���u��i��.z*4����'q��Xf�����:����|�;ޱ����o>�&��KB��WT%�҅�E�GS2�o�Z�����+ǖ2Z@�L�i+j�5����Qm��~�$rϓ	iz0��wM�o��o��mo�}�6M:y��6*`.��v6i$lB;��k���U����ӏǨ6��h)O\)���9��w�4O��		����lG�hp���u�!�? �O;�4��P!4O��)�{W`�ygq��;6��Tpc�6)�'�޹u����m�J�>h��M����B�#&*��.��<-��Q�������;���A�DV^9I�<A���f*�/�
���&#?-?eP�Ŕ� �+(dom6���G�?�����?���Y���L'4Gpk���#d)�*���ͽ�|-ieY��@D�J?�\��Gn��li1�4P�~����1��X�k�(�Ejx����Gd ^�Fmɰ�
=�Ǥy?���_.v67on,=0��F���C���ۧO��n�c
2@�����s�v�5/Ys%�����G�}"Pڐ$��h͓��a0�X\����񷐝�Τ��L���y�Y�����EL_'ú Jq�@��*{Rr�A3o} *�X, ���Ӵ,J���d7����k�
bՁ�9k����"w�����m9r.:ͳ��rF!m��`P.--x��`<ү�i��e���u�����}�9Z��
f�G��8�A��q��i@��a^��t����h� OM��jkf  ��IDAT$� �Y���Z��5]G�T�-G]i1�<�� �ϜZ`�o߾��u�t�d��C:ܤ*�،��a���6��tEV���S����c�Mn`�+T-�*��!"��yX�c�y�=��w�΍7��^�j�9R���w	�<ׅ��$^�m���L�nl�sKQ��6[}���v<Y��r��J8o��4)r��u�WI�@qE�[H��NS�A������ɓ(���D=�;Z}��;y�$��׮]�'��w.g���ǰ+�A��m�r��O>����/]�xqii�N��5��$���h<�F�ŏٻ�G�^���9|��{�@Zv;�v	݀���`�؊H����������_��6����r'�274$����1oI�q1���fk�[�n�}��7�����n�O�&��%�Z�5��qf��}�2�y�P�g�~)��1��,G	�I���W�nll�@��/(������!=�ړ��B�z�i��vj�<����4�h�C�UZ�|�HX����}�[>H4���r˦��ɗ,ZB��?%�"œR�%`~�Sэ� ��)&B�@�}�W���?��#]���� ��T�[�!+.���˭��ӿ�6ɔ���bY٬o-�@����.����g�T_������� �܎�X�_p$�(^�kf��j��� ���-a��Ґ4�$#�Ņ��Գ~��+Y�gd��)�.sPc_�P��J�1eM�]�s��FU��i@�����Z�w��xX�T�w���v���jB�t�:�xձT��)�"Z�w7GE�>&c^�a��[Y�RF \[�|�S��z�1���B�V���I���q=���u�]�Cy}���i_�.���Ӂ�j���í�[W�%�V��QI�H��%�;Ҁ]�����	S��Ld2���H�Yr߆�ٱ,��f�a絬@��I\��$`i�/.M��ڑ%�h�CWT7ސ�<ݽ���I�qAp���2��m�DdK�����.i_R��B ��(�F�s�{!
H��*�$q��m����nG�۞{w�J��3�2(_O�$�۽����+ׯ�ӳ|����� ������L뛓~O�d
M�U~�h}�_����hS�,P-ӽ��e2'�tR(��*껂���$�hõ0`3�3�=O@�b� ���V�a-u�V�H^�k?Hӓ��J��l����$�g�g.D��!�.γbn�KK,
>	*uڠM8�S�uYk���G�Gۗ����#]�L�[;�냭����N�;�
w&��%�IW+6�񐅣3d���2����;�����?���r�O�{N�"K�ƢIl��aG�25�wk�%}=9�^;{`��hrX�W�#��4>� ��ب-5b�ͣ�Mj�<E%���[B�8���ȶ�";�6|�2 �8��IT��MF��N��.��<��Dn���;��$C>�ӌ]G�8��x� �aX�W��C�B U��D��.Ψ��.�Hu��vhK�rTue��P]���g�`�*)���r�k'U:�{�޻L�M��H��S���'����\C��k�YV�}�,*�����t:�F�4�C��A�f9��p'7�H�mA��-�g�3s�����ݟ.��xQp�8�ε4���\���(U(VTJ�M���~�S��q�0�q�&����
�g���g9	(��[ةp��+��h`���>]�V���6�Q{Y�g3�޴2���T�YN�����1�Kg�Ĺ�!�^L?\�{;-ߛ�f#���re�g�Q������p�F��H��%ظ�:/ȡg!\�GH�ђv#g���D:��QV7Q��O�7�iy����(�g�Q�u�8�3�[g'���E��h>�x�F{�)=/�e�h��~�Or��g��quU��j/+Sv�%��ᢧ[��Z@};�/��K2�@�E�!�������Ξ=˝�=)�~�WH�d"6wLG�ߔ)g��Ad�!��h}�>B�`j��]�!pp�ph���I2�f�ƿ���| ]h��-�
h~�i��T�)��q�z6L&�!/��5��ʯ"᜹g�&����#�5�6�ՆS<��u��Z2�� SÛ��K�%�W5���<!���Ve��F.\C�\�oO�M�\��Ή5���U,�`q�W��:~S�>q �)4s�uL��Z{XA�s�7��^ɯ��Ԩ0\ݛ�t�;��/�/�>���\5�R�u��f�17�Y��B�O3cj�Z'��Kw�n87��+�+(�X�Ic,�!��9�dOb�9�ƴfǶ���%�ވ
ț�=o����F`�z�* [�}xZ�!}�<H�+�U�5ܲLU�*�Ü�9W1���z�o����qM���6ǉio0R���?�=�������f��S�&	�G�3��|J����!�0���3��P��&����D�66�$W����-�W!@.��c��8���S�
�"��j�4p0w����O��84�t�E(�r����Б����q0�ސ\�s���Ik��>�z�/P���Q�i����իW��������ߚ�G{5�� �M:��*�r.��ћ.��#R�gO�˱����п0l�x�Z><�Wu��;=ظ4��N�8v��)�1//�&�����������|f�+�HԒ�*:I��$#��iQ�N
���d�f]#�Ezϐ�������/ Ľ]M���E~� |x��T1�P^ܺu,A�g� �������Dyyr@�7�G)=y5����7���3���qB��C���k�Ɠ�>�d�'�=����I�Oe�$����B9"6=��������m����&H3�rB��+�B�l$h�W|>r��D��K��rlu8:����Lc�b�z+�i4ε���=A�k� ��'�(Э>�H.������1�0����NP�O��4I�)�?8%UN��Z`��/5��@��	�=��-����~ L���~������om�{c������Kr=I4�Z�@O%����Bt��N.�ϔLpT2ԙ�;c�7����r1�O9��V�-�[��k
��ƪ��l$�$�T�� ��՝���������ν+(�?I���B�@K�=�]��G6%����y��͜1K��_��O:�V���v�e��&<���ו�h�+�&G~��j__e|J�ˈ�{�d3�L��S.l�����x��V�P=��!�R�6��E�w#ȯ��*y0�{Y��d������|S1	#�{E��-!;�q���4����P�K�+�I3A�*���c?[W���V�Bh�>���{��8���s��Q>S&h�8P9P�Ŷ#v��|d@�[���SZ��0! /�L�;�]4���,ɷ��%���������gi��x"����m��4Ȏ�;�6�#��j���kh}I�7kOM]Q�0Xo{{����Ś���a��Ha4�Xp|�H��G�d�+����<&0�3|��g�%�]O8��;�J0����۷�{��{��H�&�G{���|�s��i2�dg�\�+:[��b�U&y]�\B(�W�YTZ_ռ�V�+D� ��f"
���?��V��~}�Ȓ�����7�cuA�/���%ݦc��۝�F����Tv֎o)U�H�1���iT�3g\)-�#���W��&����XM���A����U2��42��(E)�����Cq����ʈ�p�ʴ\է����ܑU>GU�4�Ɂ�w�bH��e<{`uL��� �^JҒ�d��U���p�_Q�v�ga��Ir*+$a�mA�jg�*��-�i�6���VVV�����JQ��K|hw�����a�����o�8=�fգVW'�ݗ��̒�\������Z��&�7���;�֟T u�������:F��G{@��룽��:ԺA�/@2�e�7`l8�`�X7�d��Nܽ�m����+BU=-��$�5@����W5�A�s�P6^8[�jz�,j���S^��kK� �c����J?e��R�鵓S۩��~&�=g����T�M_���TJ~\ X�@A��Z�]�bZ�)�zW�;&vlDa�N[
�����a�JS�*8Q��Q������ޖ�ӱ��;z0w��Rdu ���;�f&�/]��v{]�$�ղn�R���a]\\$_F"3�O'���MZ�������N��˿���{�t��<I2#s̙�B�J���]�$��jF��"G:�������S_�/:�<�I��ާ�?*O���� ��K�:K����Ė�
�zP듯�9�� c׊�MW�BTL�C�|���G�h�K�Sp=���3`d�my�s"oW6
=)i�g�y&M�,8��Nͺ#9'��H���Ӣ��v>�W� %���J�3�I������]��:�Y\4����8�pw�R��d�eŹAm }��.M���C�6�{�����doo�kO}=/\�3�v� �p�,88��Hj%K�Z�;d��&m�hN�i��ݲ�SD�=� � ^�jR�)�	[������|�i�R�^Ef�E[Q]OөO�4��BsײR���L�3��uN^�Èw�(]Zɔ\����^l��pj���6��.� C��Mv�4.���Ó���K1���ʫ&	���pW�0���R�s9f���W��؜���/--�ဎ�VuLN�%T1L��g�r��	8���B�_+��׬󼯙��0�H���Y�a�=��)U���! f/M��W�O
Y��,G��$;^���Z��)c�2ԩ���w>����� Vol�Kg��}�XGM9R����;����3v�%-�Sʹ���l�[� �ߘ��XN�E���*�*v�r}8�����cp8�$���n����:��W��}G5?K�#�*�%�)kN���do�UܮS�5-�f�R)�Sp�S�4/�4�7l�4-s�-ε|�E�q�p��厩
fr�\:��_$�%}ǘ&P\Cѕ֩f��Ђ ���Z�����/�=w'�w��>`���|��~�$�I��˲�U#����ܹs��`mm-/A��v�~{߃h�Ѐu�ы_~�e��dsH�ZI�Lc.;fk���FE:�FH �G���w�������^��+m$uq������}$������'>���������.K,O�Hf�4+�ǔ��<F�XɀZ�H�!�P�,���ʄ8�o�dđC4mCQ�S��os�4����%�L�?��?�я~����?s��(T]�Ë�����wd�p�@f�ñaIq���d�/~���)bm�^#3�K�%j�!����>͆��!�Rq_ z"�UѸ��:��SlX	�H�6�@F4Ò�"���ի�} � *�d���
X����k2At1��� C��&�D������ͤI�6b�bU
�K��[�3G_(��vY>��Ko�D哽�"�sĪ(^KV[!e�M#����I�v{�?����TFتb����P�d�;�u���ۖ��y8@%,�3�3d{�-��m��ɾ���f!�X���p��sيc)ʰ�^�:(�M�U�?_oJ[�~bly�%�'~��=3�J�K���*�����:�Ͳk�o7���P��~U�/������Sߕ�� NLȊNѯ�W.�@�L�m���Q��o��6�HQ���
�s��"��ز�Q�#w��j�D��Aۈ�'�u�đ;;η�k^R /��U��d�� �L?p%���Q�������c9��̀�Y�E�#w�Z_��/� U�t���@�ɨ���G�y�����o���O��o]��ʩ�gis�I�b�E�����jY�����*�*4�Ⱨ[Ý�,������镗^� ��8)��G�o��u��s7W�Q�������җ��{��`��?��#� ��=V�����0pN�X�޷��_~������	�{Ϝ��ڎ�L���h�;��򒖼�oZ:�u����^ var�B֬)M��D2}W���qf�z�Ή�rX�a�ۯ>�Z�������U!�i{��窘ʫ���?�����~�g�_��C�ə{ϡJr��2�.�s�֭$�>p�޼H�xz��=dE���`�%kI3��.�2
"�O��/�����4wa��c'�^KБFϹ~�������W{�����o�(��S�jo����7�i��7n���O�����߼�vkaqQ9�"ȞL������U�����4�n{i��M̤;ץI��g>�ͧ�uωSY:A-�dt
�{���mߡ�Y�y��� �JSh /@��x:���*�Z�N/����wVVVJ�H�R��r����������s����s'W���[ѱ�76�{ ��:=��!_��^��lD����}p6O7Fk{�w��I%�n�y��D�e�&���|����;!�;p�Q+I�����{�����fek~�:Q�u[�k�^=w�᝛�V��x��{�=��8~՞���+������w=���^��u��^��=���5�www����`d��;I��{{�xRNH9nm��w�'�:�=�V���vGn��ԋ��(�̐�hy�MQI	']7X�[��F�HZ�%n���ˣ�%���62���2�灟�Ct�n�s"8a;�`
i���OV��`�܊��q���#YŮ�#~�^x�}"�bD�BVэײĽu}���,)�I'4I�,F�j��|�|������� ��`'Uu�C���65ݖ���!d2fg
���"����7B(*a�vf)����j�jIy�*��;Qts���.nUfI�@F�A�U��}�N���=�-s����*�e��T��������k��(pc��\�>^�_}�Շ��رc�N�j%�[q�I�Q�
�c��3�j�H�q=��rU����e�-fa��t�D��	T�bz��sh;n�s�F�ҿ<�*vUocm���O�F$U�ʞ�����l;9�4	{#�\��nGK����D���	{����i�Ot'�g��N���;�z�y����7�������4���Ҹ �F��Z�|Q��(�l���2Y��9䔃�S<@�fiiIc$�Mg�>�ct�u������4Q 9��/]z�[��}���,/|��
�;��^��<�%���$_��En�c�=Fú|�2Ig��m�ZH)�B,�� iI�÷fNct%�{���7�����k�h�PCe�,��/ ~���ׯ_'����/�OL�ځ����w~����������w��������>غx�"Y4r�V$�N����0�Z蜩!����ܮ�*��zY�ȍ�w5����tѽ���<ɾ���ٟ���g���H�8XB~��D��ַ���g���G����O�����/�ғO>��7���ٳ�eifP-Y�i�H�3�fDZan�{(ڂK��4C�_��:b�ۙ�_moo��s]T�I]�tk�f���ҥK�������� � 3|�Eg�cV2ZS�>�!��o�Ư�Z]]\��6��d�(�� �1�3�{�����.����9�ߌ�ڐ�E��{�Wx�l ��<N���'�x��~��"JU
Q�C=4X�?��������|�_?I��~�	Z��Ѩ��8���'��r4�4^�q��Іy��:#��f9����E��x�f��JAJ,��������/ޟ�HҔ�����A��M�z�{�����o���."��\�pa��A'k��5�}g/S�����`@�zkgLO=��%QűnH�~��0 ��5[J�k<&�M�93U��g'���͛��a�U�H �!q��i�vǁ �U<	e������߮���F�>�A[��q��1J]�Z��!j�y"�G{ҠR��������U������<��j$'66��;��XN���;�{w~��h$෕�u��Z2��[4�v[�S��&d�?�ew�h��%�|Z��HK�MQ�~�D}7.�j�Q�Z�6�Ep�Rn0##�0&_y瀪�	��P�K���,ـ�D.%�'�#��hw�x�A.Fb{y^�0��| �\��h{��3,-/�u?9*>]��dݨ)x��Hb�g�������0�p�`���^4w$�I6k �ss�S�ץ��x�����.����O��u����d:��������Je��iG���iw����!{�1��2�TfQ���A���꼄���!�����O���O���؏���u#��Խ�O$8'O�}�����������?}�ӟ���������i�\��2��\w8A�<\�lL��B����dj�1�<7 �wm{��b䷋l����h{﹯~�#����=���� <��"�]�/�n2����p��?�s�Q~������=��?����~綾^"ݿ~c5�R����srkk�ʵki�|�x�wp+� iEH��I`�;�$�Ǥ���I�� ����I��嗾J��+_����x�nmo	��PEYQ�-�/l�n�B�������?���,�㓧N�9�� 6$�6F�V~NsS �!�Y��^\��'E��,1U�6�� �A	=$1F�����?�f4��	��,-e���������oٳ��V���.����ra�����������������~���c���[m���hJ>-c/pM8��?�o<�`�h0��:+�i �P��f �~��i���k�@�������lݤfi�������>�>����v���ގ��R(Ak���~���e��~a{�|�;ߩ�1�&\f2��2X]�u�N7��{�`L���p}s ��E��P��bP��"_�N���+�U�u��N�����=T0&a��W^�Lf�t4�����No�o>O"&��t����d������Fӿ�e��. �n̯��5 }�+>cW�iv�&>���|�>@A�O:� t;>��i�i�Ȩ-��s���W_����}���=���no��V�.LBF��Zdy�č���WkYa4c
dÙQ-�Evs	����=�!�&U��\gR0"��'����=(~M{'t�`sgyy9h7M]�,.�7��dDJ6
[q얆L�EEZ��lN_���T���jѾMX�W=�}݈(w�����"7�B�9� 8$qZĝ~k:�';I1��V���j'�����h��ߧ"3df������5&#��@3`f�%���c�y���\��(��B���[XY��$W�Vw}7�:��N�,�`�'�gԯ�������&뎎�.���r��3eA7��O��׋�+E�T�)~Ʋ�(������W�i�N?hX:�����Er���[k�c>�D3)V�)6���yG�/kBU]s�ȵ��`0�����n�>w�FZwߗe�N�N"�D;�u�+�R�����,5`�S�cB]��e�/���k�0=*�-��$��ޤ�=u���&�O�4'/g}c�d�?��w��]s=����jd�`�{��,���o�Lc���/��O����;���_��;����[�d$�L�{>70��A��W�}���<a�KX
��#=�=���W��>���~��!��������#@#�w��tl���z�Ξ=���������7��M���s�~��I�~����gΜ���@^}�`#'�|qiN�#�$��N�d\����i}AO��occ��'�|����گ������t�R��D��t��@��\A.�p�̉_�L�O�������>��s�*�I5$�ab�a).����02��܄�X��Bĝ[ɜB-J��E������}��hz�"���v{<w��:�߇���~�߸x�����������'�������7}�[:K}l�Y���o�����3�`E1��-���ڝk�x�AM�n�ޑCH߾6 ����~����>{��'~����?xQ��#���ROp$44��'��Lu2Ϟ=��������.>r/�K}��y��m�oЊ?�fV	�̫��k[��q��*D$*�-���[]5��\�*[|Y�ؠ��ӑw��ߣ�>�H����@ڑݾ}����p����';�/�Y��﫪��>/%�lp�l����\����Ȍ#�J�qb!h._�q�SdCo\��-PJ���;��O_{��k;�h'(��쀑�we���{@��s�${�x����Y��M��Qt~w���$A{0�~��珑��1�~XY�[�q͋��M��t�(&�3�	J�a��g���� ���5��R'���������ֆ�NU�Sur��9L��Ğ<�8�� H0T�z��K#`?ED��Dr��&������*}�ڻ�g���}��=�k{N�S�k��z��k=�4<�n?�+����6�����"L$:x<�e֐��D}�	r���v��`�gaC����oa�BkJ�;�)�ě~����)�Z�����@������8���x �h��V���D�`����礽�02�z�]��A]��vB�Glf\x�	ẹT�$�����Ѷ�����#����+�l�(2o���3���꫚�C�s���B��vK[<��x�N��c��U�-*Pb�B�7����Ǚ=��3�{z�`e�\i��ó���:�Ad0�[���޼���~��W^yZ̶L��Z�/����&�J�W'�/*��9Us/Y�h���F�2::���t��޳`lb��'�]�t��w���S?$���:�lbU����K̝�Jwf�á�akצ39�+��u��^���c�<�;��f�R�����C�G�t
0\��E��̹n��Sb��bUʹZ��tɑH�3ÀFcT�+@���W<�ԋ�ͭ�n��>C̉����'.����n����Wu�R�h��b����`dd��w�sϽ��SO�����Ċ���/�U�醪m���hn�~M#���Й�5wl�8���/7�s��C�s�|2�E�\v�e�_����w��Pf�O	�bT1a3�g7�:cO�������Ϋ��9c��?���]�S\G� kZ%7�;|~���/��t�T6�c�Yf~�n�(MN�D�_���n+�*ҩP%5L��#
E)���5�5��ï����`����VS�㲭��Q)佚�ɤ�n������v�v�Ig�v����?�0m�6B�&|���(n	G�!o&�H�*�l�QT�.�Ԅ���f���{�)�E��^7T�\,��n˶$V���)�^��j�B���6�ZU��d
��gT�u�t{#ު��妦�~PUc�?e(�&<@�)� ���L��a.i�A�e�.6�`���m9$v�,p��|��J}��Dy��[�L/Ĳ\�����22�!��:e���^����-��G�-ˍ�V�m�L4��R�}'t{F�$v��8p
�B���m}Ҟ����d��Su��Q-��ּ��d�UeuV���5��軦�uc�*�-R���ƹ�,�ؽgW�n��My���y��ɴ�u�f�)�r�C���Y>���<83|���ڎ��~��'�r*pC���!�c��$�%%D��5�'B�#�yr���L�R"�h4�+j[;9X �`�������;�U��#&�s�
sq����	Lj�Y]�7%hw ԰�B��	D�Hj ���Ģ`�{v��-5*^��*0�<�-�R�/!�,��X��t�.�|>�`A��FI�
u#�cͽbf�ik�#�4[,2a��:,�O 0�>���i�>ť�:�K�UI��	�#r�@BmB�yl%��5g�����ڷo�ȓC����o���hH���'''�}��^xa�e�>�vX~y�<91Q��D�Pp��ٚJ�;p��_�l٣������/��%X�B</��H�5W9i�YOO���0�w��ضc���������>�赇�V]�dr�8�'?�y�ҁ�����<�?�b�qP��A[[��3�J� �l޼9���ڵk���١����~��c�=�⢠�����죏>���y��_x�g��F�ྲө�eްK���y���fQȲ#����g�}��)q�E�<��y晿?�8�E�Pd9�zcn��I	��`�"����j��ٳ'�/��h�F.[���>���]�e9�C5\q� 8�Z��@
9j�`' �4[�ծ�cc��Vkks�D��A��s�UW]�i�Ma�)���H�;�#䥡�p���|��z%x%	��
e2�h4��?ݿr�J�2�EM8�k�CQ�Fz��jF![�55AH0��C#/��r�g�ʁ櫮��#���OO�ʁx'�P�<��%��E���Gje@�ύ�󐈌���^b�z5�ى���T2���{�r�՟�贠G��%���{n�333I�h4ʏK1�'L<�}C�J�ԧ?��3>t��7�<96��$�:������M 
_g���)����r��˴x~>i(��3�i�<KãA�!2_`̤��
����*� ���Q�#c�oٲ�^����j�����0��}�6b��C���Q��U��<}��rׁqY=�t)�b���vQOa�J{c������;tWKK���>��۳g4&Wٜ���-֟�3������պ���+����94���y1�w]�w�޹cGj�3ъIKg�����]���`O*�V����b Q�%���(K�H������s����y4��n���K�ܵ�� ���L+ְ�U���w|b��'�>��c���/\��/����$�B���*�*��!f+�����͛���e�,���خ"K��<���<����� ����utt̪��������!���O��b
���s�iNs{챐p,|�#<�i�=��%`�o߾J���Ͽ�����_�v��_�$zY�2��칥��)����ݳ��������Yg~�߄�:b�
�"���.�r�1�Ret|r��]��-x��ѱ����K~�ᶅK�� ���ϖ�b'��(���=����s�9g����S�ͱf�k]N��%>5=�v�1GG#a콇z�@in@$��c<4$2�T�S��y�w��_H�膝-�k��wd�k����_�D�v6D�j�,�Q�Z�|.��A�C��Dt7�p�2�m�������ٴ魕�����s{�{�㎍��R�U�(��s�Y��0���jVq:�8�0`�x<�	��N�ѭ�vn۶mdx�SN��{�/X�p����ǧZ[�Jk75=Ay�T�� �S���Ÿ-�\���5NMMͩl���?��[ny���0��&�I^�c��a��ʥz�����]�/�ql��j���2nh;�)�`*��\�կ_v��_�$V��rH
�<�5��K����/�&�Sr���I&��.�Q+W�۳�ou-Zz�G{N?}��w>��c�.���u��/�Ԉ�D�w�6��)5.$���*:�5�:��
�	��fu�",�^�5���੧�q�-��IG����}ި�Ú	y3�I<eS<Z(V!Q��:�wc2u��_0�`��������?��c0���}�+K��K�*A��T���m� ~i��M?��� �4��A�%�����N�(_2�gM�\Q�[�z(�LRZ\(�
1�61-qf���D���纻�I\�Y�7^c6^T���:�PC/�LsM�?8�o�I&����ƺB؜-�6�:���y<���X�0��6���΀Au�N�>F1	��Ysi��5 ��JELf2T��S�����Jw��j���s����;Lq&j���gP�b��Tc��r�P�3M�`cc�<6gܪ��N��>4�{�)��C(���*��љ����mkV��b����*�z�"��j��4ś2�����ή����#�K�0�@DQ",f\���8:x7ۃ�,$�y�Ɯ�2x�:�%z ß�XLH�&m���#�KE;���K�rQ��mj�fz9���x	���y�j�@hY���gk/m�{#��1�Fq�0٘y��,�r�t|�ܾ�s2�?c�u��KqɊ�#�iqr�!�Z�BѸl� ����&�;��p��3��L���}�H�/9tȴnH.'ث�%J��F
Ȇܺ4�N���rU;h���=�-�1:�)F"�),��tp�&R�!��O(7ydt�P�,_�*���9�Lg���JN����	�+~>�?����סyl�RQ���?88U�?��0��`{��㎻�� �a'��xddd͚5p�_���yh��չ��m��=sz|�t���%K��塇~�'}x���]mt�_.Pr�Ⱥ�5���H���8���l��n�aŪ5s��R>4π���v��ݍK��/��?�Gdhh��[oݰa�Yg�%�K���+��ن�X�t�]w���>�o=����j�!�s~?����p�}8+��[�v�S6�:f��;^<�i!�{�4=3=1A1�'���?��?֭[w�i��.W�嬔�,���+����������H֮Y���~�W��թ����u���{K%��-x{�R�p�w�s�����SN��k���eiLNNAo���TJX������!@�����a`$̿��I��ۏO2����W���/}�Kw�}�w��S�0�PLI�\�=s%N5hden���������n���/���ޏ�D�0��_����RqW+�-���a6� ��<Qf&���f����|��~��;�x��Mo�#�w,�te��E�={nB��gɬ����uC���I�h�χ�1��U'���ou`�����V*S.�_����W_}���aCuuuqg�3G-��`br��c\R#���8�x���s�=N��#B�i������Y��	�s)/�!�SҁL湟�zvO��WI��cci<Q�Ƃ�MM����t�D�-kT�����Dk ���T4O�Yv�(Ys�o�|P6����'���W���^2�K-?c���drU�%�$��˜.���H�ǃ��l�2�V�1A-$���a}�@؋��3&>[�ݶ,f�Y���5��Y��_0\�槪�JI�&��v���x
,q�Az2�E�ʩH$Հ���Ֆ���U�������g�yxϦ�e�+�Cu��8$*���Ĝ/Xqk ����b����1>>�Ymo��-�*;"a?5X!�x��v��q΅`�GL��W�pɔ)�lH<���ѱg)A���q�T��f��{Fx޵�%q�r�ᣎ9QV�%<~���{����f5�d�9`��U��6���g��+V���N��׷�h�`�a�a�!��Ї�@�ڵ�����͛1�+W�ܴiӋ/��v�Zn��x���ʎ�D<	�ܱ�Z)}���?t��n�N?6@�Z��	Eb ���׻P�j���#����a����M�%�s�9����$�o<���_�
';�

2�[M�R^x�o~�/�˘q��Ed�*�WGd.�����i\�l�����OV���O����r���U�A�yj�Y�t�zζ��-۶�ڻ��˿�����QT�E��,���:�J��aM�j"Τ�1��}=��_��g/���c�?���t�����v���n���Ϗ��'����%�M�Gƺ������O���Ͽ��k�����IbшiP6S��Uj,T�G}������k�S�x��n۶�����tz�d�rKedt�����%1<<��hc��,�$�H$*�[S���?���p[n���3�<�ͤ��"��^���u=���}މ�	h�O~�^t�W���?�����LW|^/���í�<%4(�˩�RI0l7搊|y�F��������=.	��ݾR���Qtwf&���R,����*Ή�t��I��k��ڥ�p*���D��XP�ba,"�&�x�{x���<뾿n����G��7o��߉LU$�|���ƆL��B�:#4J��f�%�RD��7�鉡���ŋ_���|�K����X��邍j9
c��:�������S��r���� Y�U+���/`M����g~���'~�����ZKvcU�ZRXg9�l�]�kU�ǭ��Ӱ9��UK�=Z���jnIj�uG*��<��#lm	a赙�b��4źB��)JN����&����D�DM]��P�h���ԄO�ؖn�8Zۖ�b�|&U��4��)ϴ�cg5FRD�S�4��L�����������,���#�	�r,� B��3<j,:�Սo��D�d#�R�{E������a;&Ǫ~�^��9�׽r��񶶦��Agd>h�l�� �H;7�8x�
kA퓅g5��HIV��ӬU�է�X�5���So'G�º�W|���SR.]�.*���D骬j������_������t:膎����+k֬�B���N�hǉ����H��m+�������;M�������@"�?�
��c�!� w����Ä��?dupp������fs�T�)����L�B�&�Ia�p V)W���n`��+{Y�a���,1��%��1���Pt����y���P�sHƾ�8f?&1G�r'�-U�Z�SY��ۂ�kE"����bf��S�1��j��;��d�XF�U��;�����\1�������/^yݍ�<�P����H�F�	�P��R�$�l�Z�]5���;KF9�f���ӹ�֤���N@�:C~�S����V�ɲem�[��TI��]oS�.<��`����B�2��ǰ��(T���D쨚V��R��|N��_V�q@ph�����G������_�"�/��7�|� # ���'CFaYy�>`�w��K.��{��>:�$�H���>F��^{�ՖD�+�x���������'��霃����]t����;�����A]L�G:��%�?����u�]��e�ؙ�\2���0��o]�k"���ע�p�X���I��۟~��۶��;���
y�K�~�5��+ �0K����Q���<:�7����A�3�yŒ�gwg�<3=����`V�(����@Q�ӎ����	`:�u�7�1��C�������+������>��[oa��tw(�nd�M�d�� ���v�!��q�����l�W�\9��z����&p#� ��ܼv�*}�}׬Y��}����w�y���'.���e�XC&'q�D���y(��	��t.M�馛N<��k��f��y�--�2�e��-���Bbl���&�[?������-y��
o���#�b����U�<|=D�{7����n��֓�Y����#>=M�^V�`0(�(ڴw"�.��x=cɩ�.���w�}w����q��Iި�
���Yv.B֫F����];�t�����3�>��y,�-�͖g��d����f����^V��O����?�xŗ�;N?��X4T��XEe��:u3���������-[��>�%���p�M�1G���6E�sY��H����8�.�� n��X�����r�/X����)~z�ʇ��3îL�G)��ܴ���3ix�D��2�oa�W�34F<AU!�+��y��?K�H�`\cub��4�?/�����"�����0o�i��N������lO�Q�Ɲ�*�$pB���*�kㆂ����L#t�]���5�
�I�.���Ǻ���>lx�W�u��$T��T3Y���n,@��o*���8ۏ���֪��	]�`�z�H9��,�$�����
@�X����26��fR����>��QrR0��T��8q�QP@�����3��4���yY���&�2�LN���I�Z$�%�s��c.qx1�S�iʐ����ڜ.V���W1�b��g��;�y�x��IS����#!�X4�jeQ�Y��ϸy{�ek�\)w�Zq�~�F��l����%j���b���D�.*yh{��75�o��ξ����xJ��G��׿>���~�=��賰ySc\����ӹBx�K>7x<o2�"�|�gg�5~�L�^�l�<��A���kUֆ�"�}�P�)��I�w,��_��"�I,=4!;f��P'��D�}A�@��B���H�O�ϋ���yOU�.˖-[����9�drj�R�c^{����]{�\ƺ:�F4�5��z٠	�utv�t*�o��ՇG�[�`����B��G{b$:÷g�"o�GV�$�@E�B�aB���ہ�{�9�<,?�4�<��s�C�^~������?��s�>���z��������4�!� 4 (���}kR��|[kKGG��������k��fKι�T�z�B�o���ٶ��~|n�[��l;���|F�`��hT�z;�Zc:�Ӭ>���ׯ�������iQ�#���궡ȶo�����Ù��G�����χT���^1�ڙ�U��	"�Շ-�x�<�7�N�:==�>��d*]ʤȋ����ڕX��}�p��y�ֽ��m����P��w��w��������oE� Q.���Q����	W�$��Zctx�5k�y��_����g�y樣�Z�`�;gf�� �h��8�
��9�}�9�|ʩs2��TMi��x�z!��Ş���+W,~�?�v�mO�s�s�����}���a�7�E)�v'�e%S��c��F����e�P�ٽK����ɭ�}��7ݻy�ukݑ�(d*~7�t�d�0K)S�;�}l��o�R��%��l����t� ~��)2��ǣ�\��nX�V�UU�?�y���o+����G�~�7�v��
.��R�\�X��[�p�08Ľ�`��ڼ������я���Y�xqK{[�ta��m��|>�U���61���t(nMvɃ;��X0�1�%���j-��KZ,U���=o(DX�X�������oK��nݺɉ�<�h�c�;�1�[t��d��	X&m=o��)�Z+����~�H�6��3���
�j
%���5�E�y 3�����έEaJx[rh��s?�V�I�N��T�P�h.���R���`d�8��%*��U��r����.OK�Zs`l�`Z"���Nx{�ә�E�2P�T&S��VfJ��rיQ���Ӫ��RK�Ȍ��e�h�d���gp�ꔛO�@�J���蓓����씬"T����5�j0�sH㚻���Ǩ��On3��֮ˤK��n|mp޼y�`��Q�z���׌$͕��!8�W����`��e3d��a[NH����J�@s��b�^A�f#9m�jnI����'^�e��r�%+�q����%�{�w���%µ�S{��ɦ���nٍ|��%
͉Ud�huƪX�ȹ�A�!�X��O�)��I�3��GSb����׬j���<u��㥼
����@Ԭ
��F�
Ɉ�Bvjk��9����76a��M����?��믿��c�wg�F!3���t��R*˚�Y�]�:�_UP�rC�)���%���ul��-� �:5�0X֗� ��j��(V�f9$���UPt�M�h�#��}�`eC׃�&D���y�0��A���C���/|R�倴�O������vd�
L���B���� &x����Z��ţnݺu�� F���������׬zP�F�T�SSЧ^x���+cg¸y�Q��Χ;K�u��J��UXd�\u�U0�@'D
x����h�Y�;hnn��0Χ�yf�ƍ+�-��v�3�����^82�n��?{��>��#��#�# ��[6���cX��#1�\֮�:�o~�Z����?����E}ݽ��J	�Ω��u(�_���P_z���~{���׮=��������*�zt����مۍ����c--\x�嗟u����/~���ai��0�̈́�Ca�&#i�$i���Dh7ś�~�x��z�Z�d����-X�䏿�5t֒����y5+�ΰ��Y�E �?��O�V;��5Odc^:ܙ�tG]�Lx�1�d8<���� N/���}��Ȏ����lr�L8�/�袓N:i��@`1�b*�����ލ������W�^�N�|�����P�,Y�A�U�������'|��O�?^5��x9j"`�����w�$���x���Þ�]��M7}���O�������%@�AF�b�k���]��|�����#wD�c���XIQ}��������RO¥K�bEFFǁ���{�yw�q�/Dk~O��x�h~o7\�`���Z#�������jl4�/I�1�Z�����{^�LlKcJS�Ib�.�����F�ɾ��=�'w��_|�	�*dEt�Z���S�Bd�߬�o��?��<^	��䓏`$��K/<������'�����$2��n`���F�ܤ657O��̕!љ1��+n�)�$Q��z�jMEA�mƨW�X	��[��Q	�bE�0�T�ER����'�ܺ��#x_c�
�wO/]> ᇪݽ{7��1���b��糔���j�d#M�Ɣ8�,�f/�8[u������&��7f/5�f�+A����$����Fcs;��+�9O$"ccc�2E&�FҸ�e��(x.<�[o�Bw��E|� �e�ޒ���jg�8�{5��h�_�kτ�Cg@�կ�%
J,���+d��ղ��Q�I�f���ۍ�i�KP�2���,ZѴ%!`ϽD����,ã
���"4���-�X���|������fK8���35q�Q$g&����4�W,V�(�]��t@mVi��N�Hb`�t��I�0�E�.5."�+�N������M7~���L�Ox���v�ģ��5��o���~E�����P]�X��@�Hi� �cyg��Ê/_����>�J��3>���f������R��fz(��qۇ���7m?��^l���^{O��s�x��;��\o��P4��ՙ���p4!�����ʕ+!��QO˞]������՝�Y�����5˱�h񲅋(?��+�C&
���N��J�	bJ'�>p���k�&fQ�_���皣�c�x<z��'C'�;�G>�A�5�l*5a7����%X��^�8�Ku{�*�d,X���v��50r�D��c��<E�i���(���N�N=9=�9������*3�_���|�%�sݝ-B��t��i���7J��
{%�Rd�s��o��w��K|�cg2�XD�]��TX<���w���<�F���z71��\{��k_������_�y}�|ꢅ+��(#3a��kz&����cQ���(w�Z�E����}z��q������<��KV�b�`5'|.��K��3�?b���#���33�R3�g-���H^�H4��H0��R�����O=븣O|��'����{G�3o�Ǔ�b�W�Z������ka<;��N�*���w��LNM�r�����$⧟�A�R�����w��3G�p$rb���4�yC�|}��������/L|���8ceK0�*�r��7o�D'���h�����[��4w�?w}�)G\x�݁w�yf��ҳ,�p�&*������G��;���Q+[L[�D:�NNQ|F.	�޳*އASh�Xs8���4��+�uݍ�~�	8�}p���阿t�Oo�у���+����<����e����S�����}!��m����?��|��k^z���{�R)��.Jě(u��c���ZO�ao���9����i�g2�����dj�U�꒣��%�ib�
f-\��6����x��X9:��4K����"��$�	�M�L:P`"5p�k�òG�r@==���!'��6�K�С��i�,,O�e�i��A�nI�B�n9p&����SNL�Q��%��R+��5�q���:X�\=�.����Uݼ�����B��=!T�j�N'���\8a_�*ե�V�����d$���G�LO몒e�V��B�y@�e��Y�L��ؽ:<�:��߅|6J�ҰL%�rNL���G<��K,�s��`0lIΩX�k���l��o�O����wll��%WNQ�Ξ�%n�b��c�[�����ƒ�X�����s�K�h�m>�6�NM�^B0���F�b3#
��7)U�Pt(j�-�e�^t8�x��fdm;�6�^����j0f�$E)jZ+2:V����4>1!�h�P�$�����#�fx�Fc���2��L1ZϲDsXDYg���2ڹ)a��}i�M%LM���Rٞ��u�T����)>3>$m�TVΑ��y�t���0=Q�%_oo߾}��5�o��)��z�6�wW]�_?�����U����=�E���3�Ų^�+�r��J��r����a���E
H��զlێ\�� �� ^8D5��MNҁ)~�Vj�Q�J��@o�h���x$�u/$�[sx����?@��o^�P WkJD��c�i�a)W�������
���^F�m��'v>�,� �ix]Py�Vp�6m�t��k?�����;�٦�лp�?g��������XD����z���_}��L&�Qe�yn�9��Y�$�T��S?�.��¾�>�񨻽T;n0o�4�0b��#p�S���U��3t
��N:��x?$6e)�,-��m�'��MLL<���j>�o��[n�;��!U-YW
����p	���q	3	�	lx��W�[߅D�s�'��1$ߚƹ�p�[�y[�nœ�z�iGu��͛����-s).��z������n��xz*�a{G��w�����~�%.W3� �L��^^(PPq����>�ĢC��s��y����+����jf�
��ȦP�c�������G>�v����G���>�K��	nhCuX;��L������G��uhhś�׬�Z���{��կMNe`Z�⧭����
��Ģ��Ɗ\�����e�u�IK�~��VNP�æ����\�~I`�w��X�ş;�䏜��������M�6��+�:����G���j�̩�j�6[�L����a5y��.k����w����?�s~�1��ͅ��i��AL&�:f��K/ݰa��~~��׿ߴLΧ���l��'�
��)&�oA?0������/����
`�����@�S�Ʃg~|ɢ%����f���|�z��"��}�7��K� Q6�h���6��ɰ�.���MFc�u\_�ݦ�C��ab;Χ~)RX�2e����`�z=�s�{���Уq'XR,o��=�ȳ��?#���ۻ���$�Z��ׅ��sy���{ث5
�B>ϛp��T�`PW*�W�����'ڂ��j�7a�w�~���R���^Z�ߊݍ�ڲeK4�vuu�v�B����M7;�������#�"��T���N��sY�ml��i�o�\A7b�ģ<1�g\����ĕ�^3�ƚ��U0�;wo��z{��f�$�Hh�T�0Zx��Rbi�e<]<N��n�`%-��݋��57�K	���E��0:Q��W�N"ReN����Ғ���� ��&I����H����X,���SI*�R5)C�	�t�68��ڦH3��qh�ȿy�q\�g�����_����#�vB��3XS*����� ���O6xӖW���=�\X1�jD|�ڋCA���.���={1�h+��NY{����ާ~�awÉ���(4Xj��JQ���1�"?�g���	�b'X(�X�dIS��\)��1�E	�$��s^Wգj,����n>�=r��`q{nk��ك����f}ʿ)4xO��Z+R$������-[��M7���p>�3�#�x�+�E�):������_�Ϟ�ө[�>G��Q�����Í���~�������V�X��y�z�-ݰ8�)l9�����d&t`` �����((��)�ym������RwW�ա�C]��WPp�q͒��V�:����2g���O��$��V�7��o��n���S3Ŷ��R����$A�n�J3�ٻ+�M�r�J���I��M(��ި�Sӕr!�<=Y�W��\v}Ѣ��5�Ƃ�-�^iLI��/[d,�r���@����#ӣs�"兹�.I�5։ikO�Z�R��o����ޡ�����Z�E^��A�������^c�Y�:�7o^!3c�2;Oyߺ�n���u����[����l>x�qV�*9���9;6���h"���ݰx� ��뮻{R�f"���B�TG#�f+J�����i˗�����O��k_�b��]~�������W+��n-�d�)����ˁ�!(B�nkz���;�]q㩧������=q�'����ܗ�j���B�n�ZJ�&'�2B�yK����>q��ýC�+��ŋ/:�ҽ1��hS���t���u[im��-�K��Y��p8Qȥ�1����_���+R��}��as�J5�L���=�hb���ua��;�Z�Cg�p��'��_X<���|���+u����7o��T*�-���3�:�����(�WK�������|���/Z�s��
���i��]�_r�^�6o���e@�i.W���|�HTf�&�0κ"ۊ�X��2U՛��k�����U�G#NU��:��{]�;���z��d4�]۳���p�T=!7\bے-S��H��ba� �SXQ�!Ϥt�_���L2��փ��E&V��f��6E].���ڄ=���,U8,:���c-���drdpo	x.\�jBׂv�=ا���i�b�\�(�|i�H�ZO��qʃ�%v�(]�4�)�(��ָn�H����� Q�
kK�uH�re�R�y|r,�K��Zt9)
X�"��f�<{���H�Ñ�x�)_1�C��t��p�^sK�b���FCWU)���֜�)�Le�����x�e	�z��i���Yx5Z(j�.����\�(���E�y�#M!S����vAa�ިa���Ԍ>>9�hn����[޻7�=�����I��czM�e�+��G1��.3Z��9���F���0)�+Q�h[A�䪫�B��<�����J�����Ùˍ`�y��-�x�%����{���S�>wpђ��GL����352<�<~�0ƒd�R0홬f��j������w։+��p�KO��	���.��ĚV)&`��$�n��%gM�*R�S�T��~\��<���p�CT��_����\����y+��SSy���4��F���Qe,�`ߝ���B�  �k�O�>g���3�u��<u|a��������+�ٷo�54�����z��t�~����N::��#�C_�����bI�~������s�- { �u��K����BS���_f/F}@ ��� ��:@��S�(XlJ�u�V�裏>��O���<�W?�}����-Mt���r�G`�%�ܹK�*===���G��[�|������䟞.,�X�z5��yV���gaFM#^���N�ge5뵃��V����A<ӛo�	���vbT�'�iޜP�D�^�3�{ʨ�h��+e�#������Y�V�_�sϥ�y1��c���5��h�]A~>��"Q+2��r�ʀm�s�B��ּ�D�c��G>��o|�m�=�����2�
��p$����&���?���.8T t��6h*�h5��^�S_�B~͚5��s��O�w6��4�P�F�����333�:�qx�7uK�����o��k׮-O���l}�c�9��_���Z��N%I/ծ���d��I�uf�P֮]��ÿ1���,(
����5bVHΤ��3��߀���E[��w�¼��}�k_����^k��X��2�r��תT�.�q�x�)���g�?���n ���W��H8�.Eu����l�� <X&l7H���	����x������B��fRmG[��`�\s"���%�~������`V�yM�og:��J�8�+�)���9]>Ӏ�Ty� l\b�bɊl)��V���.0t�R�_Sp��m�%o���o����rXJY� ���Q���h�v�z�t!G�!DY�=�R���O�v.�-I�>�E1�'� `��FMv�C槖ɝ�Rvo�.���]�|9�^��rg�̻ZNB�u��pu]�Q����E���)x�%�=��=RٌEMo��[���۶m+�SX�%K��*f�z=-����ׅ�n��L]�Kg]�)�������	�t���-�xp�.�c4����x�DU��N3��J�0�Q*�kT-�Y�9����7������F���:::��uZ��.XT�Z$^B�ְ��pw���':��C����ۺ��s0��YaM�yⱷ:�v��Ȅa���<��5�[Q6 ��2g�|����N[2��<@�H�<�p,�t�0���:w��}�)�|�S����_P��}���Td�3�y�n�Q�[�k��y�_���=��o�o���z�io�8e�l??>��7�?1��ξ�N��y���I�1��i��Q��T��]�w��a��뼾{0��s>�73ۃ�]���9ڇ�C��l��������_x-tʺu����~o4ܸq��/�|����/\ ��=���^>��÷��#�շ�n9|��.�
���_~�g>)�d~|6+f3a��"i�N=(Yo�;�����<���T�ܿ,K�O�:��ƳO�lٺ{&9�0LѤ*ݨ�K��F����^+���l8���Pd�fxU�W�$z�W���\��;����~僗~C �#?L�)E∢JW]R,i�̌�;;y6�^�LO����a=m�7~�K_ym�؀�7���t�%���_-�O�Q��hW,l�{�$i-�L��$�E2JU���0H^ǼX��9��z�9�	�����������D��-��,���ON��%�ә),KK��<n8~P�����J�m��Z�'�/���=�O� ���#����ݦ���$�t�NN4�Ô�b��d�kz�Rթ�v��Ls�*�=QA���/�Э��.�л�����|��/~�����T�"�Ñh����⁖	+_�C1�YJ��n��[������BG�\�K�/��Wn���=n���h-A�y��<Mr�ZH��}�â�q�E�/;�1�k�X�]���7k�M�K>��Ϟ��,�Ec��'S�|o���oׯ�ت�ܿ{vA$�y\�j��k�`4D8#�h.M�)��Į���>z�:��Tj�#���^s8]�֟R7첮K��l�u��Fͺ�Q�d)^�ִ]q�4�C�U��SddF?�Y��~�>x��R%�z�����c��U��g8\����7,)���?����k�"��)zA��5���{���i�V�ƔhQ�^�ٷlyCfE8��>����dQh`��[э�S5,��0Y�ހ���)�F澖�m[�mӞ�o��i�&F���D3$a˖�@Q��gR;FBv�S��ko�k���h�ՠ��y�jI���11]
������}����R1c��%�V�-�W�ļ�8^/�Ն��3+9��L� �er';]v�
C�8N�`_'��zzt�s���qMM�Y�\�D��Eۤ��X�����{*��-���%c3;bޘ�e��0��e��Bex:����0�_&5��	�U�d��D�]Z�,�ܚp9��P��}^�{O�nZlE�9���x��--���F���Z��b!�ѱZ�U)W[D{��`�s����:`��i��`5q��Rl"����`y" ��h4�B�Ȳĩ��Js����4����øiAx˴f�Ir]S��/%�LGIr0EAhk����?jT�X``�R!_�Q�9��ڭQ�����N��]���{����+�R4���ք[r;D�Ҩ��A���ŶX8fXnh����}�.:���\2鰽��ͤ�j��ޔ#�h�I��L�Tcn�ig�d��h������O�z����]v�Q'�3?�\�B#{��J�h��2��)�8mj	W�������y=헟�w�q���s�H����&&]!��ڬ�T�S+4D�\�+V�/]j��35i��=��|�Nɧ `�x3f��h`���j�Z+q*Narr���K,+�����Վ�s{T���Ԋ�
�U�S�ښ�Q�-H�(1g�<Vᐐ9g�æ�	�s���V_`��3�x��l^V��y���y� �0)�x�p�o�c�Q� β}�F����7~�<��#�>��/ֹ�&�/��\�W_^۽o���_�9j��78�&�N'd�
?�D<�A}�t���wL�mK����<� �,? ���sK�[ߺ��g߸��K�O]sx�)ܷF�v���v�V��j�L>cL��;:��^\��]��s�M�J{�r�4��@/�.�>��o�>�Wf]�iT�j����=ޕ �)2b�H8�C,�ZK{�7j6\{�{W�H5�L�x0�*����S�8��%���^�:�:2y���/'��_y���#~)���6퀥Le2�)�(lsR�K�k,��'�ذ4�V%G�B9a�̸�ፈ�ǐ8	�� �W_}�/���n���#��y����*N�ļPè�d:�R���a�ߪ'�U'>�5�7��?�������tG{�̃e���tV��=j�T61���U1����8�����m���k���a�\rɒ�j0(��P*ͦ���YҞ={Z;�q�B!C�z�8/��ְ��_\�t)�a�H{g7!�[n���_�j�u)��0Hʔ��p�́uh$v�4Q�o�[ae�64��q��[}|�������7n>���}
B���P����^�D|�b!����-Cl!{N<�HH>�����?1ipC1���^�@��8].���)�Sk,(RJ�֯��u����!�#��=�J�b�Ni����7�|��7̋a��Bj��Q�����ʑ<�:�H
\I��������X`g�Y
�Z�����؁����^�	��egSss�9�+��Q��]�vQ�_@Þ�g0�d:�{�B1�L2Iխ�2e]�D1	M�˺UjW����&--��cXS�rNpT����{��]��h����C���Yg�Q�K�J����+���E�˗/']Gd�z����"B��M�P�P63�1ph	��j�����,G��-�s��M,y6��D`�����O��j���w�)ϥR����H���0*��1������k5��e���)IV,/U��T��LP���h�$P�N.������z��jej��Z��X,�ÂI��|�g�����c���+�.Z�?����e�޽�r�
�T���y�Á	��)SjA�^�vN�8���or�S$s��T�w���8L���ݔ��
c���L���+W�+�ԏ���l@��*c�<��͂�I]I!T�ݝ;w����yy8�W��45R���1p��#��`����c,��X}t�(ˏu�]�v�̀�v� F�q�1`�l����o�}堼�ѩ,��VJ����Ƿ�l>���~���6w:�N|I��\&��NSK�w����04H�D1��n�Ґu���{��k�*�hS����aұ&�����l��$V�er�� �<lQ;�7����G����߸�k�.J�&V�i1��/�sc[�?M$$�n�����*��tE��e��|3AQ�X�F����CSdӵ�əp \.T��i��Q����l��h��*��n���xá�?@��!���nK,]���?=��O���/]����O�)d�0E�kf�F �=���k�W��i?���@��7�bႉ�=��=�=NEͦ�m-�����)/�o~}S�3H�Ґ�26���%��O|/պ��i�V��"?\�ƃ###0���'�p�	'�w���{Xg�w)9^v��)m�ݻ�V��>@ٿ=� l�-������d�(��v�3�hZ6��j�VjXi�\��aMʅ�i�c������:���b��7����/��G/��ܐOu	�^UJu�%���z�#֮L��C��!?��%A�=�ZW���Q�_ڽp�¶N��zˍ7�pC&WX�v`d$�	��/h��uy�Fɬ����]PD��zU?��R&M�yVY7a�1{��w�����S�?��۶�y�і.LX<��5�K�E��7t�A	�L2I�=͉���)䲹B�qc�o�}	*f�JxH9���9�ӥHAAT�MlG�fȦȰ-�~ʻ��SX�%�$����mb�����t�Ƨ�]�|<ּ��yT�YY��nN�2�G�PZm�#c~k6��߿[U)�S�Z[b��[�u�*� a��b�����ղ%8���Ӕ��g���`��v2�� Jb��4��U<ezr���v�+��ҿH�f���Ք)62u����kuCٽk"��.9��&�c�!,��ݿ�7B�w�놞��l$�
���U�*�Y�������`_���TxOv�mxC�h���7��Z[{kwWW:�����%}��^h�j��jժݻKm���Z���_�zg��^��4(�����\(��t�h���M`�� ٘�(>�:��Q�>2-Ơ�8�� Γ�K�`Ȣ-Juxj@����.�&�����pl���Ctz܁Z](��>h2��Rh�I�#1����U�Z�"�˼�s�0پk'��y�m���FZ����lki
F��153�]v�%Q��m�(z�n�ޠ6
�*��-�/�s��_x�y�_�����[8�<�������n��}���j�#��7m��-X����.����~��͏d��#�j���3O��*���K�9��M�X�A "����6Z��AZx%<�,���&��"�/��}"��p�����j���3��";ג���<���>K���O:�
T��̋�!F���իW���qz)�:����f,�>�I��-X��������x�-����=�h�6mz��ǿwӏV�x��2�w�� ���R�����]��8�#q�R8�X��r�>��3Lvh$9�h���������+P)�cP�7�t�����>�1HT��H��-:���������0fI�������5�寫%Ĝ[�w(��pˢ�SQ�Y��"�pS�$ź�����U�{CAb8�Sĭ���D[�{�ڵ?��]����[n��}'�
��:�xF��� ��m����7D��gӽ����O����~y���������e����̽	�m�U&��{�g���Û�W�{5�U�`�.L��M�XJd�M[�-KaHD"���D����D�F��F68��'�*�����Mw���g�;�Zk�}�{5�lh���[�{�>���5~�[�f�{��a~�l2b�y��&�T1չ�~�(z�	b�M�b��bs����7>��c�����/���O	�R��H���=ܾC�t�v��}�������/>?7W?���'G*hդ�X�eX���>!��3���Y�=���p9���{� �A��_��_��?���������~����q�֑�Gw����I�d��)ho�?rZ��1uO=�=��'����u��K�./�=��cϱcǨ��G��I-��8�����L���7����5�$/I����"G771���|~����|¸�W�>�=Lb�Lq\G�[�S[Ժ	~�>.�a�8��Y�uΝ;�0^'�M��D=D�L���2ɒ��d�e3��
���D��8�[��g�-[[�ͭۖM ���q�*�a�����.����3Z��[ZH8� gD��՚s��ѥb:�B��!yծK;е#���HO���7��G*Qo�`�H�m9kk��_����ܱ���rr��q2C��$�	��jyI�z�%�sJ�J����b9�a����=���s�`�FB��>�Ƥ��0da���Ѳ����s�M	|�Aw �??�HU�e^���L�B]jC�X3�HXzl�f� |�l��E��3 �8�u'Cϴ��?蜉�A����
1Y�z[�KK��y�on�����WD������;�ԉyb�S�3%�gSB�!�5t�C=T�-�7ױK��aX�q��o����f�)$3�ڟ��]#u%u��S�b���'>��O~���|�#�WW����sgr�bU�'��������3����#++?���똟�8q�4f�.]�y��|���"Z�ǥ�L����[6�@Z��D��bc�-���x%�İ%�"���z�tQ6��Ǖ��pq!;�����?0SX��r]b����H@lq�%�g��ԩS�q0w�I譅�e���c�A��,�m�_��=Z_S`������\�V�Īsxd�����t�C�x��S�Z/	����4��p6���2��C	�є���Vĭ�2*�LU᧷��<�j�����_[�����~r��ؿ::�~���9�F6�9��۾z���������M�G�����[^�?y��`�挗����Ań�pT�Z�p����I��8 *:�L+��p�#	�A�"m$8�fu���GAw�j�n6�g��?�����x���w~�wO�?���}��&�j�i�w��=�$��^��|���ǍJe��Ϝ9�y��+ϿX���I�V�^��N�0Rk�mGg����9��uCݹu�t��~��ױ���ʤ��J�6V0��_������ʟ��a&+�گ�����̏�؏}��&�(;�6eMz�.$�-N$Აw_���������/��w��W���^tm���ˣ(�J�7�h{�Jn�ڮ53c���1ʻ[�=����˛�d>��7/mT:�~��O�
����������?������8{����kQ8�tf��L�Ktf�]���q���毿A���a���֍��������9�����`�j�t��S�X\>�Ͱ�R�<�p�Xp���d'�M�Y=�K��zy��ln��7۬�X[�ַ��������ܳ��?��>�`�:��y���v��[�W����,������v��n߾�uy��9����_�ҞݭՓ4؝�[��}������F�nڢ8��N50u4F3�:�%,^�b�nc��Q����A`Լڱ�è���=��rZ�yL����G�H���kG������������Q����j[�ZJ����y�{i{��8\�`��. ÉÐD�I�t;gDKn��T��}�*��ۯ1�b��6�,��N�柨����u#^^z��,�ō�;^݀du����]�q����Qmv7d`k�r�gOQI�n�J���dͯ����(� ]��'b�YF��x�7b��NsM��D���m;�ť|4Lw�.���S�7ַ7�Je��V}����C>RZ|�z����6��9Q����/,U}ϻ~���;V�qz�0�rF	�V�;.�I/D<�)�g��L��s"��|_Lw?�6��[Z�F�anv{�>p�q�aW��.eF���;�s����Fc��W_�����O4���[]#�y0̫���G[}�;���9XYi4�A8|e����[��F�%���tY~`��X��I8��w=�m��L���Us����/_��O��g��������C?:��ir���GN�L�h0%#��ygs���}���Y�rև6�޾�¸k'Q��,O�~�Fh��n0NڳUѻث�Y^��aG��ĺ��A��a8����IYhOQdB��9���.S�����9AI�Z���δ�<$s��y")s�����uX׀)���*_J�� �TQ�77'�^'2�b���V|AuAH�_A�
�՚%�t�Q+mۡ��ʨM2��rQ�g�ޔ�ǒ�:bO��+VWB/��_���|��I���av<��e|Kq�Z;q���6�^�+��W8�!�
�C��>�Ĝ�3g�x�y��X-x���m�x9��o���:��Z���e%FCZ/௒� �x`_b�\�x�~���g>�ş�����?��J�!"�Of������`�Aζ�:X
j��gI��2+uj����g?K�T��k��������?1�ػ�l���]�M�Gd��Z��KSTB&������7�>wi����}����S_��Wp*pe�H���������%D��W��,.{��
fUlgA8cYa/�l<X
�����և�\���3��goQ��Qm6�n޼Y7�ǎ�z7�}��Gy�'�'?�����_�HJp&濳�0���F��>p���_��_��O���O���� vv;ƌ�Aq��r��4%|����cQ��h��$��#�P!o��n������$�v����j8Ϟ=�v�P����������Rhڦ}T��L��0�<���,�,������R��?�ӕ
LĞD����{n���4c��Rr���C2=�RS}z�05KJ͎�N���@Q��W�`e�=�=��Cu��4[^^�����&�ϚC����#�`8����9C��X��X�dl{�ه6%Bp�Q2f1�K��I����8�	eU0̆P=6닰�ms;_jX��KǸ$��{��릢NB9FX�E$�Wj$�y��7L����\�@Q��x,�\j��#�[`��l�¥���8�=��ӯ�|b><��.
�����=��p�!xs�1�f{�QׂB1��'���̈́��>i䭊��Lep ��A+ռ�ۃ����Þ�%��W_!��_���w�	Ȑ�AO��82�^����H��g��lm]���z���D�p�pk�Q���f��/�R���j<3eG2]4�1W��#�lN�aƧ}�'kme{{��ӟ��G>�S����sW�ݺ}��7?C�[[�I��X�8xy0�nc8.ZB\q����C��Y�tE�q��KQR�j�%��R� ���I�u�P&�L��QLno�b99�$adcC�PQ��[��,�j���֏:'�4#���0&IH���nO@"x��'sI��N�٨�)l�8��'�p���-1r��[F���r��7u���T#�U�)�u�x�����\����$��$��9AY���+3��fFH��z<æ�L�\%�,ɢq/��ۮ�G�)Bufu	�_�Ԍ��Vլ]t	��w]K�j�V����]�o�j���6҃��_���6�Ԏu��[j��{O<�03_���xЬ�|Q���H�.�i�I?ʂѬ�&����t=�y���)8A'6�֜�7���~�ݺo�YubX��;�s����זN�T��f9�����OGy���c�� ��
�7gmu�~��yG�`����v5v�&����2N���n�꾍I��
�ԯ��Y�W �b�C�'�"��&`:�F�+~�S��*'ϝ?����Q=��3/���׾��������^�!W��A��Z��K�����9�ݵ�,��\]��Q�E4t���is�VhsE�^�9vR�^эE���r�̱�yO��F�QQNՌaJ�D�aKd1��/@���}蟪$�a�Q��?k��������?���?��<��0.^�L�k{aeqi~V�>��#���������`��؇�!������mϮ2M�Q�8yʁs�\�&�9'ȡ_����֧t3E��Isc����Q�u���1�w�pb�g�,��*���.<��������?�M׃��Ӂ?T�R_�`�=O},���_��q6���SKs����f:1������@��&��ѪP�1�5����� ���TC��dy�G��K1BeC獵c؆}�T���Wz����K+��,�S�m����Ǆ?]Z�l��{�>��71�aB؝Z>��(9�G$�L�?��S��:�D�G2TdT�;�Q��\g��6��l�0�$�n�R��Q�.��Ҽ�4?s��s�ַ!����S�y�z�ҥյi�77��PlF�Z�����.bf�� ތ�l�l��ΧsCjX@���n^+��Nw ��Øz�E�_�j�[ĕ1�.w���T�(���Μ>c(����A�����c�.]�uzq���V�:��<g�sffl�S��zs6N����5]�8qv�P���vf�*Q�R�!�ѾɃb>T��HOQ�x��`��ӱ�����ln���v{c���s�V��w����#�f����q.��`Ѡ���(q}�i���h6�px:��*q̥�:���/8*�q'�MO��j�0��J������$o֎��\�pgl�I�8072-(��k/;>�t���k7����ɿ�����}����k/�zmk�T����0HqV;���ެ���4`x��	F1aG�[i��c�!��<���ϟ?����bJ���G�B��ڠ�&*&8�h$��xRe`�ap�x?��H,�����߰�*�ssZT6l\jڱ�:��({���O�f���X�>� �H|��xI�����G����Mit-f��:����:�V�}>G�&`���b�jƩ8��f�&��%�Ԗ�Z"%"�8C�wJ�Y|}2ML:]�&5MF��}alxS�{�Q�
o��e�<��!�`�b�f盆J1���1B����o��r[�AT�@�y��W�����wL��U1N|���^��Dz*!W/�N��I�/��R�)��p�<��ss��$ Ŭ����`4�٥	T�߇��u��U<��l���J��3����<���b"*�t�8U^%FDn+c8d���q��K�ĸ>� U���i�~�:��S]z�a�8���	#㈒s�: �zk2�d�JHcܠ$���H@<�T��K6�C%Wr�a�R�m��5�E����aD�ވ��������o�P��
�V���paa�7~�7�N|����a�0�pb~�'~�Vs�7�{�|�0L+x�4�MY8.I�)�l�4����A�5=W S��$��(ɦq:dE�C����W�w�����+�3�෷�_��7��?�#?/'�	���K/b�9������o������j�mAKy�Ƿj�C�%�b�H�)�r��ͺD�ki�|7��uU,�R�<�غ�iQ�hZ��.]t<B4�Ϋ������Fp����K�'?�0��oQ]Cs�/>f��=\�c$�� ���8�e<z��J���]R������Su)[gyh�6q�(x1Į�OS�ۜ���#|�:�}{s{iyy�{����y.^�0~�s�G��(�:tX�C�X�R]LηyLeis.H1���BB�����2"�w��������`�p���+��"h�V��ʵkPc[��1L�ao���0)������*&[vBB�$�ڂ&I�[%�EW���K���$	�>~�isl����>��3���ruC�Da�{�u I3�m�IA�=�׿q�y��P��A��_si�5���-"2S�!T�@	��GJx��{��YjPm����9UR�V�V?~�xg�����ٯ|��~�����9������/�z��ǩ7S�����!/�ߔp��۷�DIH�Ņ���a�����&v����o�}�<�,0��yO�p����լ�D>ݻ� �L+SM�&)ju���թ61ӏ����M{0G8���Q��(xܞ�/V	��C=���� �jW�M����95��s"I5˄�$Hd����~d��_�]�cc�Ʊ��q�0�^����v��H<��+���NgJ0�pa$��`o{{<�ha��6�] ��K�Awa�jţS+��>��pW�?5猻g�.׭ܱ!�0�,sp
W��f۾���������˱�x��j6D�fj��w�����q��V����Lu��؀�]�i�k~��EZZ�S�N��]���lǔLJ�U���_i�D�:���M#'Qtjua�;��o���\9��[ԭ\�p�L,V��Ey]��,V�،������g���Xݭ�NK���q��҃5�$qK�?��Qea.HҪe4���L�bѶ/�6�<Ӄa0�9�e�F�@O	���N���G�G�2�֝^�c��ӻ��қQ0w��fU�;�eq5���벰o�I��O��#15���I&�A��Y���۔���l�`tS~�ݚ!���kq?�f���'�ZI��A���*�"�	1�YV}mi�����o\��+�U|��+��taAt;�z�R�U�7�][�W=��̨���h���q��N�q��q�:w+.d�^g�b/95�C|�Vfǫ�m'�^w�1��t��!�ygW�*>��l{#�BM����^�6W9��q���r��/^������ssG�,Q��
�
�^ǯdx`8:Mb��U0̢��}]�����G�Z��\[�R�K1�(g��p�\2�	���.�`q� ��*F�3|2<r4�փX�Ν�+�8�T�P:P���9��sG��|'t�_j�Z�d��y�������c����5:�/<x�� m��j�ĳv&}�I��iUC�.+�Xδ��ط#	�V�f��J�N�Z�yϓ����Z��+W�tz�)�����px!i�J\�4�1.aQ�Yn��d��mU�C����ٔ�僐9~ġm���ձe��Se�cf���=�n�pb#�?�D	��r���ݺy����Q�����O��4���Me�>�-w?�T�?��e�������YiÕ��ys�R�Mqm�!���̳��^��4t̃�o���ŋ_��y�ɳ����g���k[-HEHW�Ls�م�W_��]�~�<�GH���2�|T��/?�i��	�P��6|7˓�~oG��ce*�3�cש��DA�f��^jP���t� ���[����\9��?�������{�<���3[�`�ߺ}��M�����m�ƻ�W����x��)8׋�0�_���0�pf������?���"�w�ҡ�(I�s �N�<	E�-~��,)�2�y�-X��M�tB\�ܹs��ޛ>�	��w����k��'`��q��� r5.���)�
["�o�IE�!��n�(R\�wF� �&�E��?_����z
�#0SHBx��J�rW�_��C}bu���Ɣa���f��L!������:Q��ۜE��<Qw�%�숈���l�8���{1�#b�a�K8��` (�˦�`��+��~	�@��"��u����o�DZ�;Ө`ix[p"T����%��|���Θ)�lӊ�lb6�%�"0V�w�����'(����%e���o�{�7w(��Z{X(��M"�cu��F*��m�c-��b�a�G���8��� a[��Ql ��=g��KV"��D���c����N�o�X��A�ק����E���S��e3W��/�)N����$d�UM92��fE\|�~�C,V��Fa�f��+���j�#!+��4vA��	��o~�!�8>$Vb*�8P:��������\�a���ǥ��>dUI�&g�p�8�\X`�e;W��^�Q@�)8��NJ\6��N�h\���[k� ��D�Z�#:�ݢ,��W���1���r0�!��	�k��0��zK�R�1"�xV�sz��u �Ns՟]ZZ��~3&>����y��w�~nQ_�d>�Bk����~\�7s���8��&�O�?^��S�]r1=��b`��Tg��䡄�hO0=���b�Xs�V�q}�N�< ��->�)����4��wT��m�'(-L�~E�)a[e�\Oj�HGJ���j���\g!�~�����|�#��Y^�i�g�_q ��۷9
K��.P"��Į��R��	��H�*rk5�&q��T�aT�9���ܺu���x������"�$\�6T���(�����7���T�1y,5�x7�J#r��`�~�a�n��A��V�ް\���.�\����7����	�Ѡ�R�#���q����;��'&[>1*�#ϒ�� ��˿���ml�(pGN�~��P�qF���ƣ�b����j��ym��7�:�<u��誙;�"�='>AH���>m��G�����sU�VK���m�pql�,�dd'a�w�ˋW.X��A����p�v�5�h�ZpN�|�L���j6�v*J`N�p_4��s�0�
�l���+U!����/-�U��j^��<M�A�@%l^�p5jM�S[���V��^=��N�����7�3u��Q3>���lcc��|Vϵ��� �3A;��Y�Ā]M��]b�:��J0VOI��=]��AaW���Z5��qܵ�Jh�5�B[=W��N)��%�X{��S!]"���������` E?�l�v�
��_R��vbg��8�p��8%[{��]��i�D`���*�b<��{��z����Kfh��37-s����6�i[l��G9��<���6�8��lT���n���(�>f,d��q�G]y��3'�YʪL�4�*��g��7��U���!����ĥ�|W��:7�EU�s����C~�@L���*->�-��N�N�C�8�.��dйKM��,�`�)b�1�"3���U�M�k�n_�J��@���u�?9���7;�����U:ȵ�ǀ�e��c��%d��I�o�E��D*�i!��0�3?��L�]��" �đ��f�l���r y���/���;]�$>� �K�T~���6��{H�ECr�zR�/����o~���Q��KM�a��.T.����)���E�f�
� �B�%���x����pƫ�kg�Sj?7w��=uhY����m��wh��),�)C���(��SB��fА���7�NJ�&H	z5�,/�L+U8:�9���]c�����}�m:iD}�]����X��|���e�%m�0�͜BL*�g��#&L�$�@1�H��\���s����/�D�����q�EƦ��jQ����Refk��0}�+�_������|�C?x��;;ݛ����]>A�}8�i<y|����_��<)��=��ǁP��"8'(r��&4�8	� �8���#�����9^N��Ԟ����	z�1�v�A�t��՗߁��[�d��\_��8�D�Jv�ńY�} �NZ�KPB0�o���	/���z+-r��������KP�4O��{`X�#+��<�x��	����`� 0?�](Q��s��L��hx0}�r}��:����&�:z��k�]�����R��f�jv4����{=�Y4�������'O�Ĵ��f� �(�t��	+~*6��������UnI�0��!0B���^:u��h4�Wy����?�y6?M�f��tR*y1E.�?1��� �Т�����p�I?HA()"�YY9v�8܎��u�h�([�g_>Vኝxϱ�
�6	������!//��*~Ǵ҈b��
Y���ߺT\+zO��-�\���,E�|NF�[E��H	`E��	�.az9�$��ĥ�q�q��<�`/Mu~?�Т��Ah͵g��K8�d0��4��V��c�0�6�+ká����vvv�ʢ�
�I�L���'1�ǘ�˗׿��/�>��N�`Oz��P<�RӍ�����v��}6�?(ۧ��e��ox]�ord� �@p�����d���e��|�S_�]��#�ǎ�2��ЋD"���2����H�rSL�+NL��Bubb���?��/J?=Z�L�i��㸅Csss�hp�탞�)��w�����P��y%�iR�I�PxBg�Y�(K�4�ࠔF#e��P�������M�O���
f��(�7�a�?K�8��b���O����k;
�Q�k����u:f��+��H`a��W�x��/��kp�U!��t@0X�Mv�CtR:�2��P\X1ق��R�5٥r�˘���9D��J���g>�X���K�����?�p���&q���]Q����ݮ��/e �̮#:$�
��[$�e1+�2B��ِ������뇋���=^���s=iq���w��C�;�Ƃ�~ê�"���p1#r����<�ڸ���]�qolQ�XZ^`�V���IS�g%\1�[�JR� %�	�n�d��P*,�D�q�#����U��%#�m�d� 烝�&���&���ɵ��v�\_jZM'i�ɮ��^��3
h��9�2J�4�po�m�y���<}r�s�r�d��4+�b��M��u��Z��^�s���؞r+�0��A�۾���������A�s��${�Y�'���YʚiϘ�ݬV�z^����-}�
g)@���ؐ�8-߮�iN����m�ťv�5���P���s�sgO�z����κ��Xθ�p�U_v\�D�I�c[���z�ML�n���M+�F;7qB�cf��4��S&;I���W���ȝf�	����#YmrzP���6�Cg��=y[�{�EGb��Z�5
\��P+y��{Hۜ�Y�:�B�9'iTI)S�b�ik��:q�&|Tr,�p��t�[u���&K�+�KĽ3([1M|}�4%Z��O�A��Q�0$4�'-=��Z',4e�<�N)�Z�?�u�넩a{.vq�A ���`tp�'$T��j¦㻕�A��2P�f�Z�r��!�� ���z���'d���Gׯ���gX�ի�F�,�!��+R
;1���S�������LR3lL	���PL>�p�0�ӄr�Y�m��0�z�9�8?�,����t�ȳՉ���ck�*ѥ�̜�4�$컋�i�����s�)��Տ\�G85�e6��Ļ=T�R�6Ch9]�N�\5A�#,S�]WϺ�3�¶�e�� �5�xu��[0����֕Ş�lNe��x�C����ȁ�,I���G�TX��X�U����5CY�(��<G�R���8�u!���(�S"��̫�Y�r6M��!Vl��E���I:3�z�4��)� ouLa�<PP�(`�+�p���1��n�|p��Ψ����#b�Ξ~�w*�2`A�=M�/���#��)d�f��"O��X�(a�-\�x$�,�9|�k'�㷉�gy<r��僭LS# �M�u��������ͅc�}�y���7������=��NB�Y^5Q�����:�?�X��*Äĉ{�ԻQKj22ΨE�P�gd�s};\/<R^!�Ju�K\��R���軩ms��-�#�����%ͷT�o���3�Z_|2��c4�\��?nR`��		?V`�ԇ@��-��`�����<GE$�!b��� JL
�'��٭N�3���68� �H��I��)��c.5� _\�7,���������e�¹�«{�-BZ�"�E��bF�r.���͑#G l�a�Ӿ>����͵ܕ���+?��?=~�8&J�V��8z*�~M)��	Oȃg��Zu����U�Ii���a�5;+�܎��ʮj���u83;�(� ��ق�]�=��I��rˡ`�6<�O)�󏥇�I���*� �Puj�y�&�S=_V����OR�8�O�uTUM��^Jw_��8���$+&U^�#R4+��'c�C��J�:��QB��,�0���|�A����DI���0�A��)��NQU�('�9or}-��I��|8��`M��*a6�����~gg�z��͒��/:	��wG� ��e��OaS��ƽ`7~��ۖ���}���O>���pN%C�|����e�Z��Ĝ39}E���VD�ad��p�
��,
~oll`⍨�T�8&;ۗ%�&��/)R��p��3h�2��mE4Q~�ٙ�*DEO�H��b'�$q��_�2RJ�J��"��_�`�'�f�K���h�NwG��I �.?]V��\�����yG����6����
�l��`N]YO'��3%Z�(��lo&�$�K�ɫ�ꎙqְ���U ��䕍������h����^�րK���qgS4�x4r,�����[��X��U9�i�P�Y�6�P;NB�q�[� �T����M! d}q��Z%ИgJx�"[�4^__׌`����/���ȿ�xU� 52î���"%&$@���2KOZ�B�bwq�!��N	�GZNG���C��8�b��m6�w��ǆ7'iK)���!�	6�X��z�I,%�Dm���M9�w=r���0A6	g��� �u����P�����f9�Ӊ&๠��$��3����݃��;lxZ��T^9A������0�mm�� G��u��>aj�d&�dဒ'J�ռ����|w���G=pg��(��׬ר[��,����^|��}��*Lr)���L���Qp���������Ӕ&��0S�����S���F��ބ��à�l��3Q�9�t�0�S�-S�����v˫:۷��������|�xow>m�Q��}p��25�����qvv��0�ڔ����m���1�/&D~^F�%�C�sm�bθ"�P�R�!E�o�`%NU�~4�A_R���wGh�Gi�-��4��P�i�ډb�1�:x�z���&��)�2B)������m�))�F�Q�[�yj��q�� Qq�c�h�ϴ����oX+b��lOߗ9� �=� /?UT�>
��fkg��a��1���a�4\f�%�R�5�,p�Y)�+ �l�00��t�`���ئ�RK��}���o|���U��?9�x�tZ����N�d��0/|�0w##�i:��k)����y���L�R���S��b�0^��c���Il�G��.>��GA�%��L�bfC�� �{�p��S�έk;�C�"ۢ�bvQ��9�$�p.�Y�w��'��~Q��-Ѧ�E59���&�U���ݾ�	�A�ئ��ihW=N
���EfC�v�(CX%��iX�!��J�Cz�
?2�9㞱�6h�C��^�ͥ�fnZU�=�Z��d�=?
��cS�9��V-F\.�hS�rk��'6!S@��l��H�F�e��Ey6�YȳH�qY��`>wz�zޕ�L��h��w�~�9AB%$iV�P�jm�s[�70�3�Z��a	G��|�;��TO$/,F�X"r;���, �l���r%��wp�Y�3ץ�I�nh�K���	�T���c��(���s+��l�
�t8c��Z�*1E�[�V+MBX��Ĺ���~���#�Y*c)��	>)-�<����,��G�x᠖�Ҡ��v�1�Z����߻����P@��0Ui�V��w��/>�cQ��v�Ne�$o�@Q.�/�u�i���sԗ�p�W'9�(q<�~QP�R�vF$Ƌs%�-H"N����\�ڈ��ӛI�4��G����'����29� S��f^޻������JS�Ev��/�w����3gμ��tΞݽ~���r*��p���:/߂O����#�_WE��f\C!��qwզ��B�Ri�*n�f�>����R2	;w�l���|�0�Ϟ=�9�������gȕ\^d�˨��C)m�a�`V�R����`�͙��9�F��"�	���ʻ�S�	xB�2�M�~�\���!����b��^&_��/#����b)e��!s��)"H����ϖ�~5�.�(zt��e{�1��gSSw\ެ��s։�	�8U�-[�HL^��1�n��؋�y�V�����׷�x��8��Q�K<��V���8x���/����g��U*���;�6��(�,����Q�z|�2\��8��g���ZԎ�D��p�%�j$�1�s-�#&�)�X���P�7�
M�[Hh����0��;��@�bB��EP���}��w�忓G9B=�"�8���\�~j^P�v�Pb�|��3'�9���w�/=��KWmz�&oyv��aDǒ&E�E�O������m���J���v�.�X����d"ԊCa݌yi<�aK��0��$Z3�="�3�=���a����o$>�#>)=��B\QrJH��c��x=�i�(C��( �L�������I�S����� ��^��+��A��n6��2�I��ѧ6����(2q멒���*��v�0�p�OC9wѤ�\�/ox�z�7}`�wwwq�0/���8�?1�dR�|	r(���G4"Wu�[�j�����ĪU]r��Fs�k����R�Խ����ZmV� z��=q�����g����8l�+�΁���3�'}��k�T��ԃ�k���?$-3������������a�-�
�{�8s5�Z~��u�WTg�fھ:�ǋK����d�ܲ�^��z��7ԧ�:��W�W:��Bc=#�;P����/�I��\������V�l�v�!<끥����߿U����W.�������`��Z~��ټu�"g�RI�?��o���6N���l3s�0��n̪sW��7�������Q��Qx�+K��v-c��X�Yu����m�F�����kć��n]�y�o���G?��{7o���]8�7v:��=������=�`�漩\2�>����$ǝZ+����o��<�}Ӭ��EULݮ���<�r��$�qb��V�����Y�N�hk�9����&~�*O��A�*�ٰ�a�������o�xҾfC�Q��.�x���w2��p [�o��:v7$�T3jL�f�5c~98�V�ъY��.�[B�'�u�֭������'��Q/�탹x*U�pȿ�`����/3�x���2F��wJ�j��I��N���	���w�c��4�ɑ�3����-��8v�ɏ�^�m���f�^�2�F���ރN�5K�)����tv����2�h���Q`B�/IvBh�{C��C�w�m7��|ط-;��"\H��ԯI�d�`�L�mr>U���f`�%�a�<#ZP膙�X�+K�(�G�奅g��"��n��`\����-��ۭ8�ݡ�7+�m�-{;�j�9��X��*>1���RT�q�$��71d��&�}AΛ�}V����'�Z�ێ���%z���^>����6����0u1oUמR�����6ׇ�����p~ʏ/e�*խ��y�V�������
,'8�q�,x���t}��0���^���d�t�%,��9���82!��0ra`<U���V!ivsT�P�V�L��p���^Â�0"j��,���w��IMK1R?����Q�N٭��0���lΌI��*c�����-c�:��1�ԧ����+�~#]��3�ۻ��������ʉw�ɟ����"�ͽ;d�n��)��66	?Ħ��t�кw+�<'�q8�dg�[%2Xbӣ�@�����1g��������#�5�,W��˅�>z�(�?LiӅ�!N�|_�,1��Zx��4�0ϹWؗ&s۸w5���燤�%J*.���?/U �e��i�^�Ø�p�B���7}0�2�N3���6[�cǤEXI �����^{�_�����̴�j�Ό�yb�d�K�C�8�X*�|�.������a�P�:�cp�'N|�sK��{ϕvPl"�z���q��p���Y�ju�:ɒ&H�PXHZ*ע���K�>��GK[�I�F��R�IO ��'"a��U��%�2Ԥ\�(`Nl;�S4^�Kݾ}_}��qX�x�ܹs�kw��y�.����O�L(^���+7�I&���Ŕ�4�db�p�(���p�J�)lN�H�=���}%�
)�8?�=��;+�8G�[��{>����Ê��=��t�˒���,!�]ߤ��C�1�>Uo^RP�iz �����9����r'�'1w'��_J�[�Mu��ug�<��̤��p�	©n	lH�^&�#&�l-���!5u6�s����{�<DR�"+*
^��-w$<ڸ���o�0-Y$���2`����ʥ�*�8�)8����M%���_/B7o1����9�==�3x��M^�(Am�pT�9��ww:8�GVk�Q�����Sl��ד�1��7�9��Kh��O��/N__��2���ݏ���L�*�s�N�Rh��2��n�I6�'�<�I1�T H��:;��Grױ͍��J}�T{A��:u�Z h�n�B�)�����ΈL����R�@�J\F���P���aC�ȑ#�zGZ�N?���k�.��q��GW��mo�/�Jt�y�C������e�U���2S�F�1��������E)�?ܕ`"(w�yyV�"smS+�>* ��,T�4p�
^���Π��X����w��_y��nnl�~�#��,�aH��Y���{0����G�(�l�v�Z����Ȳ����T�@[f��tk��#Ҋ�_���QJ�r�>�X������G�)�.�1�#�ΐ�Pw�Qr}�0��*�H�q�Q�o$�1����J3wH��gϒ ���� ��[<]6����9,�U��Y�z��Uy4����Ҥ�Q^�pY'��*�V��M��$<a(y��ib�c8���Obd1�߂[C��m8�q�(���a�9�Rp��̼��Bq~�'M�c���c85dmp��b�H�u�B�Wm�%I���
Ӭ;u��)�䧢�;V1Iа�&ˡ9p�$T6L�*3�S���7\�SmB�V�Hh���!�)��]4\��Z6Ci���֬q�KD�Q��|��!�|U������9·A�o&l�J���#gt!׵�W�G��Prj�Z�FԼ��(�ew_��8]���etqnĴ�+��,ͧ`Mz�f\e���>����M��%Eh�^C�j8Q���/���$�qH����N�x��W�+�?��b˵�)�k7��Y�=6d,�ܻc�]8��	s@^d����R�N��SԀ�ANe��b�b��4��T�\�YM����N4�D^��21��XdW�R�+P�
���X�I�Z� -������3����l��P��D0<�dbC�lS�<�5�ڝв�,���Ș��3����$��3|*T�&O��qq���	�ޙ3g._���8D8Y��o
��b�<ј\3܅�p���+fG����I[Z��_��)n	5I/<xc�y�����ב˾���Q^_FpO Q瓴�~�ϊCV�G�[Y	������5��/}���.]2GJ��la�P=M�/��\G�N�p+\%U0��a�G��ǌC�H[$�=ډ�]�_|�'���Q�MԪ8(������|���$א����o�(���iwf�nQzN��PR�=q�b����.�u��z*\�ZMy=bDq9��ے��7���,e�X,r��EM��d��b�VGQ�4�d�z�T&,��6p��mw�:čU#N���/P��!���/�?)w�!m�IU=?�Z;���9��v��,�ԙ���$X,���l\d��)��n�2�_F'���Z�����U�*��+S�)�'h�-<��F��;g5��X��w��
&���eۈ���ӓh}A��6%��9y�l?����qD�(YM����8�豕Pk�)Soa$�\�%t`z�V�L���,����2p(���˃&{~�ő� D���NQ��R�@M(�c7�%��-� W�ןFz�>��/��C��af1w��{��C��θ�h<�1��VC)�$ӯͣ����K�Q.����.�Vq�˚���-A����N�38���T��2^��oTe����2�A�̯�qb�7�_aW�A8�v�s�%Z�z�QB�!l���Z�N�&�K]5 �
����Z��$���W�u\N,���	�,��و��'���f$��rx��ׇ0QV���V�dm��Gog�LB&�,	w��ʣ��94<dL�����^�x��\�t��-)i�lJ���m��sLF+:�RzW��ߤ8w,Ck�߂.����G�vw�io9��������k���78��`~i�Fhyv	���&�Z�G5�j��t�����aT�͔2���l�kN��jcur�s���2˭��FSK��g�,q�F�6��-[@�iۦTB>R/�Z��}�3�����AB�(�2��G�ʔ1)����i�P��[Xh̴L���{aU�aD�C�_�t����PT��0�e�Pj	%23�ն�Ą���ږ��\�"f��PE�ڰ�ƌ��bk�>�ffw�;q�b2��+|�8y��F����Bs[�ˍ����I���N9� 01����,bR����ՠ����<!XhK�9�4ٜ��vl�Q�֒� �fb4+`"|O��9�O�Þ|\Opg<@-��</z1j|#�<b�]�"�5h',A2��f[���9T��S	�젳G,�Р�DMJ|��+b9ƒb��~�P�E����{���\�w�A�m�jl3�T�E�={;͑��n�G�����pC|N8 �Y#]�*&m4$,WZե���e���p��H	q�'���e��J*�GE�m��>c-j�@��W��0�ٴqb�����)�h��k���������DJ���)@>��x���>)\h}�PӴ���5�ʋ�|�l���A(�	�b>�5@2z�\�A�)������"��LP$���l
��1yV)�@�@:V�͈:WG�m�4�
��BB�D�G!�,e3B�C� ��fs,ea�9/9d���a4Iţ��$|��m�6t��:3�}(����Xs���*[`AC�8.�V�ϝ0�z�����666���;j�^?;gԽ$7�L���ח�:XG`�����'��f�h�w������_f��>����ޛ��i}��1)$�ʽ����\�L�Z�;�H-��o��� L&��&�6baN��n߾-���œ�ƣEb�G�OUI�����W�AI�y�'�:�i����8�(��3���k��(��C��
o>���٧��d+���(��
�j.��|�R�f���9�LT��PE��|��>h�L5�l�ӵ��q�t���%/z$*��Pnr����
�lnn�:u����� ���K/nn����f��RJ�?�,S���u�k�@al�M�JȔ� ������޸Od���e#?@�̲�O2M��&�ā."I�0�������B�L׏�^2h86�Y�ƌ���^GPK��"R?�*6��X\�D�G�N�����gZҍ��L(ޜmzObN�e$��(%����yF2R���YFaf�����˔od3+�� b"���A(g�l���u���<��L�A�h4kw�߹E�t8�;Q�aC/������i�1�6�%��[�[❔��2uX�����,�_��F�s���ټz�@�ĉW{�>����w���M�49���x�߇G�Jq�`\C�])w�xˏh}h>�U, /���Q��X/bUi���/3��L@���%����p��Җ҇�����Փ���]O��l�ж���M0�,'�fTzg0�B��:�7�0Q���������p{bӓ�>��� ��Z�j��IUNq,8|���=y�$~Kj��6u8�b:ܹsG(�0o�8�e������h1�I�0��R��m����!�X
&yQL};�_�<Y�t�'Z��c�����`6G���ŋ���0bL
��!��A�G;;�B�+��Uу(3��u��hL��ƿ�S��vz-�6��h�몬]�+ڳ���u����c�pp���͙<>BY6I곝K� ��,��$j�[��bt�S�3��v��F��R���aL�[�U�%5�=j��(�#��:�g;j����9�%l5��r�L�g��8�k0{�smmͯT���x����N|�{	��K���Hyq�Q]k�������O<񄔍bBf��/����杍���F*!ކ���(
$� Oܠ�K����8o�	��Exjm�b��Q[�e:0�p�&9������e��Mxa��m�̭�OCD��37bQP�&���Ex�$�� ��=¾�+�,J��Q3����iļ.�]'ʢ�2���-��H[�3̓	��t0�u7�vg��<{q���� ���P.��&R_4<d�v]_ζ�#jr����_�����EeH��ӥ,	]���M,u2u�<͛��_��C$�S�2���yKl�rks�z�Gc�5|�F�YN$$f~�ĉ���@H(|%��j��יR���7��u%�c`U�d�xbjcs{��a�7�`���97Ixl&���+"�h��&i���\��p(�3c2��ZX�k_��R���k���r:�z	�xPH������ر�/5���4# �+g���׏�?�v���Y	���Ru�
�M���Z���(���2M~���fY��9�p$<��9��eu��$�����o���Ո��*�Q2�"ե�TN��63c�7N����(&���(yǢ"�\YH�L��S�_l����ne��Mf�	����a>TQ�������sJb�,ݵ�l�vrJ�)U4҅��8� P�Ⱥ������?L�rcB1�ca�ƃ��L�]�ϊ�(�U�%����>���w�a,!�ӏo�G,Ӣ��&��ۣoW�w�֗G��4���GS��ӏ7�� �h�Lü����UI�W*�s�=1,/�r���sΣ:�{�?�����ܻ35b��r}�:\���+"���q�ׂܞ�=�Ⳗ�F��V��ݕ��RPީ���'��A�0ӵ����a�dB0P8�j�ȼw�i�gR�3�ZsyYqOz��C�rqlO�9$#3j�'�n����\s��]��y��63#��kLnC��)�(��]�5�z��,�RJ�&�%�U8�Ř�D��Yȕ�d���=��iI]4�QN�"q��j��"8�\�M�@�3�Põ�c0��8tġ-�~1�:�ۤ�U�:@hPʗ�C�|�.��c��q��b�(�HR��Ae�PTWIJhY���g��f��9��yƾeƥA��S�h'��J�i�K�&"b�U����2~��xL�0Äb(�� ��Z��e�Y`�!(���.��yp4K0�q�%��Y�-���M��������=�CrF�W2����oa�L��O9�#N��'��Z$�
f��o(~nJN�����*a�	g�m�z���\������a"Z�	�u��g\�5Ç95���R�2��-�u��?� o	�GOE�M{�c�>K|:Q���3��d���~oԯ�[��`��'��	!#d��
a]�vm~~~uu�_�p����"�N�a���+Cm������*v5���ܜ�~�P���w���4�X&����Z����|�ʽi�/���A�g�<Y�4+�fʋ�⇥��ޕ�uu֓u���K��\\FN �᝘_L�ٳg1�dY{E|8��y晓'O}��_�;�b҇��@�VHL~�'Յ��Y��Kܺ�	׳?q����Ο?_˺�cB�A�lݼ�x���J�JM����`��A��v�԰�w�]Ek�q�n�W�VU9�� a)޼��i;~����k^[_�}?����,����EKYA�5�¡8����5Q3p��(��QR�&Bx��^�/"	"�ˇC]�Q�l�F{fccCQ
�>��o5Z��N��׮\��z�׸�P����?g�\>����/w�O�~�ٳ�/^���ٳ���@�ԯ�H6�3hΈ�m���:��b��;���<+G4M2���R^�ƍR��y� ���l��!M��)X�KNQ�Mr;p�;���P֐�O��T��%p�gۅ����n��Z��1S�F�&�(��0�8�zQ����Y�0�f�O��=�+\뜚��?���L������`���Ν[m*\���c[Q��j���Pb�-~�V�Q.�t���(!�������	3LW�i�Q됚99.�r��x?vd�{kw����رc�ԉK�s�(����T���wd5�`ܗ�@�q���,9}�D{a�Յ�1�8w�^~�w{~�`woa����q? ;�ՙ0�"L�O{υH�t��G���=�q�Ă\�]��[!�f}iy�5��bkB풹Lf��#jv;uM�#�lF�!S\K}�a�b���P��^�B������:����;��-񠷣���I���[Ԙ�M��`<���^6j"�QF��Yj��>���	��V''�}aaV�s}�j�fk���hu�$��RZ*Bq�'u��5�P�u5�n�JM�5i;������n޼G��=��F:մ��N�ׇ��`��b���3-�3���F�Ɲξ]M�`�}J�`��,�_&�K�B,���"'���3�dIQD'#��U��,̷�5�rth�N<������D���y�:%ѣ�}2����]�U�Tu���v�AFq���Z�C��33D��]$L1�$�p'�|n{{���t=�����x3����Z��s�gn.�@��01��D�"�Y�pҡ� ���;��L�ot����&�&0�{=Q�g,�<+/I.�o�iM:O<��W�'�a��Z�� /�Q��
y璉�S2��z׹�Ǐ�<�cl�E�8�������S�T�N��;����<-��]�ʌ���VX�(�ukmm��ͷԴ�5x�1!�2�!/���2?t�����8:2w�c�j![���mlP�7�/"*��,�x�r�/,$�*��C�G������lM8�F�Mϯ��77�5J��$Bq�JO�FUu��'a`��ܬ��
�n�$	��x�_|B+tɥx�v�U����~��$����;�$�,u^���/�� ��9t�x��Z���}�\w}���M��6۴�]uɒl�ز�����b�	%�HB��Kr�;8�p�́M6�ٸ�-[.�l�����������߻_y3;*6��>F��μ��������4�����.���wl���!2�B��:72`~�Y��K�8�K��Ŵ"mDw �.v�aGl��cL#�'�Өb�'0��<Z�zU۔��om�d���u�@N�L�M204�-	4��$�Ka;~�������Ư}����	��	Jd��SÐ8d�HY�	Rc������,u\EM��4�#���N'��m����i��V9mV�+;�u���#��+r�#����N�o|�Qce8��2��uv^�eGdH]Q����v�u�g~�{#������T$���d���"=:�6�KC>l�p������Q���zh1I��!�
lѨL�N7L)c�X�3���:7�԰;��	l`7�x�] �yX40<�_a@ �,��;���"�_�Ķ]�&w�m�G�ax�%�\�mbb��'��׋j�3�2�3^9{:s����{b��!�"��A�����g������<6����#
5m�3�M�#�)��U�d�6�mp;�����V�Q�K�Bp�C�<5�%p�
��j֚5��#�}���e���D�:�	rL�u#��̫%���d��THmx�9�
��Q���겁4�x�tL쩩�<��+zȒ�<?��x�N�-�
BA�`�`��L�i~;�e�"o�f������:ʪ:37vp2�%�]f��ߩZ=�u�2�.�]�}�=5=*-�m41P�֨;�+d2����\�{Tp,��Z�E	n@_C3�W)i���ft���j�L`�ۖ'�"�����������#c9Ԕ�|����
����-��5lK�T]��Q��bT���%z��%b�d,�J$�!�P�tPb`Z�Lqa�99oU*�2;y�AvCM`�b�=���5����9@�GF]������ Xo[l:�#����³�mycMEY�:���$�[���E��4��g��|����f2F���8���LF'5�%�M�(M�Y��UMJ�.��g~Ֆ���:a�1�FWƀm���E�V)�f���ъ�A�LpE���@���[��9���/����ՒY!p�R�P93�O���Eb��!�4��Y�ٺ�l�G>:�Y����b�2�"��׀���N�	������GR�b(6����i$���Ė��N�6X����Vf�캆����C�������(������`�ͣ��g����Z��Z����">�!	��-��>�C�z5�"�#%�#�5%�ɇ�/
���j����X�rFV�V�mˏ���"cD�Kx{1lA�;�Q|AUE��hAW-���nv�D��5=����<r�e3]�k�D�� �M�E1����UW��%�E��{������'N�[�^a��C�����CO�z���̈o ]��HQ���-�~��m��o�姡���2�;f�i���R�Ψ��ο��v-�Ю��Xdou�e[.g�

�R�q�	�Y`H$G��0
~�	��D����}ϲFIM�q��&b_7��'^���.e0HEq�/X!0�F�m�j����q@A��\i��$B��k
�*77nY�@�	����8Q���~��}���� ��yz��ф���h2Ũ�%��gtt�����/���t,���v#텀j
?�q�Q�,A�Ze	���I'nD9p�f`��rdBj���EJ��8�V~���S��98^�����s��ݏ<���`�s�~DZ�5��G+�S	��Ҟ��Tjչ�0�Cã,;��I��!��-i:��L8T�$$�~��zL�.����?`{ї�IT1��k<r�mH�����W,�� b�m��`
��~�B�	��w�GZ�e
6�%N�g�������,���u~�G���|��I��Bq�۸��VSG%bBۻ=�N��i����E₶1=�Y8#�,��.�j������h����H�s��ȭ�m%j�ɽb�j�ŎJ�s��!U�V9T����B�(�w��-
=�э����_�b!��f^��]�;��a+M!�~��Ӕ�L���X"�}@�H�.E�^:VԎ�a�L�%���[�����uG_��x��/,�RG�V��(��T�DB���S��#v�}}�����
# �[�W�,��>0�ʵ��+�8��X}d��ᄃv�W�󄿞:u*��3}@�-���̃� �R��(�!&�&�3V!��N�	Vl�-w�{��q����&���K2���/$�ѶJ$�z�T��wD���-��ӎ�!�d�ݽ�E6n�S�~p�,�V���F݌ǒ`:��ͩTȅD-�Ƥ�z<&k��ݿ,ɥ��9� %:�d��g�K�n]W����z_�@td�j|�d�K���m�'���U�\%Q�z�P�=lڪ����R�PT������	#���:px��V� �6TE=���2^�i�bst"��Q�K!�l��4���X-����)N׷D�C 2˱ʋŁ���	�^뤞M1ݰ����7/��d��P?�M&�F-�N�G��*�4Im�"��������"���T��*������/��x�}�B!�J��O�_�๵B��%��lT�^�1=��M���!�~a�\$"?)� �{H��Ŷ�7�� i��Of��԰����aJ��4#�e
�h)�S��
U�c����@0��:�r�Tp���X�����p
�^�D�mh���=]82,��7�p4~*&g`����"�s&F '|��r×�ӕ�}�|���S&K�1��E4$$�rB������h�R��k���%&G� ���F�3
�)h| `Z����ʧ[���v1����U�}[�aF^F�[�hp����Xt�"gE�;ku��T��5t�0r�Cb�"��[�����GȨu좁'(�.y��T���=�Ř�Ph��'D�H�K�]�%��◰����EA��课^,ft����ǯ&�d2@SY�h���8��n���	[7i�#�+v|���GI� _�b�1��FN�24�r(2BYCQ%_��B��ѣ��A6�>uJB��''Q�C��o?����͌�����#�f��?������`F�F���A����
>AO�jY�f(x
٬֓7A�XZ�P�ZX�v��\�3z��p������&��l������tX��1��	�9������ ��\_�ׇh�ڮ�N2Kf�uQԷz]�W066�w�^� �/��^J�w��A��W�����v&����ω�t��ZgG�B��;v��ܱ��9�4-���k5��6�ɀ� ��)G�� 2`I�&"K���*��D� �<�u�K�uw�p\A �\6��*Hlٲ~T��E	c6�`EE2n@x�_����$��055�5'�@���E�š��e�_[���	�Db��9r�B@Y!ji_��4�~�O,���#�^��ڑ�i'����z:�����i�W�"��pq/�:x?�`�U�i	���߱��=,
�=ގ�)��CCC���v횝�پ}{�{�}�V��Č(-��CN?�;�Y�^��
�1��/r�ٍ���6*Ql�q�0�9����%�jv���T��Q��k5hc���{�MxƋP���{M�T� ��bͦ(8*�%�=y�t�9�a��]�O�\���G��.;`[v=�?=߱2���x`�0.�3��e,E�(&�D'�gi�~sﰽ�����pH��]��`��$b$&S�~|����r����Or�O��l��h�(b�ۣaD��\%��w�}-�J��ی���h,mZ^J��揈�u8�w���/\��R<I>��[r��K�
�X��TzN��L/��}���G�լ�ě;�~Q<G�_�V�a)���rFq^l<�^�$��l�)9�DX��U���'��LXp�6�ZT�|�Eb$�X&ǘ-�@����V�!E"��v>C��\S�(:Ƥ��e�)tT���Q		c`-q����_b�N���;з�o�fd;�<�̰��(͵�����o���?r�yP���aʎ9I����@��� ^]`N]��z��\�!`�$S)Q��)�h�%�A��؉x�8}��|o�ڨN����Hhv3��c�f`�`N�9�=V��gX��Նi�]�AH��s?=}��矈놮j���wrb&ט�&O
�
�*����[U1�f�^P�(���2�|s��h�e�F!z�a���`�ư¯T��h�0<�K
3�*�� ���3��	憊PT����j&��2oq6H'-`�M�w�ԭ��Q�UaP8��0��*U���cc+V�\�L���@%����v�kZY:��X*��c�C�I"�=z�-K�yj�C��!��Vo¶,6po4�8�BOH ���.?���U�+�葯��h����cf�����F��UM��A�)e�X_��]�h5T�w�=S4MA�ᮾ����Da�J�N���:#~BQ".��f �����nԱ8%ȥR�m��-Ƥ���.�>lMc������{`��8����TG�;G���x�rp�?��-
��n͋��u\�5ʄ�g����s�0����8�)B��2a��`j�qLa���g(�%f��X��U�R�1R$.�6�S�nF���|1�%RV�r.d2��5F�����ZQߐ�ް�gA�3�>U"�nuux��@�A.PHؘz@���-������u���_�k���D�=N�c�Ϥ{_AU��ܠ���Ŏ����6J��U$��ɩ�@3bxS#E���<��ѐ�oQ�4$Q��~�!X�Tx&�<���l�P�<	�@aiC��K�z��|R`;Oז�j���4y5JTp��<V�2˸���IP��`os��o��]�R`��Vr.��}7 �������:C����tF���>���/�~��g�vh:�v������+;g��ēπO�7W����u��u��V7�6��G��f
,�L��W�ZR�X�
!�yjT�{�h�d�К�:h�Qq �*�H##Չg��.I�7d��J���E���\T�>G���`iώ�V	�)pg��n�Wf�kox��'''�+0���ׇ�4R����O6���-�ZW{�Ά���]�-���zz�p]$2"�Ц���7��I��@. �Iu1<<:���,���фZ�l�s�_�֚0 �C���?#���dG#��41
�p�Ν4?Yd�$o/8���un?�r�	�ĭt:ms�f�O�Fs���#K�-�4o��[�~׉�k"��R/�P�,>�F��j�*D" �fuzb	���1�H�օ<��ʟ�?#F�J�Z}��>�.�@�/��a�x�b�?sN��+�P�@�OB���A�Eh����0l���^<v���t�( �@2+�E+-�T܁jx� W��{��\�"���sw}��xQ�ڥ�����C&'�?rP��faG>������W{�X%({v�7��ח0����{A��n��Vh�����[�a���N�PH��<����l_�}[y�$_�+X*��Y��Ɋ
�(�&Ӎ,��eu�P�6��V+x��E(�m>P[ �`π�c>���9V�qk�K��C������;�Z�Iy���8�ǯ�-�vJ,�t6=�Rڑ���y~a�?�8(0xr�\���e}��
�K���⏳�e�'��9M0�K�_��۸qÕ��2���)��I����Ig�n�}ݏ~�#.{[,V��ɩН���_�||͚5��>�;�����p�Uj+71���}��k:�y��4�5Ϧ�g��bs����w��P+��}#�z���+׭����,���]����f�#v��ƭ7~TȦ��%�>Db�.�ڥ��������뉘:�Xq���+�
�ʼ�.{���~��!�#�]qeMî���7
A�I�;B�P_zp���B�`_���e�A��.7 +J�u9�cfZ��S����L�wu&�{���LMZwɛ����x�[;v���|C���(ި�ʒ��_X�ˎ���+��'�=d�Ծܖ��N�Q�5��b�{��Dܥ��2��셞T&�%/�PX�@��)U�-��ě+�զU(U�T�v̡�,�م�����������0P^���]՝�l�2=Q�q�<ɸR-W��/5jV,V���eu�L�!������K�P�W1Wb |��tXZ�@��*��Z�'a�6^����Y,�P0w�ȿTM�$��	������@-^�fE�Lbt�0��^�U͆�����O5jeI�C����fI�zZ���M�j�@���m��j�Rub��d*D�n��8Fz4�?�U�����
��A�Ѩ�#ѡ�;�Ru���#�����xs� �]=X�n�*�f-�e٪#���R�e���f�']\@�_�t��X�����V���ʛ�Fɴ�����S�׋�y!��y��T�EE�G�_-�2E	�Z�A��KhyOD��Đ��첗#;¡���2o�V�� #�	d�'	f@ֲ��Y)����|4T3z
�i��*�^xE�e�ٌ�z����H�#t���DC�!vj�(P)�ǂP$[!L�������>���{[-0MY�A �3�]�&f�]O���d�������!�`�1�bA�L�1����1/8���:CV[��:*�[�w�у*<�%�<�ćM٢vXk�X	&�JbMF�V�r.�l�i´m:��V�/�rb�Ț�+D��C�B����"U(�Q�F�Q9?���e�	�X�7OΝ������
�x�l�'�SH=�Tj�lpdE�a6��k��庆�����݁ށ�ǧzR�)-S�ќ�0g�G��*� �r��Z�ѩ�
X�޵T�%BV)֭
�f�Fj,�U��'�i9ە�[NVu�F�MϒB�}�h9H�ˋt��j#�b��d"�A�> �A���	Ţ*li�,XŶ��*�Q��i����y����L��(lF�c2zj�Map�س�������uj�v�UXZ8l�>66ƽ�_J�wBgۯ½�+9_P�]F:;:�>l���^
<!����@a�w����ڷ��m#��/m�Q9��я~xjj�{����J>?�5�� �����\x���eGFF�o���Z�n�N]Y��-�
ˤ���
���ӈ��������p��~��o��&!C(9r�+`4l�#t-_c�浯��j�ٷo��灇s�,:�"���U�Bv�,���W�?�Eźj7�~��	.6kBǈlF1�X�b�ѣG1m�� ��_.d2�3L7�/�]����ȑ#t`��|�`!�Q 4�����/�;o۶+a���G��S[���"::vC��"�/�U���Ko���/|�p`V�\	�߿?�s���]]]���)X&�R� Ŕg�`xHkS�8n@5�"�FNi��/9����ԺDXQX4�S�����.mu�E޺P"�?jk�5{�
�ؕ�a��ULL�p-��`]�?~��kዦ���;��κ��� ����QY�5�S�"��\�q�0L_�,�˕���jqm���FU��T
�d��AO��9�2�"a����T��x��?��SSx���k�k�@�/U$-�J
�p��\����*4�|v�\^\�Cef�\)r&���$zS�	m��R��?x;8�b�Z8^��>U�Ғ����s�@�vH�$vzƺ5l��a���tQ戮Т)��2���Tp)Y�\�`��x��DHQgc��������zH���g�����NtBC~N�C��A��B�����w&H_pa7T+�	��Hy���S�V~폰�&��S�ah�`:b�%�BP�kI�*Pn- �{�
�x��
T����E�N�� SupxlTP@𤠀�Tr7xN+�5�����+���?8s��j��W_\t��^�mKmd�PE 4A�2^	D�CV��/5�nh�qQ��&�ɂ�k������_����tR�֒�/���=��Ѐ�l֫�����C���}�s��?�������O4p�xw��xwtI�0��������.3�&��q@�����������יs�#�V����s�3��㯻ir׮�f�o7�o���/���!"�Td����Ec�.�<|ek���׿kω����u�-�G]Sn*��l,g
آ
��X����'@�	N�K}��
�!!?���'�d"�=�v��]=CCBzh���T�[������ �q�X�>�|�|�X��~�舞���h:gyR��M���O����O-�ۗ>p`�*��1x��Ҕk��j�f!; �Ȥ�P�}	|l]�ɓC/<	ܑ@�BĀ�)��/J�*�n�.v�m?�����4�V�
�,l�O~����.B� ���¯�x�+����7N�8�aÆ�Ї��ao>_��`+z>b�<�oZ�����D�AYQ�-���5wq�>Q2�*�b��3���ue�PA�b"~����0��+>�3��Pܾu�p�W�P�L�+G�g�+'�N������q�C��p����>��YA6�X��X�խD*��` k}�J���$�{�R\��;>��p�l�Y�L�Ѵ뵆KͦiYv<��\�t-�dA��#X��_Б'�ڬkF27�y����C��Ε�-[�������YEOLM���.B�^3�N�I�{j<t����&���3ʴRw2س�'p�)�8�/��u����ҿ�x}Уpt$��ria�X�dr 4&�WOLN���˃�H��H#%�#8�5Y���I����@��NI�!s�R�6���b�q�v�c��GHb�F��w9�f|G��(���"J^�l���Ա�ѕv��b�ZK��g���4��w͈��!����o�	��{؋!`1�Հ���
�=��݉ ��nl)
������=�0W����n���PZ��QI0�oǅ�к�q�=����Ol��U�C�Yu��.��ѡ5R�>,��I�BITzj%:�
?p�!#�����J�d�)��#�oa�����{\ ��Oh�0�X��~L��]�к��O�YUttERq�B٦�r�����H�=э�f��byq��ib����/��� ��Y��=�����&�o�� ܛ�h6�����0�d$9M*[B\;���[F�Z?찍�*,���˩�U�V	/~-�Q��g	%���LOO#㍦J��ıc����0wp���]3Po��7�pC.�Dl9#��O^��*��.���{���{���ڹ���׃2 �3~��O"��������z�5�4k�J	)��&���7��R��X��M�6=�\w�W\q�=����񎷼��o�����σ{�t��(��Kd�Y�j��I�-�%��?߶��������II��	���I�vҔ����1>5蠳f'Ϡ�o~�*�ȼ���x��k�33��|�;7\v�̠�CU���L�����+����F������b%����������J}{Ud;5���`��o�T�j�D��i0��&��ꮄ���<t�Ƚ�����}�
��Ѿ�Mo�馛��^�c{���q���?��?��?�Ї>���~7���� �{XG�+`Ya�1WM\���������Qw;M�H�S_�b $2E2�ٻ���
3`��j�&o��&�j%��"e�{��É��ҡ�|�ۯ�����ڲ��V��]��'<�-
�Z��́��]���دĥ��6�\%<��c·�6fL"��]�#Y.��/ɭɭ^�z�ƍ|��(��X�ϲr��?��?��_~������(��S~؊/Q�2�N��W�_"Uߜ�n������s�/�:��A>�~��);�����2��S��##�h�$�������F#9�c�Q�����<�xZz��� �rH�񈈭�2K�i���6];0�IG��0�3'�FGG��/?_�ch0�RI���K���9��y���ߋ^Qc.��)h��o�E������Г���l���hj���b��������:)�fѣDAV�S#ҧtv���7��gܧ�C��+�!�p�NP��搘n��Z��0-x���[��N�����p����YڹEP�]�4  �\xt"��?�z�V�p"PR�u�@�`﫩)�'a0\���M�E�"P�%��:oo�3��(*@?��{{z/�첐J�9��bג�oG<r�`4�I�_��&''�vLL�XX����V��R~YĖ��re|�X��௯X9C+�vܘƺ��/t亢�cx0�~$�����'�]X(������TyǏ���"C��\*ޓʭِ$�����3�����c``b�CAW�ES�����t�L_vd�h<����Ǐ.욨m�t�{��5K��51��>�{�Ԁ.�3�	EmY�(������=���pLZ�������~�h��~�:� ơ���ML$�@f��Q=9O"ۅ�	BK��-�GKU�m�V踪�[}���Nն\7������ӃH���b�j"�ɉ��
A"�Q�-�(�ѕ�Җ!�`[������MOO�\�j'6(d�Ấ� y���]�'�izB,#c�i��ו��0_}șE��d+\�����a�'
�G>�8?�v=��O}�#��?844�^�kP��&�B������eY`�L�Y�����r��oz��va=  ��IDATo����{�G�)"̀�H�`���#ԧ�����7[����y	3�S:��w��I��7,Ĥ *Ç}����Ph�=�\8b��b��x[\��\<I]?奰��⊾�5�	U���C`���=�ڵk�m�Hqj&�ɮ��'�r#�셏/2b0�������r��+h1�	4�2�1H����Ӛ�����ݘ��l$��^x����Vo�v1�sZ,�����$��\��KJ�����w�X��S����	��͙t
��bق�$����l�ETI��Dp]��|	&�tdb���V%F�X����5I,�R��ĀN�1��{q��X�$�j��T@�V��+�샇O�>Y�=y�/h��l>��A�4���������2�mM�UhB�Ɔ�K-�5�	�_��t�ȹmz�:�ePѶPK���@�Sl#;o �|�ԾA���j-�*�*{�{_U<���K>kԛ@kߟ�3�o�z�" ��\��q	˙љ� �-FNa�T���{"y����e�0 MK86�_Ǐ��܃Ѣ/��w1[�Y��́Y��`_�U�bZBPb�_e�����PdHiy�b �X���F}b�<7P0��Ji�^Es%����F,��&��;?�'���B*- z��� q��0B�!6��{����g���Ӵ��ۘ�,�]ǚ=CG<��h� �PM�����j"���ky�k���H������вap?��%��6Y��d�Q)(P>�s���E�{)���=����Zڝ�Jb�1��.�N�)���:xh����|�L�ܭw�sj�vY*C�W�`�p� x�ä�m#���6w��	?���u�0 �Y"��R�P��?�E*"�������qn��9Z랏;�a�:P� ����Ǆh06�0�숈�ry�'j�z����"��,/�[�]<�g�������v�ӟ�n݊r�#X�:6?��B�T� �P��*6� ���{��h��/Xe�L�NL����f��V5m�c�O>�䩣G�`K��FZ�h9[�НՙX�@��$%z�E��s���ۮx���� ��J%�bIXY ^����I��L�-���9�m���9]��[*''W�\�D��L�v�C���?��hx�VIAF$�KY!�֔�E�Y�>˔���л����<����)n�$��ʁ%�������G�\}�����>���|����ޙ�]�V\|!`Dj�2�Y�F�;!lFuS
M��!@�5�H�O��r6lx���6��ڲ0nċܛ@`���&�����n	���y]wݥ{�>������?��x�H�� ئU9 ���{n� Z��������::�`��(��,��d�B����N�,}�|�+^�?<�SJ�{a���,"0Tx.�/?��W\���~��/~~�u�A.�&�4ta�Pve$�U��SL�C��c���m��h��u�z:��]���r�Ag�q3x�����(�wN�`$0~���1&F�֞�N"�����F1���"x�@�/=�����0�� �d���(tǈ��
2�]Ol�`�Fճ1��`���~���m밗@Q�2��*�\5������p*aeӉ�xg|�vB�&��/����K�ZOqƃ��$lPdmy�(T�,���Px9N��J��(R��Q��-7k��a��!�� ��Q@5�V�f��Mt�Y�IX���<G=��!&h��jp�]�|7�Yp@`����=�C�_���̈�hԧ��pXx:_�|~hh�Ks9���~�YjC��V_��g'�Îs���,��>KQ�&��u���x�pu/6$%e	��e� ��W���<$��z�z����~��R�6q�i��9�bU8>�x�Ut���|"����7�6G �*�����������ǧ����x��%M�/ �/N[a��}����nb+0?0� /	�|�,���.�|՚�	�#�;0G�x�	A���h\����^Z�@�T�l�o���`�=58��©�97��lX����4/��b�*�|I���pG�2�BY���gp3	�ɹD\BL8�ΰ���źS�_zQN!���+؞9�Mvq!��Q����,��j�'���#�ǘU��&F}Y�u�P�J�c۶.,�G��ɣ�Aƙ�R�T�mc���^�Q�V��v<�:p*A�0��;�`�C�K�z׻~�\w�5б-�i�W��}����q[�kN਀��Gepp�����n����~�����7��":
�=����J]T�F�9]_�B$1�ů�2WTL����TSpZ�"j���p�.L��"x��_�z�ڱf@M�VլۈٞY�/U�Bqq��1�Hzgg���1�g}��IU]}�E��W�}�M�}�ӟ~���}0!��jY����;�"fQ�29$�"^��
d�G9���T=��1v&+���<�LM�^�ʯ~��]�}|�Ы�+ WR"^��533���:5�M�Կ���u�����O�r뇾��;��û���a�*�zo�a�lZ.������R(���8BЅ��H�󐊼��;le���<I��庣Inth�N��T�'���c� ;ɂp��r��q0�z{Ə�6�X$���m���?=~�_����&L1�仈})�F�
�_���O"q��A"�!SE+�鱸k��G��]���y��v�MQ�}��A95�͹$�~�3�>�}��\6s����|�b��s��!�W
]�t����EzM��j��5KVa	��!~[��,/}JAP�E�O�Q�;̵���,� M�H�� +e�%�θ�n��](�̓�ձ�n]I����qS��xdfk�k����ag''��Ӭ��k�[)xNi}B{ WA(��I�ڞ-�q��3&X%AM�L��CQ�&��c;�E+��	)O�P�}C�A̮'����ǡ@��~��R-]�Z|���B�[��݈���, �;���$��1#�T�a�,a)2|�B ��J���O�L��8� Y��9� N�ށ��:u
���ϋE��Pmٲ�ĉp0Yⱒ)+�� ����RC��fi��m)_ ���"cFx�K9ۊgt4�Ul��X���tx0�z��Ú��YxB8��"�+��r͚5�!��e��Bpj�⟜<?�����?����\�[Xܸq��o��.��v����)b�Do_���T,���7����w�}Ǐ �=�B��v	�6�~h�jDVEާ�H�aeAS>|��o��+���РH�A�$
�*��~u���6���ˣ��.�v��rαN�F�G����/<����뮻��A��3^�1��H׵|���ʰ� @�)�������/B,�m���F�l6�g!�_Tt�vrFBh����NNN�6Z1���'�,MM��l���G~�~��\"��O0�l;Tb<6�0���h�ǎptl� ѧ2Z��?��{��7/�6�H�q�]� �����pA��e�� ���6���ȗ��%p���o�f��ݰ<�?�x�yu�#�����9a�,-�˲���>f�g_�s��n�z�k_{���<L	!ȩ������'�`Vk���r0؋�y�Kj�:���Px��a�m<�������u/��G��������O�sWm^9:�L?�w0��N�!*={82 e֬����׫�](D�1��}>v�������`߾�<r�ȓ�=�v��?���]u�U��˿z�GV�,C��VĄ]��W�N'��;A�b)綯�~d�JU֛B�]�06��ML����R?��^>�aÆ�g�y��Gzߟ|�������������4��E��Z�M�@�S^��"k}�X�.0{�p�<g��K������
�
�93��N0G`n=/~�ŗ<��Qx��4�)�c�ܦdI�]���Rθ��[3�D����&H�|o��i�y��7�'���Bk��+q��o+v�9�Krg���Z�|X��N��s��O׉����^��ܭ��N{�Ƕ��S��GmZ�>>j���_&� �:��)D��){  �X*�M���I��
|�M��ᯠ,��Ax�7�8�G�1�x��Axp.���6$<�B$�qn]hQR�
����Ac�\\�%Z9�� �@���c^@�vs�e�=���LeO��~��Go��f�T�t�<z�����v�Rin�םN��?������|!Fŕ������_t�E_��ߩKl���������7�c'F����S�����~��O=�Lq_~ A��mCƆq]�s=Ě#�\5˲}�	7_t��q���cKPt���W�����c��6��<��}�kG�N���¯�뉑.,��m���J��t���tܐ�[��9����������������@,C�m�a{���1$-t�}6�Tmۓ��e�ݽ���:�d{�\k���x��,I/�K`���.ط�&%�H���U՛��+����>��ј����Wi>�W�x��̘����.,,Θ��K_&_���ܹ���+n{l����>����4��\����f�vlU�j4�V�u��r����l���ѓ�/|�3��w�1`�1�COtO.�ܹs'�%�>A$q��D����!׍���7������O����ǥR%����FU�8��֭LF�bCp�]�7�4OE�F��sq�Aگ�z$�B�z��?�����{W3�AO��؂��!�V����d&	'�R�Mk6MOՍLwR��H�y�<��E�r�'Jp��rӎ�n��7����?�9�+����a��1
&��e�ML��q�9��&���#2t1��Ѩ�]��6��l��g>w�;$�G"?AD��xy?L�T���6�͜����b���皤��T2����<�Hռ�6^v����O~�?y����W]�Ŕ�7�ɉY ��J2�p}	��J̳�a�0��AH��$�?p`�9�=�c���>�TB۫;�Nt�)V��zʹm��9'jv�0�����dc�oH�r�98�e���)��o��?���)��T���d�`�w�è:οeb9k.��<�c2������j�0�Y������}�if�ݤ�4ϵŐ�$��@_v�3�>�Z�˖-[�����d"�;��&JE�nWn�ɓ'�a��D*��iN�����a �梀�������)#��QXg)�y�":`#g�I7�C�Y�����|j��qpmL2&)�:bh������B/�N��-zz��؏��1xS��n����{�
_�-���TɆ%�^��1�S��ub}a�l�1E��{��ܢ�k��|OO2RŮ�8��J�*E)���d���krӤ����ή���c�>��]	�kfv�vq��m۶���O?�{;���]�
3S�J��,..�����xLh61c�+��]E��xsrY}4��	�=ҩ"z�`I(�xq`d`��'�/Q�(F�<j5���M��߾}�(+{��en��g&���ra� ��&���4c�)Su�Ig�Sv��o��˗/g���O&KR�ȇiqc#����^e�q*�~T#@�!v���eBG�INu��?�%ޏ�ɀ���*�����1�,5p��Е��%��}ya�1�����=��~O�lp�I�@J�i>���_|1��[�}�K�]�����Z�ܿ��ƍ���>7�ַ�u�ȑ����p[�`.�����hiڔvc��J�	������-�?J��tM��L��4�e<��?���������'{�|�������W�����i!(� ,[6�Ϩ�-�E����Z��8^ą������D�����'a�(��\2�4_\ �D�x��1�F��#�|p(���'�ş����G?[��=@�2�&h���r"��e��2elɪ��◿��g
�����6��V\\�C�k�+�f�cZ��T�|��+�����o�p˶z��Ld�_
� ۭ����ѣ0-�7o����/�5	O�cǎs�4w�BJ�ɟ���9�{�}�-���}�����]�00��z��`����+d�r!��E(.dŊ#wf�$��n���/O.��fga�&��/��ª�k1� ƥp���2LI������f�7߬���L$�.��P�0����v����mp�?��^��o|���p�W����h��n��1�E�׍��N�#����I�j�(	B�#����|�0�C̔��h��p9v�0�[�<�m8�b�%(I�'�d7�z��c�=�՝}��^�������;���?7E ���u�W���Q�¾�eq;�8a�ਁ���q8V�Z��l`�������b�а�ߪs��z�O�s`�`e׮]۬��,"L�R���������G��Q���Ȑ�|�:���vb�Cg��;G�*c�O�����$�G��E�)��
EN���l�z"Ry�*�X�
��ch����Tխ��`�a�d ��\N`�؞S�����D�ͣ�	<�a���7���*5��E�ư��6#��ba��7_�V�eT6�nUN��K\,���`�@t�/?����@��Jt����@��L%P<L@D'|�BN9�}�^�XZ~�Y�"p�$�?{Q'\��]҄����ܰ�%*e�J'9�@�NtOO�P�/nڴ����`���D��PW�W(�&�t-�F�s��&���q�v��*?�s?�O�j(�h!�����6���~O�U�Z�>u#�����k\d���)M�E���.U�HL*Ϭ�����	�����p`��P)V�&N4 L|�@�ĝ��CqYw�A0�d����g\/��A0��0� @"��w��l,�b{��y�k^����Y����E�"(��1}�?��^���Y����v璍zu���4}c�)4�t������;�񎫯e���f�TW�J��+=>1	c����{��_����?x藗\rɥ�o�n��Vr,�
R,�ы��,�fb� ����ʋ$�	��,/<��C�=oZ]>9���w]��L�s�P��+��t^b	ae.ޘ���꛷~�C���jyt�F������뚮�{�'�
sr2mV������B��5����$RA ��Z��˕��i�2t6ʰ��ꚶ�̯Z��*[fE4k�&�zm��hn�Z�3������-o��G�v��ڱSWn����-psz�Jd-W�L�H�j�+.΂c��*��|�P�jX���\GrU�.�� �ɮf��b�$��%&���{>&_�ڱ�u���%�]�<I�D�eb���0��5�f�暫�O�η����׾���+�|����w�3�B��i6��Fc�<���`L
s�Z���~�+��z�w����w��}�<�XH�<]�7qK7�jyV|���j�\,��۾��n�����t �Z��ޮ[p8/��U/���܉� �+��/{9��w�����on=���0�;���%-[�Q��S�XZF�D�����È����#��w����Ё�/�f�u𞩩Y����8���H�1r
�Ss��L�D��#Ӳ<w���W�b�_~�S*�J�7`!��B�q� ��L�R�y��&�NZ\��S���?<8(86U�R]̅d��@�1<���o���[?p٥�n����B�X6>�r��gD�ζR�̍s$ #�LSI�DY�#f�� {KK%{@PT�!��$tM�8��Z�D�Mw��J9��+�{S���Q����y�JK)kIN��Y��y�|l���n�V<@�`��ؕ�J�J9JQA�"9FtX]Dr��Ϣ������$c�
$P��@L��J�C�=1�zF]��j4�'�H8)`�N���겑�����Ǟ�����zC�[p�	�w݂m,̉=��%xY
q<�;�S5�+��� &�"�*[1P�O'��[�4�&B�?!�x�p|,3����h'O.,�/����e�JuVd����C��Vܷ������2�O�W��Գ�Jl,�J��X�B	��'�B�cK:,a��n�u�>e�}N	�ߨ`#�~�	��#ɧ�I�Q��/t]��$7?л\��''g��ਥR�Xd`U�DR-�%�1�)��7�.:|t2�GG���G*U<�lQ�@�GƓ��Z`Ț�\�uwj}	�dJa˾�Ao�B���Jݶ�:��nD��^��[��:�������e��@�͟�q�t�'�'�����������L"͋~�li1C�#iO���{n�	�?�Q1j��O�O��!��En�Tצn�����!�H]�-�wP��靏�b�_�roIK��g~ �����|�=��U����G '���T>��bmq|����;�cߞ'W�\	��)���r�/X�Sc٘�ݿ����c'&������5�9x,_]>���c�`7���7oٲ�ޟ�J��*�P�D��� [��|4}1�����C�br�nĎ����������cf 	^\a��\�����p�SOyGJ�)9���@�U[�����XX���O�'�p6�	<˲�Y����I	�� ;VK�'Nd4잜������^�bE��vO`i>|�9;4������J[�eKfٲ��A�9Đ�We˶j�
ޞ!��YkUgÆ�z���"nc�N��ª��hdx&�u��x���������^d��T���7���/���P\X���{������x�:��y��6�C2����b�>�m�Ew���W���_�����6�E]����;�(���W�¿���W]~9�����h/<�Ȫ�h����׏=�j�eC}{'��������իW��_}�g���W��p�f������OiD�UÝlY����l���7�x�����a����U+�}��T
�:��vm��4l'AB6���|�X��g���7��{ߵn�z�긚VC�*%l�D�� =t���0!�[���O?x��w��۶��o`0��XdM��@�R� �2<�=��|�:�k��;��X�X��n\l�#JpȥfL�ą?�cX����15U!Y����}ð���^���3X�d��T�y�`�������u����$�$B!ccK�8�m���,��C�K��f�ܮo��=��$��&v�v�!\�xj~aα��e�����`V��~:���0��M�8	�Z6���&R���9r��G�6���Ix��~��(���&�4����H��¶���B�u�d|�)��9v�V�\��GR����Z������D�` -�����~n��T�x-	f	6'h������#�k_�,i�J~�����u�T����2�mċa("�0��@߃�47lT��MF���QjG2㜞*��C���L����?��s��>�]����2��`��L��1$G'��2�0֞I�\me�3;��|X�n"����<*�����'>��� |��K979q���8����@ ��:�p�U8���Mg�[��@&;�A+�t��R�D�+�'�<|��X�w��sj}�w j��D����m"�p����mۮ��^����
�Di���	K<*��7�x+˻�0<�����?�w���r����]����cՅ�K��j؎Y��7�z$#�����~�㫯�����#cL�,R��&bm=��_B��p1\�vM�����7��� &R�lW���ذ�T�	�������h�L$.? +4�~�9w����������>}�����y�nZ1��+��±9�DddF5�tɦ���(��w�w깇�o������8�_����%�n�K����:ϮAi^����:����1��劙�e�c+=��;;��[6ד��%\Ks
�&�������>�Y�=��#w}�U���]��jFX1���*3E3\��zEq���� �w�ߡf�*\1Y�ؠ��@�=ם��tL�����j�����,W�D<�`E�^�x��A\��W���T�J��m7�;��KMTA��ť�	{t�CO�8�.0"�
ܱc�m�o`m���{��y�'n��M7��?��k"f��'&NN���f����7�����o���Ν�M��dw"�amO@mQY����#������$�?,�Ɍ��\�֜ �QO�ə�''����r�H>}�����o���j���ggWl��Ǯ]����}��^��[߸qC���:��gۚ���Z4m�Y1��������ġlvݚU�����'?����n�)]�=t� 5D�:�K�,Q���|,���-o��~d�����rjhaKj��,���A+�JW*>;;�i�J���M���;�o����,�|oX�7]4<���H ͮ��U�-ՊJL_��؁Ɇm�n3D���*����I�hHڑj� ��y$΋��'iR/���G��� �*�r�^l6��JѸLj�ڌe�dy.���IN�(�����}���|�����9Z���Lw��j����|6NM����zc Lsݣ`G֫'1���USW�����"�,�冃L���mq����+��#��6�g[`*�Ai���,��,Vv$�[UwNJ����ֳ0;s�����r�j����U-Qw�B	˴r]��م�\��MMÝm����ˠ��~�U+]>�}��Á('ҩS9 f�e����E/�Z�fu�X8t�8U)�E1���ܼ����b��N�9y��Q�=�~��[�}��`�X�<55Um���t�Z���?��Uq�4t�
�S���w[Z���R�f�j����!a�@D�DA��蹽��3To�vgi��Jns7���<6>�ı�l .�*��Eӭ`�ܵ3]�=O�(���_6V�.NL7F�~�S�}� o4g���5� y�h�E���L�^����$$K��W<Wt��l"��BJE׌Zӝ>uv�y�.x�[�������j� ��TXN��)f㆟A+���j��-�4Sl}2�lA�53 ��������y��#|2 ����"Ho]0K����-��ڱ�/f�P�l^D|�/R�yn_��50\���_,p�v����ב֘9��}�.��WЍ���\���?���>~�)��`4�=ѧ�l�&�Œ���2���7n�� ��u�����~���������_��+��~HM���1�:axx��Ba!S���ڙY��fRiIZ�ѭE];������͛�J�g?�8s�m�Y��7�����]w�x���,��.�V@F:�/L8�����ZXXؽ{��������NS��]�y2&i�pP���*�a-���H�@�7*�� ȒU-��b��jV+JyƩ>[�������i§���x&s艇�9^3�w�bX"����!�|bb�޽`T�
�7���~���d��o{|�<Ը�R��Ӿ��V�\Zܿ�zr˖-��E)-��r�|na��|D�s
��@�tuc�����w��x4��7���/������	���"�M�qǗ~�ӟ��]������V��O�:�!�f||��_h���}�Ϯ���;���������[��gO�_=���-�ߒ���`z1�䣼�eEM?�y#�?6���PE������X���p7'� �I�J����uמ�~p�m��������)>��`���Ā_�������߹�;���o����y�鞞����T�`k�:qh׬׼��?���^��Wr\ʴL.(�i�_����靚A�)�+`?1�x���@�����5��Jd�������m�.M������+�Wz��ē�`c�x����Ad�a̞�ѣPV`�؁nU�q�H)�i6똝M�zu�eO�옟����dU�7~�[�+t��ݓs���<
�������꺫��#��u���QAEL���KF&29��t�]]9�����t7�(��}���~zj��n�{�{�t���#ٮY&��N˘�=p�?FpH�I�X�f�L�֭[/�;�����Y�{����l��L�	�+M8p �$��&x<S�H�K�ʖҒr��iG  J-İ� ˪I��Ϩ��%�I��w���@�:(��j3T25�nݺ\�<v☬4�Z�J�âEagN�>�˟�[�;��ż55��FvE%nW(Ra�o�ϗ�Z>�+�X���[Y�wj|�ljꀏ����Gd���#�/
>V� a+%�mX;�OhpW�\Y*P�85Mq$ތߴ4�ZcK����MĽ��g[[�|��,�[Z�L �<z��[��+s�)��f��\�}�P<&h��dA��t��t���ͅ1���	:�QM�3	��>���/h>?�8�v�%|�f��5I��a���មJ�*���6yAK,ZD>�
��+�� �S�3Ǐ���&�~�%�ʦ�{�nM�cf��
a�w�	����j^��I1x�7���+����?�ǜ㚸�/lU�4�\����}>T�vĻ{�*H��j��������B!�HXl���X}>S�7���/:�d�Í����2A"�(s�ߙ��]/��{`[3�D�%����ʵ
��"C౲���$Q��Q�Tjnj�Z1�u����9{�ȑ�o���;��]��iV�yx��G�Z�E#�F�!M���#,"KSʩFE��k[�|Ʈ0����}�7X�g�㶰t�Ƌ���R�4�)L���dӚ5��0=#��E�ת��.�BiN��7\u�_���?|o(o"x]����ˤaMV7���ug˖-��#��b1��O�� ��� U�rmW��X�A��V���4f�l��n���(dGο��/��
��ۯƪֺ�û��t$B�F�}5O������N�**�ڲdpeK�����ܯe&n��?�7�v�!K��C\���9��`���X�*��D%�����v�K��A�=1�DX��ˬ����E.�-�Q�J�fﾗ~��_>|�:�-�����E�o�:m��-�E8_�җ�����Qx�IO�}����������~W����%�������}����[D���zB!5�1�2s�T�HB���eH���$�V�k�h�f�?����~D�Aɋ"��Ñ���,�P1U�.�p��ٓ�⾯?��'��o�n+�X߈�щUW)~�P��A��J�S�=���r�W����|�߸��'����[����=���|���[����R�N0HuOã#P��M��[�C��������f�ƕ�괋�dj
5�)�?�g�����LM�C)\�ƛdj��ֲ�k����b����"�G�&u�*(R4�O$����Gה(ԛ?:�dVZ�U]Ǫ����hs�ԙ�g�F�,CǕ�y�KQ)�8���%QW�����\w���� �Jm�=���4�Ew��E[�X�}ݎ�0;S�,e��J�����E�k�7+8�S��MMR[�:Ah�����0�X��8fA��(Y&���4R�:�C�v��Bn���cZ�+WX'v�M	���"�9��	�)y���KRI&��ç��֭hnlEuŪζ�V�u���2]B�ݜϚ��\���|�*=Q�M�S���c(��ٝG�$��&���!~��io_'ud� ��h���$O�g�*����p���:�C�'TA4oc]�&[�sğͭ+V]z��`��E�M��*W1%�"���tE�j�r��Ũ��U�/��eWE��Ce����S��B�f[���~�/	��p��E��	�R���L�V�C-�f�*ش��J����ݸL��RUH����L�q�)vS!�+ϦgmF�d�|��Ç��4�ׇÚ�F2�t�<Z���t��1���IG�4�"�)~�|b�������������M7�0�R���H��!���)NN�[:�<������W����'D������0d��{G9�~ �y���Q�x �H���\L�s��Я��M��N:x���8�1T������$����[}���bd���<8�	e�>�&j�`>�>33�X"���O?��3� �}���k��	�1��H�y$B��r�bj�`��s��9����1Y��غ[�l��A����w��w�Ny�dN�O��;rP\�F}Ғc{oWN�|!Mمh@oni9��?��t'��8zQ2?�ƼÜ��� d��֋���	U�!T̐L��'�7��lڲ>����׽�uюU�@���R���8|`�8*�>�Z��ʠ�s�Z;!� �5�L���䮮��x����׻��S���/��C�	� |
(t�|��G����Ͻ����E�����c�@`.'L�<p�u�;��F�9�CffR�O�V����B�V���+�?O2` ���', r��p�o]'�q�Z�↸<x ���O����w�T��P!߰�?<EkG%K���"�U����W�\{���Ї>�����x+>�㢈�� ��[���w�����B�����ښ%�`�2��]q��u`�y�l��s8�6�K;¡Cg���Gĺ.��Y��9�7b�(C�hˉݷP�T"6=x��Mo�����m���'[ڨs��%�J�g����g0TL;y&qOMN���������=w��G?�)$��!���}���n�^4+c�6,Y���ll1?����Y;?x��|�'�:a!��Jd�&%�n��{�+ΩS�Ό��o���h�F+�T�5٤��t�}A���� .K��-l���~J���p�eV���С���!G��*�xT�����KR���q*^~�)�b�X�t���C�]�v-���(U�)~��4ɭ�@�������7�u���$�aPR�0�'s���5-Bp@z�U��ij��%��*Y�rN�}Ի����ť�+D�YN���n�����殹�z���d��4�4�n�T�G����BZ�*�Dy�K���^���yn@a1�&Pa�Aնh��Arjz��GJ����9�+>��ۡzzz�j��]��R�rl����������^Ʒo�xɉ�'*�*Ɵ/9*eq�CC�+f/����-�q�3�����;㡩���D쩁�9/k���M�i��	��Kh��EÆ����f�ϛKϕ
��kw��l1[)R���>�����Q�t�@������z9[��(���%��.���b�??���Ʒ46�(�S3S�Y�r�W��%*����kV�tʾ�M~�xt�g?��72Bp��_w��-ێ?J0��2�O��f&gx?�C�a�ôC]�ݻ����gN���s�N��#u^з�:�UfZ���� �y<X����E��?��<�������l�}�)�l�~i�MU0�N�jm�`��]/�!
̓GN�NOg�ӑ|�L��f*��,�0�?�)�N���J
u+�B�=*�R"�x�P6m/��'�:_ ��x��?:�����q���8�Κ=�	�Ј�e�W-��b�'T�q�ԑ�x�?�̗5k��c����k��l�ͥ�_�tu
��7⃧�gk�\vr�e�>���%�e�f!�P;�/wU�RT5UN�XA�3s��X��^9��ǿ��;���x;�#jI˵\)j:v�S)��#
�Ȏ!5W�-�����6=KX��S�J���k˻̩3{�mp�ȹ'���w�j��R>��0̄i�uv
�D�41���i��X��Z'
Ղ�6m�$xz(Z��M�m�lUBY+�������_/ĨDcY�^"���N͕���j9���\���*��	BFs�G��s/�c�PTd/����>��o}��v�j�8|�ٜ0F�Fn{�صg74�G�����|��%ɐt[�$��%TR��������'��w�_��>]c�bp�l�>$NT��Wb��t�x~��u��H�JilMŭd��jŬ�IV���½��6qaϤ��>�QY�nc��QG�|����U�v�V�y϶��p=�ئ)j�v�־��?���>r��[n���Z� �����m�L�|�x<�ԥ�������Z�bӆ�����vS��t˶�e�N��U�hת�tŶ�J�5���S�������_��)ʣ�Dc�%1U�.�Z�Wמg�Rg;B��w�x��5[��4w�ݞ����IEu��֑�����t���_����l40S�C�@[�Ù������a��n�mn\���N�r[����Z7��^d[�LYlb�W'l8��b�"H��C�[Φ���6Oy�s���6_.CEa�%���I�)�J��^B����'G/ڱ�,��,T��P�`&;CD�F;f��mݧ'��L�f��QeQx���2>eٕu[W5֗Fϟ<q�<>�- e�-��v*/��G�����\mۺ��x%u�P0�����tE�|~p,%
v(f�~�?�I]|u��l�J ���%�qEzt��SY��K��R�a���`8_�=iK���[(��i��4I��|6VW������;-JEM�n(yЖ>LՕ5M��hH�`KV��_x���x��ՓS^�"~Cשϰ"Y��M5۞�hCcc�R��׿ޱgeE��1���L�W����P.oÍ��~/j�/ "�XoCO`�`�r���d&��I��g����^��C�+8��*X�U	�Q�2�{���8����ۑh�E��q��-��#ǎ�&cu�h<U�F�����D�h��S'ӹZ��˪�h�+f1��|�O�%��сG(�,JcS��7��?����u�00ЏU��M���X���:U��Z�_zI��Qp�?����~�I�֋�����ql�/����6�%*N|���E2�ؙ�Rc3�0Ƭ��ƧRC#p��gǶ�!E���i���7�J ZM�U)X�>�VY�-dֲj���k�dC��E�Dq2�j����d`_�������+K��3���Q��fL�����o}�� �:f|z^s�U�-��x�M�|��O�DY�*T%�c=��j�23+Q�;�'�x'�
W���]O��/ܸf-?y�/wA^6&Of(D�8$����j�Jak��Ç���twÊ�}�*�d��q�Z`��>�aq��=��n8'v2�rٗ��.]�A΀݌�.���p�'�-��e���&+��\0Y�~�;A���.S�b�@�ӄ����&F���S#O�@�n!��>q��uvb�p̈́�B����B�ym�4
�uAVaai��=F�x�WO�y�g����+�di����͖�,W�����:7�c�]�b�ttt�t�261����;��u������P���>}�]���榇~�駟��,�5��h\�̀ s��r��;�|�'?��{.�d!q��1T��@M��CqC2'=�-��ʕ"�r��Vd1���2�N��S>��+����ϟx�P�vO�s��U*��c��M��kV��̳i�ą�O�һz5n��{������{?z����퐚+p0Vm��z�>LD��ǟx�;��ܒ�W�C��4�^�b�Ύ�B��~����$�C�Zn��������wt5nڴIeH/�,��y��A6��x�
o��>|��e;oܺu?j.2��8f.�1�q��{��C
qj�IBaj������Mu���k*%E<�K��CׅcѮ�]�,���p����cXP677?��#CC�K.���qk4�3Q$��=�eVu��Z?��S��׮��9~r?�`H����Y����r�<5I�ڒ�A*�1���h7����>��ġ?����X G�q�
�RE��$�{(,
�P*��{����[�U������L��O�F�̆�ݸ���L�zPP��IҲ��v"F�*�?�O�D�nD�����1����l�9�g�bv���8� c��H�R�
� <�߻�����7��[o}WSSV����G�P�u %��z��e1L���c��5��� �ة�A��R%
����\��3��zu��D�sj�ڑ#G֬YG�]'_�̘2(�IR���$�݇o���H�fS�T]�ؒ�G��	c<�M1(���3T�1$^��׃�F�Їk�|�喖��|�++V��������(����Aj�1�</W
x��K/�UJ�>��S�}��0��2R�x��O/^}���z��:q�rh}^�������uh��
 �["��8q+�X��*�5�{).��|�-풒��H�)k��0s��P�<|�Ձo'�\�������.D�������Kwl��u;�julb�X�JH�X�𰸙�����_V�B�	�E��F�Z��Q����D�EVj5���?h��Y;y�����#�~�ګ���[�/y��q�ZPTѴx=�9����!R�U���X�G�5c=z�-��ڊ=� ��Y�������77'�{�	M�2���3�.�$�@��Ǜ1cYU۪X&A��R}}�TL�=���+��`�٠,<��O���\p�����1� V��6��J�D�����L:;�U�M�!T����XW{���0��U���Јq��,�}C�0�jnl*5HN�>I��l��K��k#V���|͞�	�|J�P�l�6��o~�{}A؃u��*��Cq�	��_�R$0��J�Mu�n�����V6	��"�CC{��}�G=�쳪*C���H����4Kv�e˖!��^�;�_�x�k������Djٴ-YF�J�Q�Q�UCkG-�������|?l$�q��#�=��#��|.͸�TF�c�F�:v3����Rq��X],؜0��g�w�Hׄ͛�,J�T��ssy�r�*c䊕��Wjh���۳UIP<�o�}I���6�_g��7��mo����誕���ĲT��y�5v{4B�<p���:�f���*C�iz����T(�ҩJ���F({�}�����?����Ȫ��!�2��Y#��K��%�����x�G�aX��(�]��fﳟ��Ν;o{ם�=J�>���~:]<~�	���cr�a��N��Mż��'Ξ�"�s��7%�!��ڕl:׷܃��TcS��9���^z�K]f�]��&�}��e�PMv�SK&�d�'���?iּB������҄�̶�l�:�¡(�e.G�ʞ`��s`����5�7|�D<���72FX~9����T| �貓�|!�ٴi5����{�j��JR�U�ͪ	���Ie쎤I|��4)��x�U��A�SZ�ַ��X(O��n�AM�d4����4�߳0O�=���p��Z�B�FOgg����չ^`t,����� Ɠ�suy˦��P�M�ԖƄ���iZ�j�6��d���kP�Š~�P$�S��;?2=�����m�}hٲ�D���_�jn V%����,R�?D�l�-�G�)YC��BZ�MG.z�;�o��'��;YF�S���cy���p�Vʏ�����.�2,@*�B�4e�e�I�$�Uf�
C�gA�򵅲s����p��0��et�V(8T�j�K��%XX�+M�� .w6��\���~��T-W1F&�p?�O�nܼ9W��3��a��0w�}��:��ٕR�s�۷n�4���]�>��t������N��k^"����砥�p�ۗ�7�MMa'���&>=:�W�pn!"FT4�Ó�T�^_�+�Ӷ�1sC�9{�-�C��@���/������?=x��Ճ=�0ݼ��ț��|���#���b�>��힏����������x��R���eE�1��﹒�����T��>HATYG�����w
E~�)����?���]�S����\���b�slXC%�+�;+GA��������7塡�j:��`�sX�Z:��p�X`,[$b�O����:>�8a�\_g*l>�X�G�Q�;�e�7� �کS�����=y�N�[��}��NaK�
łU(��N,_�ON�:13��hc=���ٱ�iF�A�b�"^&��,i �����/c�k׮}��硚q�ɱ"vE}����Щ�= p��z���F4������x���E��y�#�Az�u���*[�2��,C����?����{hd��ʕ�1-"���|���O�?��/��b�AvED��'SvNi9Κ"b�
y�lڰ��w�����G_������Ɩ�H�kx'L�����B�nM�}����2xf������#.�?���[m �	-a�н����V^q"���²
�L�e�`��
w
A��Ͳ���޳�y�����O`q{{z1����#"�� �6�{OO��!��@P��	O�+6�]d��
�U5����NcY����t�4~���"��G���]L�8���G�/�E��Ux��n������E�q���\�ιE�X#,�5k�`�2S��ʕ+���{3��Ҧ�F�!(��-�\
)���D0Dx�Nm�����F`�¼b��j3L&�g|l4�����׿���nJr2��Q;���X3	a�X���M:��C���.N��)�S��{�ϡ#�>��ϟ;ws+TGH�	T��i��b�B.��d��.:�	�S�>Hη����9�iߴ��k��F�J�hV�_)Z�c�P ���q֩����ꨦ}z�f5k�s��Q����	@�[�5���1��(����� ����/gL0s��2̋HR���H��N�R��*J~�*Ųh#�q���?�|��W^u�W\1;�:{�,$�bdh���e��?@�V˖Q�F�,A�_s�5�/ubttl��^4ݰa���8�Jrx����Z0��cgϜ߁οe��k;�B	��m���-'$����U"������C��Is�<�ᕫ�,��'3�ۻ�zj������u�����Ā�p�RI��4j�&�9b�e��c�*EW��\"��������W�YA({�'�]汸�8v	Q�DqZG0���կ~�E�/_ֵ���__�)Fb� y0��4ep���2��@�H5�v�I��2��sb��^`)y|'^��Kj�~��Y
��-4��6f��bŊ|.i�5#��7�555��]��()K	.�gSG%oi�Ă�rT� 1��*��%tMRu��(W�5&4%I���9�X�n�����x����Hݎ׽�	���Y;��]ȧ�����_v�:��ts)�p԰x�%�:==:55ӑ��F;r��T���\�B4��5���^U���5kD� �j�>(E��H]4?7)X�Xӯt%#c��gǇ�#���m۶%���ٽ�gU8����v\I���
�ҩCׯ]I:;@�JO{S�'Ōk���CL�� �v�ʕ ��B^��<��L���q熦��ǲ�F���wl�\�d��T:_�ȑƆ`T��!jL�c�����Ԩ��'i�K���c�iɚWm��5�H��՚�0J��<�Z*��P`!�<�����녟q��):���M	��,w�R;n`��;�>�k;���ټ���2�� �*�X䂟ٱ��HҴ�s�OAv i���������w�����=;v��	���k�u�o4�8D��Δ�ǧ�2��+�l�#{
ب��L@~�7��"��6�U�jS�$�#iW2�AkΌn��؄��(�Y˞�PE�ؖsKT�+V239�{�p<��(����g?�z���o���[6mF�W(�&'�&ڇv�fp4'���:�u�R1�Z�����u|��_?����N���u��!���by��lbB19�7���yB��ĳk,�oϗh�� ���UK�4�5����u��۶m��n�&��D
N��,選�x�߲��4����&&��jmhz�����a���>��M�/0ߔ%I3��L��2���)f��H�gL'���'@�ڞ�P�l3i��<��S�!F��;r���?�ϟ��������T�� �=
�����&h���i�㎎V�J�lU]C@���d<G����f�����g?�ٟ<��_�^�� _C��%��.���zeתU��?�zn��p�kCQ�)QW�9{��Q\��%�Z~�����ֿ�'�A�D�e�H 賜ɑ����*�P]��эE��,k�C��@@a�Q��)d��$J�dC_O����?����~d�V�_���-���:��^]�\KY��.�����Z��֞\x��p"m�������/��d<FF��0of�����@��S_{(	��:r<�+Cz6��.��f�/(2f(?6�;�bEt�a����o����D�"á����R�6I�Xc A<��<�/��X�g�2U�~�?77;;��e�����ZC}��#�M
օ������iiԗ��.ZM(���?|⛮��0��j�`�.��17;
�O&㍍�sY�:k�G���RA��'��ϰ:}�D[%�y��{�>�!g�
5�T�l���	�P]����c���'�����=z��!���3|���G��K�R� �0
Ŝkۮm�MO65v�	�O��.�ӴM�R;�-�]g�=氧�Eč�<E�p�*ݟ8��/Z��z�%x@��n���>���U�{_��Y�u�SN�(��x���}傋�E8ޔ��I$G�P9�C�_�6��T&��~�xa�
�_Ӧ䆮����������Gy$�x\P{��)nY=>>��'q����3��ě�n��#�nŷ�&��	Yh�g��ؔ�<L:?�b�8�qV*��b,�V7:���������j5QߛH&������˵:�R�im����>�(�Kgo�|j�Vܭq9��>2�&��`�SM��AI�e#tFy����;��LP,��<�=a%��.@��]����A	bY��T]��[.��Z�bְ�-�I�����bP�.�=�"�&�ܦ�*�sxx��������W澭G ��0��C[#���H�u��L�[�����O>���O"���?�b���]�nyllh���"3����W^�*ϕ����}z"ѱl��z��!�%�������X�Ǐ�}�]�- ��.TJVz��z�� <�F#�l�=�/ Zݽ��[o���K.���h�w�ލ���P)�P�8��Y�`�0!]��_u�Y�|��>rh_GGB=�t���U$�rԶC�R��<��@�8�d���p����?��`.p|���Յ�u��Q�Ozd�ů'$[Y\��ob|��)�`e���22:$��`��Ejh�����yN>��e�#�r��%��<�5��
��W��x<�QA�Dq*�{Vc���K/�ǝz�}�J�UyjrҶ輙�**�t`�������z��9��o�5�(�"~�_��_�ƼzM/���a�˹c�/��w�|#V�=���']�>�e����
�:�X�l����}�&�bNƧ˃�������}�{���Ub/�0$8T�j���Y�3 � �\���sE#<��}�L���|���}����tvtPϺUX�F������A��D�Q������Ν;��g `?���7��W������������v�,�Φ �?�S'��.�����13�E�[1��q0�QS~����]l3C�ʲ=��k�X�cv9�R\Bf�������	�^76ձF�Μ�.�'�1�����KԔQ-���,��,'��G�uT&8�/sa�Q���i�p�ڗ�t�����&��q!�0;tv�0�FUZ� �,��AV�F��R��_�z�ʵ��l����=�b�M������'�b#�H��9��� :=FN�s��7m{��B�_��`j��ͷ�5���X�ũ_�5KS���t�?���P�fَu���\#S�Rզf\�ʲ���b���h�Y�S���#V#��j�ɉ�R������y.E} �ϬUj�2�i�yF�t��(0_�v�^�~��ANOOBy��L������Y=2*�ҹ�s�Xb�U�������!�`kT�0I����+�+��8UeB�\�o.z2�Wr���r� ��t/%c��ܴ��~���^P��V����,�n� �Q����'��*�޶֖}2-M1\�R�W�n]ďI���^��b�2�,��mM������e�mM��t�̩��3�T*=:>��#�^z�Ţ]	��HР�������+8ӓھ�N��P�K+��<T�آ�^��.+~ϫ�J2�Diګ���g3�R�͍�X< �f�F���0�Tqꃇ�nm� `��2���J�7��S�O�-��ԭ_�fn|��ӧ�r�2�褊h�����Cxڪ�v+�]*�=������T��kX�ft��Ç���\s�5�������*b�.��zS5��i*h
*w�u�7���
-߼�o�q��*�a����s�pۃ�Ԭ�՝8�������G�Lf�,j�-QU�a�&1�P<m�(4�����|;,��������w�r�-��˷o�65�h���D�X�B�A܃�ʆ-TM������#?�5/ض��g�R*�<��`=,(������YFPd�a�7��G�ec��Y��+ek����%۬�#�3'K����>��'w=J'D��=jh�?}�\<V��:4x��U�9r�.��D���Y���Ra�R,�T�Zݚ��i�͹X���`����Bkx6�R�)�\B�<{�|![B��7�f������?���_|���u�]�}��4654�7�]>r��,,+b�@ q]�P�1[��|]�1�퍽}}f���.��R���)�z�J�X�Y_��΍���ww?�^����⌌V2Y�ܹ�R{�gf�x��I�:#"���<���i
�bj�/?:�ѻ?v����Q�oڌyF�ohs[�dN�$�Ŋ����w&?ֳ�o͚5�_����W}��ge_/	cC��y¨J1ECX�2?����fB�Ю,Q[5m؃uk�o޼y��CTu��J������w���_>|�{���oljJVʥ���C��S�U����X�T=	�=P���S(�-[���B� �"R�Ҋ�	�'��]���Òl��AIO1[2�cŢI^���~@�皙&$�p4&�5��Q)D�h�r(�F��tzptd�����w���g4Eu�����▙�9�����D��_�R��Z����D�etE �u�����>��o}+��5%�LY�l&E��A�h�L�U2�E�R6�Z�S)��~�բ�:W�g�����e=���b��.�z����	�iΦ��$����単^���jo�oc(R
��o����R�]�H=��k�ͣ}�U��W=��x��7��Q��LT4ʇ���da�� ����D�)��B������t���ڭsZ��L�'^�GD���Fa��U��(e�S�p��� �4�j���b����V�L`��j�q�ѣ�{��9���d)'*��0x|V�0��+2�A�+��n�7=�;wn����.�A=�Pg��ް��q�P�x���G@��A��eפ��\�Ӟɰ">�9��N&ṯ[�.!� �&��x��a>TVG�L�#y��L}�+a����d�iqn.�L�C:�{���0��k��	EB�L��+j�|l��{3�=�����\<(-�?�o�>�隫_�Ik���,�߰QX,�����5����D�{~����F�h���~���z���&��ëT+�/��
�Z[k���:{{7l�N�%B�7�8����R�@��"$�`N�[����@��T��9�5\��1�*�\�V&����_�~pp�{>������r�5�P3�sA����Nq��'�ۇ~�  ��:O5��O���R�:=�F��o6�JӪ�:�"'��Gq�M�-^_��j����g�tR�����xkkk pbH �?X8�u�VA%GpRI�����x?v���^����	��'/�5	:��ζx��m:��\�y�y��h�k5�3�i��"@y>ݧ_|��CC#�w�����O|��������6ՠ`rpw�Ll%à�uX�owWϖ����O�s�=hl�g��ݗN�Ь$9)��`u�E:��p�20H�'��� �>�vJ�(���Υ!BO��+������<��C��я}���ˍ�63�D�D��i��#�Ɂ�ݽ=�IBT}������+ �]���6x���z���*�6�l�1ʛ��Y�L���s�����w�Fl���/�˽�}X_�?�03Vwww��-o��+y�.ܲj�l��T
w�$taC��U&���1RK��O�ű�P)��,f&ZWG�!l����K�I��c����''VՅh}v~�   <|������Dⴂ�F	;(����ǆ0��SI�BԤ��(�jR�f횙�قT�p�����sO~���ϧS�ׯ�O��cC���U��O9-�P�w���Jbp�9��N�$��q�
�d�X��?�gϞ�x�mk׬�4SQ����9���� �<r����)\�CWpK*��c�Tni5ƶ|�r��*qF�b�����ߘ|޷��_n�� �PV͈��K-�^�@����m��s�ٹ47�MiH	e�5�/$�Gl�qX�1����L�1eD��P�(�����1?�A��
V�QC��E����|A�& ��^)�tD��E7�R\W
㉸>s����r9�Ԭ?�O����c��O�>M�����A=D<q
Q� ��7j��[;w�l�ŕ��#d�Bi��k����უC������5*�TD����G9&�"�,r��[E���|�R���C�H�A����+U�Y���G��9���Sv����)������sí�]��gΜ1Z�ƨ!Ԋ��65`넖6��������ɕ
Q%`��Z���&#���2����!��/�j�z���W\�z&x!�P���)�J����� /�y�^H!�-=)�h�:xp�e������
�����Lٴ!�:�C���8<Ό�L�$ò���WuܦNi�T�wu�F�7��v���`�5��������Z�����+/�a�Xi˶AJ� qSU���\�Pu>�e��t�A/��W�a}b���$x"F:8�����!�B����e3��3fr�;;ZcuaX�}���Ϟ5��Fד�kHyH؀�Ɩ�����{C��Z=�,y��';v
�2ˆ/cf��b���3K0$cN�L�����ijj�!V���1��ˤR�X�^W��R���=��=v�3�]�}�휫TOa�W�H�����'Z����!��+:|����f����@���K�wUr�~���T��Ө�̫z�.#�zG�c� ��1�\E�6�)�%#We��J��Ec��t:��N��ݩ�Y-������&�ř���ۿ��_���V�^���;���M����C��x㍍MM3ӳ�y�����p(-/+Tq<1���s5L�3��\�h��a���_E�X�}�F�h�G�	���L��U!El%���C췬�7w�=���7�q�}��~���a�N7��������9{�������$�>u��_����nW["�7�R��Z٫U�����.��5�&��@��~R�:�a`0�t�N8ߡ�r�y��/���UkU��u1K���rjftݚ����u1��>���>��+��Q(�ϟ??9=KT�;;�QM٤ �K.����*w�F��j�N�
S���f`�U_�l|5L���ɰ�̒��b+u.����0�f��6�xA���/G�vb�[Q�^�j�oJ������������L��57?�
ś$_;��xs���ohL`6�ލx��v�44p��_����(�M�4�,i�蚈@4�\ ZD��HP�Y�I�9�G l��C� J�"V���e[j����У�<?i��V��N$���O�Nrt�@��ȫk9 kM,3��gg������?��#�W��7��܌��ͣ)�9�/�/��P�:M�-r�oD�O�A8�p�����f��� ���/�g�8�SI�Wtu��G�"��#���3BG�Cg#&ME�3�z�\b\/��G�/D0<�ɼY����aP�i4�;�ĉ	]dE	A:ј��A��۸�|F�|;��͛7���!ǩ�~=[�\���R�@c���n2���f��ʝx��Lt|�
U֯�X�bGD|��p��KVQ�աt�ؾn}<NPC����ہϾcǎhOOz�a��ͷ���O|����mmm���<�\����X��J��5119� ���nP�<��W1wGO[��Yr@C�Oz�󖾸8~�x[��^���)��Ʒ?����[�0c��������4���c���7,��X�"K"?�X!!��y.O�8����ˉ=mQ��˸w���ln����o��0������L�,t����E|��� Ǌ�H�ƞ�͝;s�g�:�T&[\�nbh�>�,�*]�s>W����8�"��1�Ѳ�@�h���3���0ީ�^L���1�E&<ă�Gs� .�"�ZQ�og�Y 'X�D,�kw��i���b�nqi�#�?��*�H�y���� a��@0X�X8+b�>|xjJ0|5*�l(�j�A� �03��7�����{:�fo�Ϸmۆ��w�'�`��^C��gϞ%�z��7�X(h����l==:A�B 2"����!紼����~N���~�>)qE'R���Pu]��L}�cC��կ��/lnj���MK�T���0�'O���/~��o����\9|�$-��#|L&�L�����<��S6n���ݻ��P�*�0i_&B��PtT LL5�a��Ѐr)��/}�N�?|�?�����
��/n�e����s�10~���A�'23�֭8��X�������x=̒�%i.�ȗ��-���p�V�Y\�)�?e/[�FCQh?V3Au�өKzS��CV�f!6�PhӆM�����;8xN�v������<>����ٯ��(Ջ�(��X�c�O|F�������k�o�8;@�V�^�6�l��w�8�h.���7�����r(�kvv,�T�3 ��k}�m��CM,�0�/��w������-�+��kAX�S�֢R~,�2�
;���ƪC@ع\���Q��k���U!�u::��s9b.�A�%J&�s
/`^:Ts����c;�'��O'~��\��V5��mؼ��o~��U��Z��PD�dC]4�}��Bks��X��/䰋c�%�,�zf.��>8��9�����ΗF"aʩ�����<�̋���CAK����*��3W����dE���%׳W�5�!�pD�����ұ���T�}nγ�h(H��pMT�`9�L6���J�z�=�fFF� �����l}<�MS�Z.T�Fbg+�
'(�X�V/c/;'TZ�����S�D�5&�p�DE��k���츖혒8/l��\�U�}u�Xf.��SO7F]0�3	���x�KA���_L"��e���.7�.e����$t,�R�/ӻ��P-!��[Y�ќ�C!�pMݢ�`gX�)�����K�e�h��H���U��}�E,n��F\��|��]�_'!b�B9|��o�J�.b( �pn�7��lx�\}C�Ln�g���5�zY!����sE�!B�Yn:[�D��n� K��3(ҧ,iMH��%��&��|�f��h�[s]�t�,ժ�N �YD�ۖ�`8��$|�?`��"�^��[�����p�$)3(��ԫ���e���9��@u[X�Z�El>��F��[�P�O4$�����-[c�,�r��Q3o����"����J����}�-_�ǻC����+�y���|�p�z{z'��L��Nͬ\��(Y�±X�p��r��I��Ȱ�+M�m�<���'��߸q��S�ڻ�?aW��rM8?4�T|bs�0�Q����,����jx`��G<n��mA�=2t�R����*^u�_�w�u��L�&�e�M0�u�f|ִ��ކDz��/��yY��h����V�D��#�w\|���g&�A�c�/��J�|��~�-���-��̐�p��f����~(�O�<�+�~�_|����'?y���=�2=M=o���]�V�SG�5w�+�V�>ܐ�4�Y��{N��diK�b=��$2v	.	;��?�$*ر.���f�H��D|�1�Q���%�iGa^�C�8�I�Lպ�m]�A0M��Պ��N�y��R�P*\�K����?��'�w�e�!?��4Y%�SU�/��(�LʄE�"�f�y$.w~pl<wcD�*λ,Ԉ"0�M8ˊL:��d�`*U̥�������e�+{z��9551Y�ؔHP=5��"���
VY���?}��&����_�,�m�O���_BQx����bF (��CE�u�Tx9ߩI%��(EB�,e�-"���+�ڽ��-��ӓ�Pe���>v5�a���),럞�`��8�U��(Ì��vxz��P����P��b�h �N��ɤ��d���r��\�7K4#�&,w���Ǥ�>�G\�����hi���fZ��Hޕ�s%,�&�CMWtìցp���%X*U�9�P�IH��9�q�(!O�=CU�677�.��	�4��Cz�Ʉ�_t�PH0, � _,Y��'q�o���+�.{�J�n.�gW�Q��!}�L�Ș�8� �?�J�l�����#iq1�@�w��,>c}o��bqj�5�9�|�|S�ڇj�ȊTIZ)�s���p��f�P��X}�1�ȶ�tKC^n���z�y�,�����j�ՋP�+&�Y'd	Kƛt:g�#<����S�ŲK��7��5c�����uWc�qs��
H#lT�Y��|>f��i�	�kҡ���q�[����</d&��#JŒU�x�*,�uO�y���t�qA�׉�^�T��a{���ET�r�m�z{�<���3)����b~ڊ9�����@�ԡ��*/5g�Ov�����[�"�;}����v����?����r8t�ԛ02�r�ʷ�r�s�=7>>�{G M�N�	?k�7�ᏻ^� �7o���7^���
]���Zt�<Н1��"ͨ�h���s�>x���������G��ɏ��څugp��@��6l� R�;a9Ћ� �1���_%�����#j�PdBRbK���*$��Ň7www�=ۏ��Ǐ!j�����3�@!`�x�Ԯ]{?����'�X���������n�
��oؾ�g���o3�i���^�G�S��;��$z^�qI�����^��^�8����ѣG7n�rm�$�U������Xq��M����?t��q�),"/]�F�06
�r�
bڼ�B���^-������Q"2*� c�E�~�����7�t��u���G�'(����m�.'2��T��=���0m�m]pI����P�5[���V_X��e�)�:���,@��+#l+�����-\Bb8�4˲���\�@���EI�S<��GFL@P)�J�5˞EdϊHIl1ErU�P�,ۆ�W�2��u��&7D窢ɢW)WُpHV����
��!�TNOͤ�fF�6�r��[vQV<�%�c�EU�
-�7\����9�f̖J�������ua)��HD��+֐����U!])���R�G������[���B�[)��F�WBh� K��i3��5(
���S���)B��S��\J0�r�hV��N�)�m���ϟC��k�&2��l^T�#85!���>#=>*�3f)ЅhP��(�ZHP��� �%��h�,�M�Ze��|�P���b;�;�8+�,-PF�4լR�9�v���B%_03�g��
	�L~I��˸��Q�)��X�7�LRT�|����f�KA6o{u-�nh�k�o�1��*H�T���Cpy��2SMZv�ũ2�>���|MY� dCd�=�i/�H<����ˊ�	g�L�-��t���<���.�s�-_�@6|��hQ�v.=SA��r�J8L�4|#�\��&LD;��1@�QS���7b}�E��Rլ��� �����,x0�+U�nR0<�ĦSTl3O���\*�&ȱHL�IC9�#`�v�{>��\��r�D��m2���Y�$��f3���{W�+��m�~���B���\%}�.��Ƨ�gg�����-Y�_��i͛'�"�]�b�IR3�ٚY�}Z-o66%��DL�ĉ	��Բ��NLl�}����T}}����\gbrhx��󗫥���Ф���y놧�y�`�q�������>���O>�$�b�)c����|�}
��e�D�� z�l�����ǅ�x�ZnJ�Q1��[�����a��?�|�X-��"$ s��W�*�_������F"�3�GC�@,���iw+8{�R�)5r��Z���N���=��x0���\�v�3�>�N�֬j��Y���==;�j�ʳgO�575&Ǐ���쌆���*�Fϟ���=k!e������ID!�cu]��Tz�F,��t�� TI<�x�} A�tT��00I����ѧI2ä�Ϛ3M΢��=�a&�d�6c(��Z"��ܙ@hD'IB�~:�Iόn߾���cC�No[C\y�W�����Mq�(�������B��l�+�"nPY��Ȇ�2\��3�ivFȖ�a²�^Ar��m;h�f��F�@H*U��G�������+z���0;�D�[N�1��ͬ��p����O�!v��%Pѝ���Z}�6 ��t��˲����sA��6��CD�I��%8���ONR�e���n4�!����lcw�~ӥ�{5|!^����,?���10z�y�_F�LŽ��zoԈ!�@���Ix����	��2�����2556B\z��>���;w�[��}?���i[z�νHq.2\�c����8B��^q�:h����>wl��d
�AV��Q�ɡ�A�]�1`��?��/lٲ b�ޭ�\{�׃?����O��*eAT�����9��6&G`�y9G��'�7�1����1dA-�%�L���)/]�Pm��q�Y��-�"�e&5D��Sx��ҙs�
t�B�*Ȥ�x���P"�-9*~U����#��vuu�b��&�(�d�.�
�f��{��[n�ڼ#�V!#"2������e�{9��M,�NfƟ� <?G���ď�n���4�#��*<�N���������2y�Z�+��y6�nOS�D���av5à|5#�������"�a�b�%fx������cl��:�sb���/߾T��W�6W��U{��m<3F��v�G4#M����gP�4b�@�G$=����ˀ�r�o_3�{���o�g�%"nd�{�M�����7N���������+�
�v�+��y��>o�O�g�Ԥ��g�I��8!G�`��'}�����Ƅw��*z�iF��9TӀ�+&_�����F���������g�;��'N����<��{�������W�^\�4Mn޼	���W�
�1��ҥK������� ^�x$� `��B�ΝOSFL�l&<7�p؉��(X1l�Φ��,U����S��ݝ���~�Uo�]2��oPW�)�Bi���>�#]X?�4���͎���@�
�����>�N���g���a�����sϽ��+����[p��ˉ�l@u�=O>�$�r�Ɲ����G�h�E�H0^�ɞ[�h��`+0��#:�J=���9��U_?���|}Q4�翗�R��l���A���8�n�F�=~g���{��{���2��6w�;v(�mn�����[�>����)����,�%NC�ܒ�"�_�MFL�-�~�O#�#��/~�O=�J���	r�������?���EV
"��v�n�e@���� ����h}T��r3�#��Z��+��j�tὬ0��k�B�"NBnG�^>x�h�Mza��t�S���WC��Dw�Yw0~���ޒ��)�)�Vl��}��$�A]��I����Zm<�V�6�n͘x���ZCZ�����`c��6�vE�eZ������W?�����g��X]x���姾w�Զ@x���o�O�HE��?�>}�7y�쩅���[�����4	8�e؜L�Lľ��Zfb�0�@�7�2n��!�$���؟x����_��`��y�}����ꫧ=�3?�3����n�ĉ���=��t�n k��&��"�Vk`膓F�i:bg�?�ʤ��JS��'$u׈Ԩ�+4)+�D�N90y�%��1xo��4;�^�����+
|���MΌl�8
�v�&�X��UG*�|u�L�C�I�n�5kIn���x܈�]ό�9�Z$s�i��VH"�������i�u�RC�,��?��ӤF�'�G�Qj+��`�M�'ڲ��N��Lj�$��>x��4�_�-����U�p3�3��Օ$o�yA�9)�(+5�����Ī?�b�XL�F����p~���q$@���!�U���Y"�HQ}p��v?Ś�Un�,���c�?6\i��j��E��MiX�π��4���4�"҆Dͨ��4e�ǧ�� �|p�RE�a������c�P7yJ&kG��a�'��q�����������t��<�G�v:3��<oBd ���dZr<�g�KS�7�}�>�x r@��:u
D<�r����c����g>~�׾�׸N����i�q2��Ϝ9��;�.�S�:v�$�.u��77�]�]Xp�|���J�5��:ƙ���O$5��������Kb�)T>�}{sO��\{	N3D�m����[}��ُꓭZ�������͍4S��I�8mv����|���&��^\��9d�V� ,�(��+++@`?����ѣ���r͙{po���ɹ�o�ݷ��V��)���u�w��� 4�v��1x�՛w����"�YJ�'ؔ+Krm�m��Z TR
�8�'�0i���\��E��I��`��!'pHfQM�"���O*�;%��,#��z�M����T��~�ҥs���C������g,�	F~ww�a���|D^wö�#�`���p�H����@Ww#�0�%�cq�Af��O����M��4_���[ƚ���!p�@��Aoq��d��93��z�a�-�>W���N��{�ojsa�{j�\�W���}����z�-l6i��GO���h}t�u�b����+o�D�ZK�Yj��XS�p4̊MrA�B� �d,.�P��5���!�L���G=D��lhO3I4ϱs�B��<�t-�� =����Hj*þj<` §��{�@:\�v�g�g��"#��>s� �l���IEa+�W�~�!�WQ�]��e:e^�P���c���4�R�HhP+<o�,�c[]�3g@�����)�×���'��-��n�Ѐ>�^�+�a�Q1�xC�r���xƳ����&����U�bTܙ$����_ָ�ގ��.*C٭K��|�Mx�x����A5�e��v�y/���쓉Ŀ�sQ+	֗����=�E%TP����V��Z��S _�����ٓ:��e�Q*�9��L���/�Z��
ʦp��dz�m�8x�����xR �w�V��,N0�T�n�s�h�D Y63 �5-)������8`���3����9Ҁ���nccC��'�#,G������V����鳼�����X��,	��$�:���5�n@��H	x��y�Y[A�̈́�oR��.q�� aW�a��5���S��3���'�'��q��X���۷wq��������!O"�s���_{����k8}`n��̔+{��� � �:��`���p&1=iٺ��b�q��8&�v,X܈���޻{��)��:]�b�s��U�~Q��q@�5���p���mb��sƟ��g���o�c �^Y��x��;w����˿������3_��$ܮ_�>�`T��������<¬�䰽�m�i�>�n� ���l�i�0���9l�@ޥS����b/���Z�&:f����X1=��_������ao�0�� ���&�Q�_B^C@~��d�����\�Ѵ����Ҍ���݃ ��`���;vv��\u��+�e%�Σ�"ܸ��oumu@=ALW��#����*�Z>��E��50d@�alئk�Qo�U��o���Wřhl�Z$Π7Vh�[�P-M"ʹ�o�����ԥq�Q���9�5ӹ5ˬ'id��-D��)��!��ңTno���<�"p
;�8��&Yd��(l��M�%�֭�WvVE�:�t��y�;� ���e�4���_[v[�M���pP��N���E������i��cs��������z�I:���ol϶�y{�=�U�Dۉ1�(B���GF���$pM�gLz��^h��x<�2�r�8��>3�ꍻ"L:n���:�*��o\�s��c"�;�hy�����!�u�{��Ω�ſ���=0�V:"nò�\�����j95�����ѣG� ��X�	F��������fuc�Mx�~<v��Z�$^�_��=z�ؕ+W�AQ�N�0{�Z����`�g؍�)=�h��2�`��Z.���|�_�j'�N�A
o��A�&8
"63��c��������M$T��pNQ�۳M߫��^7,�"�ո{g�Q�B�����J}
��HB#KS%����	����d8!�vp�e�Q�a�PHoSo�-��*3J�vfz}p���dog�6�U��xQ`F�=�����-���Q�K�D��V�g�����Ro2e��@��W����S=��r��6B�?2�l��u��Z2[G��Q�Tld�q��ت���h�54��Y��)�=����y�뙗�Ify�,eYIb�>�f+�QD8��nQ�C"��Uܙ�M6��%�A����Pș�ԅ!��K"�l��MW%��B�'���~�h.�d�uZ�
��݃};}�,<;��c��F��3�_�z�����c'ff�0N�T֠�I�˖R;{J-���6N�i�a������F� CW ����tԭ�G�0����Y�s�i�ּ٪7�EK�0�
=����c`y�lʮ���<*i��4��C��1σ�z�vN:=bvj�;����O��ԭ�׸��t�W��U�D�D��'��?=d�J�ݻ�	�|0z���_���]���D>G��(�qf�+Wnߺw���g��^{�k�ݻK�b?�VN_]�i;�N8����g���&�A��7�L�������1�}c�Z��L��������PMk;�@��sM�^�|]Pax��guZU'�.�p:E�v¶R��5%!Ԃm�Sx��N>�a����=5 v�]Jp^�f��H� 8P�2�ЋL-��/p@�	�#��F����.#STɠ�u�`�G��_S�ؤ�h`��q�h���"i2N�ˮ��[�x�����x,l+�B4�h٩���8;@�h>RwF3����2u;�]�|�ر� ��w�Φgi���T��y4N��c�������6kU��9MU��`ƂRN �}D��5D+��������
�xX��4��)�w�T�1L�����e�O\@}�VQx�&�j�p����ͮ�'�_F����J�^vݮ녷���}v渟���D����{1P���,�r����:-��E� ��A(Ak�� }�i{��s�̲ Lr
ٛ�]���TA T��*_�r8�p*�f}�"4�Z"W�"�OV�:��Il�#.H�XŁ�;p4�R����X|�&�40R2;�~!?�,�����[�!/�����h���|^�sŠ��i�Q�$iV���t"�u��������ZQ����_�鰲Z�fĵ<��S�Y��`O�Օ����0�� y�#[ý��ϵ���L*�{i>"q�ӇW�T{�������{�9+OS�Ұ�Ȗ��{I�ă���/�ñF1��u���M󠀢j�8��]R=<�3|v���r�����T����P������'N��w��I���8�ڋX���B��*\B�54<M�M���8MY�>���[��A�e�����S���R��.0S0%K��� o��8$���Lf߸�C�}�6w��E�q/�k��������e��������9OZ:/�d�� ۀ�:i��P�q,/��;�Z���}�$�e6�u0{b����#��f��@Q�ǁďr��@ �����PY2Ŗǫ0oH%5e4�~�.9=�\_?�xbzp:	=Y���b)���R��#�#��QLUN��X�q�!p�fp1���!���q@��"ZVM�?��Skk�"�����s�K�`on*�Z��a�|j?�)�$ź�������� �o���3�tG�=D�&�c��(����`�j5P�R�������OHv�M2|�� Aɍu��BJ�;/����Է1s\w�ȭ�p��ȝ~��By�Ŭ�~�Q���Ta�rBP��v��G�@ ��8�|�1��ɳ�COd���O}���ŚfX	.&-9�@�K+[M�tQ�1����~?6Y�I�r�z#onf�ԭ��u ��V������֓�s����7Љ�>������{O�i��2�G@Y���|�<}��=�A�3-Q)1tx3f�����7�푢�	0"�*�N��
(���5d́�Qex2Ȣ��F2�w��n���KNdg6
�ig�)x=����,�Q������6��;v�딅�#l�˕���5p�c�����TxJ`H�_��5lQ�sn�֡�Y�O!�����@E��d�ý�2#F&�y+�+��*�1|'XaH��#��/s�:��Q"I��bP�$���y�RHE�C�S�]V+O�O���V�W]��r����=�F�K��Z! ����bz6DE7 �Y<8��1�i���љl+�Ȅ9��K�������'KL��`m�e�\�5�������~���gJ1>++�$�ٸd灷�J�P�c�x�)�b�ϲ(�x�rW)����ԞFǥ�s��m~~�ִ�j�R�kX]]Q̸����\4=h�O~�`�o�3��N��� �ޏ��(�pnYj�n���PG(��I��'^4~Z��w�m�M$Cj9�f�vF� M=��?�c��m}�}tRz��*Wέd�rq�F��\��[7�A��n��������*5C�.��@Q��Z�Y�aA��}�h���a����TZ&�;�6��L�@.Ĥ�(0�L�b����}��rv�U'L��>R�H*�|ńw����-�.m�^��������gČ*p���zU�3{ �;��K>�Q69�5�����я~�o^�&���d��RB�cݜ�I�j_᯶�3�׼N�r��ڠ9Ğ�Ƹm`������d������a_�g{��$8}`ϵ�5�^.j�W��D�'�জB{�*�َ�o@���au`�#�Pu�(���R�l�,*B�M4�ִ���� ����GW��Y�t�҄ҷ�����2A 2c0Bk�n�!X��(;L�˅�����=�\����&j�Fh��"9��Ԃ5�����g�X���"W���W�PPF�fp���.����[н�(��_��ߔ�N`�\�1��T���6�\�a�v�2cAP:I�ư��Y
�\�N�؛�oZѥ-�����w�F顂�A1#!`K���hp��,e�#���A�sYoF3ӸB�ݢ�����Z������X�U�h��y��S�O@�#�C�)��ʯ�֣��Ur#��_?W�i~F%��1q���
�ݙ1�����K���5O�ҳ�n ��7���(]���j��`�XH�\�S�#���g�NF��FN�#���#߻w�����%�׿���s������<�QAeї�V/\��9 ���C��h���Ã����WN �;ux��1ٯ��[W��D�kQ�����v0D鷰x�{���'>�	p� O�E��b�N��_na� <�M�@��1%ΰ[Sװ�V�&�=@��|�<҆�P<�5��2~Xu?�(�@b|R�y�-�����P�"��b�n���\ӂ�"zWĮ�6L3����uE(az�ʨr��A��)I�~�c�}�Q��u�MO,�oR���xU}��TS��
��;��ۏ��h��X����� B�3=��3Q�)�����h�k���SaKIB�uN�>}���������v��^\X���{w�`h+�T�}8���'c�Bӂ�G���!#.�P�. ���ayݞ�D�?ۦ�v�����ollBI������z�*#��{�Cˬ��H��̜fX�1�U^荆�$�A�����6X�v�ڭ�Wo^}�V艻k���8��ȵ~>wL�da
���G���QmQl�>~�t�b`)u&���~wp���Ax��=۪Im4���ec�P�&y"Ng~ٲ� 1�N�&ҩ���tf��{sx,n޾����ñ�}�A c�O��X�9.xՊ2bЪB��it�j&�\:~�fye���>�|�{	d�Xf��CKby��U��z��k�Ñ��br���5ሑ8H|/44��y�Sm��32 � "g�a�g��ے��6$�XE!��Tߒ�4_��TkHsQ��ȵ],7A�75Iބ��9�'�G��Q��yl��a���ߗۊ����4	��{&4I�4AX닲-Р��<R�J&�����s?�>�_���G>S>t�xE��3�X	u=6,��&�c[��`F�����)��b4!Δ�"^M�Q���M62�ޘA$�X���Xp,ʨ '�U
\������vZ�i�	D�ܮ�=n��m�4��f�F�n����fkFT,H�W���[q$�A�s`��zq�"�Q���MM�/)�/z:��+�^>ތb��f��;,NÓ�e��������l~�~��������Q�9�-Ӥq���%h�L�$4<��hMT!z����U*L�pⷛu�2]e�b�\�T�</�s�un:Xup�(���xc+�U�[5}������?y8Nc��BK>���dr�XV
��[�dJ�3)u�$)կP-0(*�b���?)Ÿ�l��
UDm�� g(@FGX�u�d���̼��k��ޓO>���B>�A�{hZ-��a)QZ�b����,����������[�Us��k���H�	�ε�F�=��2���	��×�����o޼	"<W.&Jb���'�=�`={8�U�_x�e��b�f�O�g�����ܘ�>Z������(B�^2l�v��Qy<}��,]�$t,��9� �X?���'��v4�sT�Ea˪V%i�\�`�P�O��w21���㕘^���K1�/�!�|A���|�2�}��ކ�b*�~��^x���hh�X�sB��/�,�,����i�;�].�eG!�3rE%[�c���!5F���a���3�8q����.oZ�}`V��O�OX1=5,���{Bt���M+��O�#��R#�(���*&ݜ��Aףp0t�0���S�Y�����%��DH��y��G8u�gZ;3�)�`�6\H�= ��T�����a8�&֊f��wmzFD�iB8�Z����EJ���C�ǧ�q��t���#��e���CPz�a����,�	}a;)�sk)��L�r5�Q�.�؃V4���$�K�~�_FkԡK��2��BeC�ߌ���fpL��o~�<w����?S��T��_�s�E���q*�~r�����fT�=��m���Z�)7�\^PZ!e�^4�1�&;��O`P�7n���w�{��œ'O���;���=)&=� ��� '���q�4&���3�0ě�!Vw�h��;�*�BX��"񇼘��6�h�9vI�lL�֯�n��7��^Y\C�9=�������j�V�s�Cb�P&�E8]�41�R��${hbr�Wyjl���<y�[�5��"�;|�%a��k�o�i��ˏ|���7n�f�iﱡ@��l"~l��Z]jc_^���y�v��	�	�s��BI�Ͱ+	~����[�I:mݫ齽.����hyy�z��'.<�v��8w�2��V]��b�0�Vp6�k�APͰ� љr>�ӄ"vq8��vk��p��P�8�5�Epu-Ό�8K��бS��l�%��� S=;��N����8�ŽQ|��V��������&��L��]ϱ��b���_p��T�!�I����!r�������D�%6��,/DI�E�����j��Y�G�6�cIÍR�ҍ;o_��B���Ƞ }/�鏝fc�;R����+,�+0f��#�߁�`��.��qS�����Ǭ�r�BE�Y"��J��{4��YK�f*�(S�̰��Y7��/G)<�L	1'h�R���堫�n7��KP��x�"�:4�hD(�gƙ��(|� i���Fa�,�厵)�0��'��*�Nɋ�	44b�����D�=3�a��{��B���)8hUc,!<ʀ�A3��'a
$�����]���%^R'���=]��*�~�(�=l5u����1��J���� e9�Լ1��9r��<amQ��ҷ�a�
���W�r��H����,@Y�S�;�����9�~YY���=�G���� ��b���?x��֭[8}��ey��Ya�Vs
�����4�.��R�=04�2U��h���hL�F�)�jug�gEU5�_&� ��l�������F�`�|�+_�����_��_e:�7������Np &#lJ]L�!d [��^�dLL�a사�Ђ�S_'R�vu8Z�X�/U�$�O�`_��u�.�B����#D��es���22�y]K����6�"�1��d��BnҢ8MB���Ev°���dO�͚�_��d��p@-�'�֪�7#�Gh�V��\x4�)DT��#�>]��޹�y����O�M�Z㡛�^Z��E~������*-$^�&-���pp�s�M�`���n��w�Ǡ�����)j�M��:Ɛ�%�GE����&�p�?�����~�:�|z��P,=��AP��R�diR5j���e�8s��t8,�������5*�ERw,�N;#8?��M�'�<,�F�0�6��/�}f��h�܎�-���{�r�hZ��+6�Y��(â�v�('��Ҥ�d,���ظs��0��`�g�У�r�g�(��C#�p؟>����(��&!'����~�ܳ�Wm��X�*���H�܄'⾎�)�;��5՟,yB�4���|8����<�?$��$}*��G�E^�j���/'�i�D���,��*��0�)2���OT��g��v���(���]��n0� ��d�_)�X2I��v:i�nƾ8�J��y8���iF�KI{������~��iO�T^�N�n;qj��X�����83ܶ�zV�&� ���ԯ�U��9�Pfy��3��uj�:�b�zXjYRz��u}vuX��L>_V���ua�2R�2��s��������:�=b��q`aY�Ä���!ƔJ˒�R��B����^�X��
a=lb2X!N<�4w�>{��k�A��=�cg1Eh8�"�Lo2�)B�"O�Vi����xB����NђX�!F�O[���S.�ש�'��k@�gJ�[�?�*�N�znY��#�WY�@�w��f�^'Q�GGxnHՖ:@<L�["r�(�/W���C�2�W�E)��q���1	Xܑgs��)��[e�r��M�;�iv����4��a;�^Z�aǴŕ���N�*H�D��<���'�ʨ
���{+KM&_���+�,ʳ�� ��f^�2�ÒBm� 8�|�̙3�e7n܂���~wox{sʹ������߽^w�B�*��&��sI:�\�L�\E���l�N~,�L�ƭم�߼�7�5G���V�ȉ�����ѓ�&��}ϩך�Y+��'���ua4�ԼtSZ��[��s5=��zsn��`�8�	��FA��/���������H ����f/����l4���6�@�5��$�~����Y���'�?����έ;kJ�[���O�C�Vmv~y��;~�����{2���cq���O~敵��;�?��V���0��$�6��� �<hNA�C;�d4Fè7��#����F�J���9��)a��eG��:�)Ə�7�=��㏝�{]��n8��*��N~8A$h��<���hB����X��z@Bp3u������=3-��!�t)|o8���I3�m����4v�F�Л���H禘N�5��/
^ecx� �Q�n��b�l,j�Ē"f�k�r����-��s�3�NK�α	E�S�F�YT��qGh@VBlx�f�N��>�e�'��̢�;���K��;1����Ik��jU�i�y%��8�=qo��L$�)�)��In%Ɓ677_���o��=��痖�9"l/t��l+� p�m��Ӥ�kv�˲Vn޼	��a���6�+"�ą�R�VR��|#�b��i=�Hp�"
ӄ!!��(�:�|�2h,�JC��
�p5 #$~���}�7pJ2e��u�P�:����׾��<Ch<�R�#�5�;�����5��>D�Xa�"d˛�t�8ƆK�U(e�
�l=oI�z&n�����?��L��_��R���s75>�5c�p���3#����h �6Uq���[�(;c� �8�1�V�m��
ΉOV/õy�^�Ȍb��U�Jz$���`7J�xS�~����������x�B�qRZE�义IaI��6AP&aJ|���u���v��M�6~-X�9��� 9�����3L��Q����[Z:�`` �K�%$ǇE���˾9,e�r$���&�c��9ә�g��l4�W>���^}���tZ���?B�^��d^�nvއ�Wi��v�c����KKK�\�f�!���|���
�!��E�s��Wլ�����q��D4��`X�E�9���E�(��$��t����%󃸆݇�J�{�y�w�@�'���� 6b�����+��(o�4֏
���2<\�q��Q�-�ŕ�����*-��m�	"��n��nF�AYѮ���B�*��E$��6&����:6DY�Y)iEвjx���}Z�]�����:@?UyD\�_��M1�]�=z�ԩS �o�@���]I	��{�ZYc�M#�����
d���ɦER�J�W)�5������4��)h1Up�lo�rG�M�!i(I��Z����%��u���_gr����<*SlYQ��[*������,��+���"Z��S�ߊ=�h�G�U���)��������}�;�X9z8��N=�ȅ���ѻ��H��4U��e[1�^8�q�2�={)�*̚�)�Np=������?+�����\��x����}�{�O��~�ĉK�.��?�?��F�yF���(f2��%7��Ǿ�o�΂Z&?��'�߹�������s���$-H<خ[�n�N���_��?嘁(��)Q*z)���W��)���T2S�$�T��
��"��P�?ܕR�V����h�MCY��P�s8�#�[�z��/��^�'*��.��"�7eK7C��A X�q�G�W��x�?��?�uG@{�;����|���Gj}�+hh�Ww���{��������H���mj��(�j����t��[[�{��Vښ��#���2kh��3;�|�}��c��FE��)։��"i4�øP,����.��B��nIӉ3�ӝ�n�=�y�X]��BOwj�c�7N� Na 5�%M�8
bP�{�����0R�T\[����&!p�j���ՙYl���VaD?�LC�K�`�E	6�`P�#!��.��R�@�m�G�{�啥PZ���j��RLb�V3?��|�p,�f����(Bŉ0����KG^Ikw/���5D?�ހU�K���V$�y���^a�hR$p\`V�[J?�od��GUfLqy?�;	ma/�tN/-64y�Q��IϠĜ�5�x�HAT6\�A�kl�U��3�䔥+��`9�^��c�PM:-�d��� �Њ��f俒O^TS����t���	��"�_�/%�y��`�p[�aws@V���Qq6h6�o9�DK���@�VA*��,|+���ɸ��o*i�Zi���W͛h���+�7����=	���>��?��mՖ���yn"�0S=�Ϫ��EZaz�8Eu�뇛��<B&�.�g;d/[إ�#��>�Z
=ٜ
);MDE���8;~E���ԕ_�=8$����G�|���g�y����_�wa�?C�#�,]��HEz���47��A�c䏬OP� -���Pu~Z��Q�`��@H�A�^���Quk�6��n@X�7����,�:��ڼh��#K�U���)d���5gWI8t��Ѐ.-��B��:;7���j���Dݩ�����TE��%i��I��y�.�Ui��[n��9�/�TU"�c����<����#µ/8- Wy��"����<Q%��,��X�J&�A�9�?�q#%���]��\y���u@Ö�[�pV�3�l�$�%�#����P��u�Y��,��ǣ�L����/�z Z���ml�����6p�� �<����ĭ2��7�8�U�;�=���lpім�"�B�+�6�ȇ{��A�p�����(��G�� ��`�z���Gz���gl
���9~b���O
(�d?�?���c�4����zZ����;�4����Ҧ!s����+�݂nDQv$��(>O��_�4�d��AH�ٲ��Ic���aQQ�et��G�~?����ا�<=8��`�O���%��>�n��4�ʨ�ƥ)"ع�{�\i1�B���e��h�6�5�$���o���� 
��7�x)x%@W-㩃�I����L�e_X{_oc촆��M݆dl��~�ݴ	ͯ��9��FH�P�Ib����v������bu~�d��zU����|~UZn����O%�0L��i��?����҇^�X[��<���N�J��qy̿�K��9ʺ�T9�>��!�KS�Y>�X�ZNtaɱ����שȓC*�9�@���_e"����T7�K
`m��=
4���o?��SO>�$���:߸q�,�8l�������t���~�ӟ��׿�h^)+�|Ě��*�!Y�qK���r�
�5σ���w��/}	�	b�mNhT1����.s�j�"������%�6���)� :/F�ӷ�:� *�/mw��˟���_�NÒ�(_��8�1��4���(m��MI�f՟�++�i
�˕����
��:G���$�h9��2 ��3�0C�<�}T��X��۷o�V/���K���@M��߻�m/����
��o�z��7����?nlP�\�ܹs[{���;��']7����r����9�u�~RD�aLT�!�&gN�G_�#�!4��!5g:�'D�m���RMn��4�>���խݾo�G`�&��!nR�j-��6L�j�be�<��bq���v7a��p�߼����A40N�>�@O�c���q���=�B�n��r�1ƌ`6��6���N�F�q�evc�~����i�aᨏ��뎛G%h���<D���e��X�0m��Xl��@:�CX-�P�f">�I��i��$Q�>�N�"%G�/b�����M��T��^a���긧�;qzE�Tg��h�
;�u����7�4�����ǌ�is���hAG&��.�?�z=�M"�k����i!g͕+MAK�OQ1<h}��$�,���m�\�V�9�;T�԰�5��	%�!�*�A`�5���\��>I.I@���l�¢�혶�N�>�Spe*Ĵ>��x^g��3)�Z�������O�oL�C�������c�?X����y�ß ����)q�eJ
�D)8�Rf��חE�*�&`���F�Vi�R^FT_{I@/ԙmI�������kuhs/;XZ�X�<�����_�M!B΄N�ZPR�;�j�s�~�C������	pu��]6��3l�QL��r�ڨ܀�@/=*�� j�c��Jw_����+�tզqqa�Q#'t=x� ;�5�R��N��ʑ#GΟ?�����AYK!]���^��cū�RB�g��r��� �h��wDV�0��0�0���(�c�E���ꪠ��^��R����E`3A��>���̱E�O�rE�l��*�>y���g�8Z�:���G?�ά,��,Z��!���i	
?`��01s<J������T=��I��I�j�rI�U�i_�afvv�ԩS�����ѧ�T�J���<�QaMc��}�������K���Ѝf_���4d�w?y�u�.E�{9Oa�2e��&p��3Gñ~ǀ�r�AdT d��6�.F�殔Pli�֙3giev�5*�������QGFE�@"#�2��
�&dg��3���~0�_x���Gk���UF��'酢��R`<�"s���r�x�F!�5,R\WXD��yw`o���@�2�>PR�֒�5��3�?[�&�6K�,U���b�����1O[�e��x�8� n�O��1.pk�;�9��~�[�4ϗ;���ZU
,"(��8dֲ�&M���$�Q��H�p}r���2gS��n�$��P ��4l��U�������zq�q�$��U�+S��o��^�� ��}y�	���0luc��H�\LP6pIq(��W�>pU��#��U]QT{�C>�kR�
��=��Y�5_�~��_�h�p�p��(@5�������l�М�= ?�!b��e���g�nQ+,đ�Pl��ӳ��I����x�1�Wd��k8��E�s\;��[o���W>���+?��`�sss{�A���x�9\�rN�>�� N��G?����/���y(n�qP������A ��&Nv�!�16�_�r>hX��O?������^ɢ?�\�Wa;�d���r�%QT���~�זk�C�%��H��20Zc�����8��:�9#a�r�����\P��
x.�rM�]�u��,�g7�\)dپ!	i�*�O�lA5=,��V,
�TM�q_q�S*�wݹ}�O�{���D���!��gʲL�bv�½��Q/X�ѣGW巵�cv��8�� �7Ⰱ(��`�X��l=�]U8�(/�rl��1���[-���os����C��&����qVoRo�b�1��ۭ)��)΀{������86w;��`��{�W�l��� �?�GIíGC4&Q2
�k�X~?H�g2J�|
����[�V��}?���ּ�~�P�cYN�d���V���N���-����I��4��ճ�1p����&##��.
ůc�4�Tja&��!��~�%h|�����2�f�s{�'I*�7�t�}��:�
�\��?-f	��3t�v��8���^��Q:ޙ��qd%��:~���,� �jc����DD
r��-��wo��S��$�?���.��P��L[�W���9��T����E�V ���2DyZ���CMH��M�&h���q,�[h������,�ߔ�ѹt��>�o�W��*�E���B�J��د�Jpe^-Y�S�-d_��Y����EAx���_�`�GN�bGp�s���n"�H)�~�*2��ԩ��+(���fJ�;��-�B��󥢁��0�%;�ml������S���[��Y�:��N���?�8��0N�
,W��]ޡ��Ir��m+�G�Y�M��Z�|�x�y��}�s��;�����p9@f>�|�?�/@��2�-i/鳼	����͛�DZQ�W�6ÄWB���*x�m&�F���pbe�b4��N����$O碩z�[[�@��1�����S����~OL~�t�|<� ˋ����/H��^��OѝTq= 
���r�������\P�s�_�Oc�9��B�~�����2k^�M��T��h 8�mZ<�X�kB���z�幦��ӧh���W��ׯ^�D���0�g-S#ؓGf�h6�����W?���u��i߆���Ä#`�;C�1��p��t�ڔSBV�_���p�����,�,oZ�%帛̴̇�Ԣ��r�hS$u�3��:�0�x�#(l�:������qnf�nЫl܀f$C(Ǎ�E�ɘ𱹥�c�]:�뗺��~E~6he����(d�[D*�N��*�]s��g�&bkGҼ,xz�`DR1����#�O�)�pZ�pA@�*ܰ�Ϯ:���1�.T��7�+`�M�8�4<x�g�´0��(�L�Jh}�8d)sF��P%�	f�M��g��/�)��a�J���^��J��J_ވ�}�!-�m;���h~�$�R�D��N�D��4��^�c�+�#�*%Ĥ�s�B��K����#��l[�?�b��a<<�¾0ȝ �\�F�M���
�@����lPW�e�� yg������KW^&2��c4��z��K�����Q�h�#"TUB���*娇�
�;[�`p.,,p1
|vkk�����	��W��������r�(w/��N��ˋ�_��Woܸu��;��U��Zo���/�/n�&�<,A��O�m,0S�~�1Qx���A�Q����J0XI�����%� �ZX�S�)���:���*9�,��P��+?Ƞ�iX�wU��TU`��"WN1!g"�����Y�?�J_�*����fuǪR��$�p��E�L�hρ�Ad�6���[.�z�q]�t���S,��{�fl��76���4���\�[Pkֽ�{���>��O ��Ȩ�Op��4�~׈ ݚkX����?���cǎZH�%�?���=�0k6����3�<3� ���{���FS4���8�8LM'���^/&>W^wg��sZO��,�����s��I0��w����ĩ�{���ݞI۲�1f�v+*6��$i�����G~p뾜[ڊe�17�0\����̫�;�0��Y�ϯ��ƥ��$R�0ZvgЛx��tY�{�l,E�i��>A�q�{�ʃ�����u?6�Be)R �f�Z&�����H�$�,�n�ܞ�;�xo��Q����B�3J2��t죳3g8ά������p��n�O"%V��>�بST�� Ik����]����Tln���<�~cթ5�����n�M�ֽ��p��x������ݑ���E������׮\Z>u�����i���jX}/h��Pa���p~��~�ԇ\�J���&��>�Բ@�4�F�`����2f:�{����{z�"�o�D
�<� ]�`R��9CMn���x�����*2��޶1��ڭ�ih�xd 9�	ʶ�$���R#>F $5�#���~�"�1�Tc�'�95B���d�r%ű� O1�E y�f ���RS�Á��s6�x�}0�b!��wkV�i�J�9�j�c�FM���̛ ��&c��a�k2L�̏p��zo0��cs��i��8��b���e�B�i
�B�9&�+����74p�d�]'�-=vc�MiL2�k`���LǞs��Z�fܹsgiv�,G��S�'�Aok�Q1��W6G��p�4<n)p�"���"��0�sJ1b�*)e��+�J��0�l��Gf����-�}��`^Ǆ����"�"�A;qD���7 #�q�;[�46m]��������lۚo6{�}�ڋW#����1`��Y�Ċ*xM��I���SB1�3 �,V����w0�&����5�l/��Bu���3+�q��������f˪/,������u����W��p��7n��������Ko�>u�<P���1Q��5"�YI�^��Ӓ�E�a�
D�?�b0���ghd�crAi�h��`�4j�Cܪ��}�'Ϟ��ƶ�¾�50[�ێ���=u��Ŀ����}����6i���}��k&8�F�\����G�״|��#�mͰ-i�i�[Mk�<u<�O2n����HEH���b-3�(�����۝V��^U�f}�!EH� �jQ�ұgJ�Tn���|�=�㏵�Z�v���8J�0�5^y;}?�R�Е�Y�4�*ޤ�!�^����e	k��ͽ�fgFj7âxl&C:�mj0�'���%���f�2��q�̴��g΀��sa��#c$��{�A��/���;��p���z����8����}�3���>ܽ�5���Px`EIG8gS����8ˁď}�c��~�����Q�TA�;" ���R�F�}��)ݰ666������W^y��.^��V#��>-7���\�b�
�����KU�<sOR�;�@(쯬�n��ϳȑ ���0cMR�,��"�>�C�8LI��
��7��=\v�vf;�B�l��o�gAh~���?2��n/�t���>���Us��G�R�;X]HC����3���p:sǎτ�����a�@�/�H>U�$`o]|�Rob^?MAxa���"܎G>?��w��k�������^��G>��}����𧙙x�y�ܹ���7K��j�2���ښc��!_g�s���K��%lK���k���-�
�����[9��03���~^E�c�����^��G���< 0����:�C���޿(�w��pNd/�VVVB��n߆}^j����8D�R�Gk��%���!�������q�(R�L�`��Y����^J���'=*Hȿp�y�d�yfQ!�����:����9~��؂��!��ţ (aq�,x�X��y��l)Mr���r)��cJ��A��}�[�3D|�y�Z'L
�a�e4)8r��*^\\|m���g���DpD��aĽ������)�R*�}Sj�J;3�D�[�ҍ���T�_�3N�>�M��^w����A4!���I��I߰ENX�5Ca���25d��KKK�ΥX�k`�4?KT3L�X��5M�ӡ2��"�FZ�ŅU�����\ю�)���+%��j���F�0��1�Ս[�0
k9�&<��8-WE�#��TTX@�kE�n�L�h��Bw*j1�e��"��Ӥ>�ľZp�b�P�N)�9��N�m�4)Ӵ��8���0F�Mk'�,P�)ʒ��;Ev��T�+������ED��?9��@I��V��$��r��}�f�t@Z������oo������r�\v�Ɏ���;Pocor�ڕO=#��隣?����xw��d2�7�Z�����ʬn�F�����.\|���>Aȝ�x��l��p�N�_
$] ���,Ӱ�X���]{����R�������~�7^z�S���B�>��́Ϟ|f�u�֭���Mwv��Q0�8ފ��7
bLrgݡ7��ٹ��f��2L'Jb�BV"x[1����A�N�(��8J���sl-,�����q&g;��+价n&��^��2�h�-�+�֒Y�%�����`B�?���;�����Ο?������՘�uG3�$EG��:��L3��;���<H0��[;{����^s���x�R�):������i�3���#/�k6h�Ս�a"�Qp:��p ������ �<y��x4~����~����O��wΝ=���Ad۵f���ݽ|�F^{(n��w��hqS�i�UK�'���՚��^>@bggh��i�\�"�PXY���q�i�ou�~Vk͂�d���lO�I���V@2��ݻ�ؚMԝq5ڋx^[sƞPh��)�Ψ����T<�`ۆ۬���K�Q8�nj�牟:7yRfQx����^�ؒWk����;kW�տ���F������R��՞��[�Lͥ9�Y��j,�$� 8,d��lc'u�⯹�E=��E� &GS�;h�3�4Q\=�%��{ I��$��M���[M��i� �Nhx�=����|sX��GkZ�z��]�a8F��[��±���	��� N�U�!�p�N3�O�(�[�86�I�O��ɎeJ�����G>��Q/����`�n�y�m������;�y�_������O�Ȅ��dop��5�`v����`7��W*��3n�BT��Q��e�l�0"HF#K��vti)���lc���������m����V-�r3���dB�R�6-�ͷ=�-0�������5���sgVD6��?��;Oz�Y�[�(�4^E���'�����-V�B�H���Di�8��U�b۲�6�����i	x�CAǣz���xE�l���$p�!�蓊P��`H�\"�I�8z���WM�ɣ�h�M���������2	C�x	Z-l�G
����F�a�@��'���G�4�e�lՁm��SC���r�&����]US���D�`,�⓮h}Y��������¿�A�|�C>e��	�������0�\$W�h���IQv34=�*�/� ��Q��x�uP냿�Na��By��gڈ�x��]��:lDwess�o88���A��4q +�7�{@�?~���;���>EP<�L��ܽ�
o����ӟ�4��+_�:��?�/>�k��kGO��Ę�M؂C����[����������Q����!�.*�E�i�ペ���s�G!Alb�<���(���	�[Qc='�fp{}�f����0胈��/�c��ǎs�n(��0��%�޽{�>{�~�^��������w���/�]�PQ����\�*�+��0d\��<K�"���>1�f����-���kS�)��-���;r�A��/_��̡�LD���|��7�����_z�;��>ܾ}��ի�.C?����c6�K�'AՂ\cK��27�#ө��\��N1�cOW��ݽ{7�'?��^x���q� x�a���v�6�������W~��ӱ�(����L�VV`!�TדZ�i�c�6��فF�'ػ�c���-'q\� b[n����Jd&౵f�`��.]��_>zfaaQQ��S���/�P��p��[���3�Sњ�������&��ܛ`8��\�v��V��򯌙��z2ř���A�m]	�6�ʘ�&e�ݹy�)§�{N�m���BNd~�?ba6��0S]ϋ����q ���&�b\[�F�D�=l��ߖ��;{ݮkgΜ9u�����s�e����I��ϳ�Ҍ&�	�ub�5)D,ޤu�P_eJZVW5.��ɟK�Ti!�=�C�-#�̔��[-�Q1a��P%�v�ΝV�P$0���$�����3夿U�1#�����P ���?U���REfZ�T���HF��5�3Md>�/��F2�@� �'2��22Q`�ɼc�����L3gt_46�}^�,Z�Pc1E�;�,��ah�
�|9���1"�.=]��TGqL5.������.�A�tk��p�OU=]�왚~�0ӕ���$Z��
����+[u�
֧����&A=M����p�U��s���RDq���@Ve���uαA����(�yc0�`�W.]�~���smK�nw������������$��,�������@r�+���@�7�x���끏�7/���{!�`�#��7��*p�ɳ�~�?�?�=�</-?WD
"�\郿O<�H���h�D1��]�c����K��Z�6�H�I#1�I꟞[��O揬����k���a���wv�΀S��a�غ�6[�pFA�K=6�̹Q�� m���p���^���?�c?����?7A�j�k4�=�1
��'��k�������������������_���/~��ŋ�[���u���!��C�}���#��f��س�M?�k����p�GA/���0�eY�݃;�ju�q���5�7n�?��g��+��_������F�ya_|���noaa������'�_��Ͻ���o�~	�l�޴�VK'N�<����I����7��o��Qf!Z��qچ	�+H#��5��ղ5P�J�jM0�BF����X����`�������_|
�6��>Rs8�>3�|���������?��/����mx���9�����L�Ӕ\�g�I����C`ہ��v�9n(���S1�E��p6ַm�z3�E��YA� +>������W�^��MbPͶ[�5,�yc��ۿ�?�����ߊ���>��,��eG^�}��0������Lky�m��@����-���V�?�h�
Ϝ��1�k�-����WE�_��xnq�rk���V�ڶn�>��G�Xh~��f��8�����ֻW��8�w�	�J���9w�'O
���;�O�&�f��$l5��h�z�(.�f�i�6���	&�4���0
��G�~��<�d4�p����gQY%V�<��� H�� �t��P����_������S_�č��E ��>x [��z���>y	�W��rd��P� �����F �o;��&�Ѥ����eظ	Z�p�bF���B�VQ �Q�Ae�[�)���GO��o��O��?7��1�����K��,%I�I6UZ�4�"s8�(�b��&1Ja��bQ���A��q@�\�u	��D��-�2�A.!\Eo8��/҈0�Q�5�I�*�Py�zh%�	�^0�2h�=R�����`�-��F��H h���ZZK���� �b��!��R�wQ�<"�X�"��� �luX9���I2-�9nluQ��Wu��+ѰHsǜ�	��3x���:�vR�#̲�Yd?Ҋ�|R���@h�$��F#jA�� 1d���9;��C��h��-+�.����ǝ��"�'�#���>,\c��K!~ДWiP���p�,�5�@<uww��3�<�/}���7���h�����|յ<������j��+6ؘnz5�H	�$ �#�� ɣ�� /B �m0�]�e[����v������?��dAH��}��O^�fg�{�i���I�hp#��TY�7b~�ᇛ7o޿/�`U5mx$R�.�v���]�vu.X ���O�g�*C�gn.��j�μ���x"�{�'#�LHG3xMِ)�F(2�/�@>^2ɂ?q�0
:�UK|������ֆю�M�u��y�g�y��^<g�|A�4���<sX�OK�Z8>��|���MMM߿�3�8c떍x��y����"<-K���=Κ��x���	��M�����������pqp,�u����~����`���~��Y��[��u�)���G)Xy�U7��L�ȉ�ioh�a���¬�}A��*	����U�+<÷���z�#����^{�٧�v���}b��̳��h�ZU�\�JN���W�:�.�x�K_x���n���NXQ�.x�?\�㻉��3ay�
U�_�&�!6�䙕�y�K���$H֧�J سo_cc��}`��e� ��M��3���
�K��+&���/��k�����s����$�Z�ʄ�?99G��n�z͕u�
����3Xc�V�0�݁�X��n��^�-�TJ�h��-��å&����Z[z�����i
�������H�VG�#�J"�b��T��c����f%��v�[,&�����Z�D���,-�X\`�o$��'�����V����ކ�֭�t�`�j-_��F��Ѡcnx� �P6�g���CL�CU���`�@��F����JHa�V�����oJ$�����F ���]B{{;&(��6�Wd'~nh�7o���g�PU��55Νq�K�� -M��ڡXC�tSՒ�(�a��u�~fE��ۿ����0e>���QEtY�LolSJ(�7Xi7�>���*�R+i�`b��(�Y�p:|��ɀ��ʀu�+'y�U4h���w���Or@0Q�H�;�Z��'�YLF��d�{�z�9$���S	lS����<��w�����}6.5;����L���+R���ih�Ps���9�2<P��rg{&r���"��9���V�9~���$����V�?-��Sykj����a���
�qdp%�#�
<'	G''�i.�p檕+z��O<���|N��-:�صw�������&J�f�;S�t,�E{��@�54�1&�����GGƇF'%���'~�������Z�$��˚��)�UT�._P,v�^����D�B���Hӛ�(KRf4���y�g&c)U)k��@*�Oe���$Y-*��j0����a��kN%�#�hZ��N>���/���N��,�X��hU)��Bl�[*�$Beýh�oq:-{����D�u���W|��G�l�J�
\]٤P�8u]��O�y&k4��:<��P�D�{���H(bux�%�������g�Qz|��2#!P��U2�.�������T|/Q���r!�9���<.wdr�*���75�К��^Z=��Ƒᱮ��FƳ�h0���;��%p��W+�.3f��d校�W�P,��4�,2�L�寚$9WP��H� �ϻ���;��}��WH[�\�D2��4�I��j��
t@MmCuM�{�o�[�p��������s�m�~���S(g�:����d
�d
bbbb�G��Ū3(��x_W^EF�O�
r�d`��t Y��R*�.I���u��r�Ygc"`,�򥝻�� 33T�WR`�VWWc�w���ﯻ��?�裏���/��ln�S�
a=g�1��x��lf�T�.�xF��Y��3�V�C'_j����Qe1������X����DN1kBS.����e=g��b�	��x8�*u&����P/�����s�=���8Eih�'}�����-jz�yu%�̎�P����h*[�4۬��
�T���?�5C����#
�F�~��d��JZ� ۪��$7�Uተ�����-X��p����Y�fͱ�N���#�hn��Yfو����Z�e<DI�?Vd#��⌯������g�\� ��Y����e+k��.0`'CJ�a~J��[-��&錐��b�v<Ka��#���74օ���ޠ߳�]����;xf>;xWC�.������R�E��N]!4��ଁ\%GEe���BY�,��E/d�Y֊e��>����i|r*A�PM\&��d���tH:SI���,eU�t9��B��BY�V�%If�_�Y%�grxi���]n�0����f�,��4Y:W�:��a�A���\0���c��]��8^p[,�6�&f	Q�c&��.���f}�Y�J?��E��Y�ʸ��������/�&���*|��~9��0s%A�Ⱥ��ef)J�#:����6��%�U�n^N�k�9|�@8�A�Ly<	�`2���bƁ��o������A0x}�콁
�P�TZ�|7E�lѹ��w��###`�������?��E����oڴ���;H;7���r���+Cs��Z��l�`�bv���X޶m��\p�M����g��f�O��_ ��E���!�8�AB�� �,�ް���������p�%�,_���-b�OLLA�3�Y܍,G����b��^b^��ҭ��C��:48r�G��[O8�T��E��0�<cE��!{�u�����r(����)K���,-Y�d钅�7o�O��f��*#!ds�MM.G�3�|��P9h�i��<�3~������L>��h��P�A]��!aHNLLB<	�V��Z� �ڣ�^�x��w�͋;��ovU6?�y�	�#"�p�y-V��Zp�?pZ|��~�[�����R12E%~�_��,e<�5�|�����ɍ�Ǉ�;����ⷿ���6�]�)���)p#���w��)��j�	�X(���~E���n�	��������[���!P������'�0�����Ĕ544��G��k�x��y�^�XKc-�d1�������Z�u�e�[�����9��Y�u�%@�`�g�D4:�&g%�b��֬I�|��+�;,�1�A����f�줈ӹ��������/�r9�h�b$�vy�
�\�0aW��4�uZ����	̯,�kkk9my�Q!c{���:�]�ߦ ��*���	�(G,�ؾ;��g��2���̽A�2!
�8�蜬-=er(Z�y�����L���<'Q`L��&��_uU6��xR�"R<-cl���׈�o�}��}��`N[%�Ow8�;_,0���G�����3!z��מ0��"�����Xz13�2� L:��F��&S�oܴw��~���M�Gby�#K�5.��*��TuF��Z.#NW�T�����:nyL�E�V�3����ט�̲%Y@�,	z��J�`�⌡��E����� >p�D�A2!�����w�"'�tRSSӮ]�����U�Bn?��"N'i����y��3ߚ��%�LS���fo����4��.xئ<�z2��7[�k�E�6�,"�p]6K]mq�vj�l�_���A�L<M�8���o��6�22:�hѢ�/�l�ҥ�����f�,Ń׿`�s�R��@_���ll�}���<��gp�����]{�8���ݽ}��LVm|�t��s7�t�M���_٬�d<w"?j�1�^v՜9sR�
��b�QU���9��X.�����[���>�<0�J�%]EEA"�M�(҉U5uPNUXtđ��B?��y��C�qa�n���0�N瞞~w��(F���{©Y�Y(�h�T.W����᱃��TFgw����_��{0�J����lY�M0v���2��7����V�ê����v��n�9�&,�b)�6[S�XWwoss�1'��֦n��?��Y���A�Cc� �ӯ褢&eK��%=>˫�(uz� ?Do0Z:�9����WX�9���d�1�Lc�s�P�o�� �f���z�`������Z��!���L�������%���hL_z�W]��o���o�98��q{<n�Ñ�LFKL#[U����+�&���@�p6M8CL죢�Cԩa��W^yeǼ%l�r��/S�	�������&}6���Nk��t:a�� ��(��_l*�J�m�)v��w\p�5�=	��l�n�ۣ��Q��	<L�XP7k�2�T<dq�%v���p���*Y2Ԯ�]�g��������ʧ������X<'�ʍ��Poh�ʫNϿ%�?��D������݌��P�HY-�~�E�{ҳ�>����X�|>�W,)xS3����
|�Dh�,�9�H`9����-	�o.���b9��狂���f���O?��T������Ң��G$�*��!��`}}}��zdSo��ڴ�Ioo1�9rͼt2f�Dʌ��(����A����KYc�_�\�e6�*|7M����R�`sCؕ$J�*�$s#�!-MLW�<�`4Gcj�/� ��q<���h5��P���&(ɷ�8 5��~�?2������d�2Ū�6�-5A;񬧢��>#(%��攎�sE/�s�@�K
uZR5"�Nr��|�ߡXI_Z}��z�M[��r{�h��.H�@��55]]]�S�uG�;��;��t�T���d�T	J�7���R����2���sfQ�׵382�	^������K��^�Nd}�� �n��v��յ��`pX-沪g����V]��o�ӵt�Ҧ9��ؔɨ��%���\	Z����X�¤����E�h�6w�ۈR�d45+j9� 46��d�j�R��bpk�|	Զ��VP��m���wl�ʴ�7M�~�g�k�poO�׾yKM]�S���x��2����A�D!a��}��:)��0`�r�k��EJ�*��D��e3�P�9�B
%���D)(�&�qIw3�(��t�駝�3�d���r?���"�;#5�G�9���@{ 6a��6e�q����С~�8�(|��/���h�l�28�n���k��{�Qh���:�S.���Z�����Q��n����F㣣j9s�%��q�i��w�~��a��h�N�lǅW�caC\bq���A�8~����[PV3�2�-��Kb4�0��؜�M�6���?6nܸk��+������b�
��6�*kT�Y"��cL�`�N�c;v���߻뮫���G?�џ�}�h����)$?�p:3p�V���944Ե��i���y�7�9;_n(7в���h�.8��(nk�)-�����ٹh�2��)�����햩h\Mu^vppT���~��S�������w�~o#.���W�4O/��� p+&0��<UrUY)��s؞��N:㌙"$�߲H�����K0�q�	����ZZf3��Bm1�.W&MP?������W��ؾ��G~��OEc�,0B��ccc�7��Hk� ��S��@��cc$5�vkuu�h(�?��w�E����G+j�� Ñ�';cf+T�E��n��:$j�v8^7ULNFv�܉u����-o����w���ݻW����Ǧ0TH�����P�.�FI˱���E�dfݗ��F �ã�x��?�k_�Z[�<i�;M����S��h���TU��	,�c9�3������$�\��z�7^|�Y��u����O�Y��:eqB�����iި�g>��f���(�9	��^����n~��?���l&ys�l&�d��J�� @a���y���i�k�rcb�xp����Ə7oưmހ��U�ԭ��_D"�]=�7�v���Δ��СtOU���V��:�@!�qܳ�����U�c���&ضhMOOOUM-aZTz0&xoͤ�l�YeO�x�+%<ލoy��|�φh9�S�(�gg���i�}Q�R$ǙP�%��A�O��A����K,��O�� CL��C�c=s�Ε�^儯�D��ɔ��c#��o|�⺎�NA�߹{���L^.T,Vʸ	������MA� ���_^1�(��T}�32iF�-|j,O����7��F�FxR��U !OeV�?ݍ[-[�ldd$�.]�J(U2�$�<%}�ӛ� 
�rY��ۣ�T������^�l��l�m9�`�}f�	H�Pu�ڂ9��=ؽv&���C�h��w�nY�P�a5�s���l8�o{`� �f��*��5��g�O+��f�x��6w���̞����NB:����3�82<�!�U��_{��� �t��j�y�5��C��pc�"��0�ۛ���|�i��_���3B�Q��x��GC���{K��k����NX��<b�޽��u����W+�l_��6,���P-�����[>��9�'?�gp��SO=��'�op��p��	��\����G[7��yp���3ϼ��[�9��J�Ev�5�$�t�%��˥\&����b��%e߾}￿i```NsK�����ċ/��;�lĘ���+���P��L�f���Vyq�قv�7�Fb�dM{�ÿ�͚��Ǡ�"�*Ngm���u�z�D$n���H��{
�S7}���z���V!��ѐ�}&&�^�������;Z_}�o���Ш��9q�IW_}�	�׻�d�8��D���k0�1M665�ޝ��h1��¼+^������������PcC�h����N�uŲ�*
�?��OKD�Tu��N��{��߼�;w�q��ឡm6G)�f�ext��c�^�nh�<T_Ldc[?���#��T�sι�+dV���V��V���m9E���e����o�=�����]�в� Y{��A���X�n�`o����ˊM��n��
O}�}��#WaO=��$A���勴�b!,��` ��L�FG�,���X�`�QXN��0�uZm���W���!�wvΏǒ�6n�k�|�'�?�駟~���$�#�@���"k��Z$+d����Y��`��Q�����%�^�z�Yg�u�1�W(+	�X
3>2<�u��b:�M�����x�*�knn��x�9W.�����-K�%�����H��Uy]Ͽ���}�'����%��l�`��u��Y����	��i���Q�D��IW2�],�+i��!P݂���ֽ^|�m����lXDbd���|IG�A����i�7{RS��e��#�X{�����,Y�d��#�LH/���XT��W.�6yqJŊ3��T5J�4"��7DcXU"��3BI��g]I�.s:��i�i����v��p���t�6�V��:�����W�£����T�J�����g�J.Y��5ZLj>��3%�IX?v�B�S��Q�`�}&����Dh�Jf�|l��H��Cr�JS٬lr�t�;��Q�F�T�8`��uK���[�j��wh�b����8�uh��kq���T�����=G����btL@����[tv)Y��ۛ�ǩ.�N n�(� ���L�TWf9qZ�U���	]N`�}�J��N�*k,wBb�U��'�T>÷lm]k�V�BC,��U�q��yr�l��P[[]��}2�߽k��7��̑TB��d'�?p�dMV�0�l��8v�,O��\��mvVF/�%��?�E�J@u6I.�<� `,���Hg���i�דL%���J�䩩���2[�B1�{h�#�=��I�>��{o�������uC��y�V>W*�U�A�b�@61�:��Ua|G��J��>>l�;��9pּ�H	�L�Bm�#��xh�����G��T�1��B���8���pt/���ǿW�z����km�>�#�KFm6��/��ܜ�������k�}��y�1,�d[�C�ᑷ�~����z�e��p���g�3:s4�7��0l!����뇛6����/b���Y��l2���?�#l.��F5��ˬUT�HM��{w����]��mmm���*~�����w��7n���^ ��أ�;|;���Ԥ������k�9�Sz衟��Cc!����i����;��1~'��b��m۶�K����X��*�s�<�r��E�igY�M!����n��%K&���y�x{#��Ds�O�=O��QGU�H1:�����	��v;������b�xY��ٳ3�`��k��6�{Ϗ��a{�*��p��t���hU�	y��ݍ���  ��IDAT�p��eG����@M�K px�c����1H؅���[xM��������;�۴�_�ꊕ+�ʯp�\��7�H�ds�ёq��u�UW��O>��S�r����͡8��@��js�'�T�],��2�
f��xA���+�r��b.�-f��ڬ6<�b���D���c�Cd�4�V��^y��7�x*m��՗_v�|Bl��|���a0[<��_�t�����q����v64�_}��g�q�/����E�&=�ש�zzʮ��ԧDӳ�{�ɡ*�~O���L>y�UW�?�tN�L:]�Ă	l����А�M�V��V����{ �]�p�'83��`�>���<xGG�ē$��۽cǅ�^z�%�����裏V��������Kc�pD �X(yM���B	�ܰ��Op�w��]GG'��c�8wpy�v12�v�����m���R%���P�\��:f�(���61녓���b��(�����5v�^p�Lxq���%NWdU~稔�*�k4	�4�5��N�hf���Ht*E���c�xS�
f-�p�4	���2�P�A�kH�l_II���v�e�F>?�����t���?�;���g:c2В��+nN���&�!t�`6ߵm�@�	�a��>�B�8\N�z�l3@���옏+��c���F���(��ǩ�)Y��v�V�4�C>��L�����fL�TfM�2L�Q�X`�EA��M4���{wArV׶�YKbV3B���ί\z���*ċK9\�hQ��^���a�(2�d��VΥ�H�|���ZPk�Kq53�˴G�wQ��ќ�f��?��c��
����*�'Y�ѕ*�:;1��gX Ǯ_�v�ڗ��E�����9��H��x�C�Q��b��R0�`���{�M7�fA��N����,�@���LkK;��r�j����¤��� �b�'	�K���\�c<��_A���f��GA��M����ž>���������ߋw����ƛX`X�7o��������җ�TS[Kin��x]�f���f�ǡ�A����>??��>p[���9�U_?��+��p���e[h<��e��QU��:����L��j^y�y�MU-�����gr<�9w޶�u��ׂ�[?��7�r_|��G�]-�3we�Y�y >���LL���[���y�W�~�y���ڕ��[]]m)���c�.Jb*���_�v�@�>g&�:��SyK_����%��˖�VU�F���/�555�Z����.��q�J�``����s�tGG;�
+D $�X�@�ՒAo4�9Amj� Sn�ڧ�	��{����~����"��,6hFW�K��JeAa�Ѳj��,g64�<���C�����
���|Պ%xǭ[>���O����뇇��������o���+}�۷~�n�Ĝ�k��2<ʪ`��^�����=]�n]C�~xך����y�?67��ki�>�/Pt§�tF��e0[��ѕկ������6e�y%��0
�Hs:m�4�jj߅W�x���������}�P�뚶~��;o�z�9���[mOc#�9����aɥS�H�WU��wh 3;2�.��v�7m�����g����x�
+�����Jm%�I�S�:Y6`�cSS�s���/��`u�&�p2������T۬�B.��OZd� �P�l��otw��
��Ⱦ]�ރ]5gn�t��Ø�RV�^6����nڸ�C��?~����{~�u��c�X��Xө,~��~N���qTR�l�]̲J��p/��tA�uN:����O�3�X����be;��&J95I]�Z_k(<��;���\�bEm�"Y��*�y����m����N:�ᱍE�B���-퐡�b�֌Ky���l-1�De�)Q�yy%����ŭ췙q��PHg�&I�ˆ ���DOfu�!_����p�0[�&�|�$N�����r^	Tϱ�-5^I��f�kXJP��G6�E�q6���x�紅�vw��5�NC9;�z;�jm�'(i�c�&L�j,��KMt��?.�Ƈi2R�K���f��)�>��b��f��3Z�X��,���{�6�I,tѺ����[�J��9�����������n����k����ԷI��X�'�ו���Y�Tf��2Ƨ�RX����1���2ko ŭ��e���`ȧJg��yx"�p�In'L�ġ���d|b���C�r�ֶF��cVS�u���+G"�N�mr*������@m1?�:Dp��%���t:�͐�%g�6�&���
�W�3�~�R`��4�&d��Վ�������.��������h��m�A6C�9������{�eL���|qn�<�Չ�8
AS\pŗ��#��t��=�AV���:��E(���+ 4��ȷ���Og�O'����
&E:��熢����?��:r��������f]]Ü�V�	�T�P,Kخ�1�[�<E�sMY������ӟ!s&'#|���l6��l�:8�@����e��t�P�]�=,�:ǃi�<�H������v�i�N���]�`��<�����Xh����v��0���=�p�E���5�g1x�8</xNn����wm�{ꩧ����,=��
N^.�u���f�iժU��1X�����q���_�x≴4}�T6ñ�~�P����y���O���=�3��%���'�4�Ԝ}�٧�x�`4
l��L�$B����r��kb2G����n_��#V�J�۷|����Z�f��U+A�h�̩��>8���t/�7nٲ���qÆ�q�@y���q���&["SQPw�ܹj��y�L-ںc�o������H4�v�!���^|�ť�C�:�h��3o��A�2�B
EJ	�Yj����5�~��J.�nݺ���n�����Ὴ.O�q��?����>�s�~�QªǭA?���tGB�wu�jll����g����bS4ᢋ.��O~���0����B<�Hgr<�c�	�Q��E�õ~������g0�x |�l�����o�8����v;<�F��<����1������c�Plk׭{��_�{{C�<.��-�4 ����4xE�B��G�[�c����(�?��@��P9��`��C�VV����_����.�3�� (��+�x<�Ͽ��f�u��`�$����7���x������۴i�}?�.��e��('c�b�6�6�58��
/I6qWch]���k��&_L"��R�H��dk�!qtΒ��9������t���=;��@��!9�0&���!D�X����"U?e�t�V���V)Ȯ��J���bi�/;����T{���,�fD+�GE�F$��`�����������ڪ���%\���������Y(bG�Bp`<^\������E�fr2���<U��+��TI�M�?�3U)����;P�Hd4���@�x��A��	X젒X�D}+�����*�O�d;��,�������r�)#\ļ�������89>��Nau��<W3�VY�Dɱ���q��Ý6a��z=)�T*MI?�tX۶����>�;�!��X�\�UL`$��(^�b��� ���,��~�HEC9�o!��8].��̳rVˬT�Ϫ��s�g&��	�K�rY��&�&��퍧󬞥���&T+��.kT;<:
7==n��ի�v�'�Z/Yr��������ϳ���770������`�S���g���x8i���<'�c��-}�g�v��Ö���g ez{� U�S�^�G����(��<2�fJ�)�W��u�=x��`(?ɯ$�(v�����Z��/��a��&_���o(x(��#�k�XAqY�-[���{�
���8������6o{>���́�OU��ܹ�]x�b��YI��YQ��D������L� 8|��M����Ƣ��v�FQ��a���w�׵����<~s��UMao	���K/?���n�����26x�&�S���B}SN�N%�W�~������W\q��ڨ��L���i?�`0�UX�&E(��}���_V�X^*	���+.��~բ�R.�ɇ��lLf�B��zäsԇ�j1ޑQ*Vٵ�g���~�'<KSus�C����QŨ���f���mnx|�w��lo��+ן|�w�y��O�wk�o���k/���
�%��^��_�U�SϏ@nh<��u��)������0�~�����A|��l��v~
�5>2h3�&�462K1EM
�w�I6�u��]A����l6S��A�L��C�+=������s�#���+�]�J�Fs,�<�s����-Z0�C�l�g��BI'�}^��H��`Gc��3Xe~�o/=��ǰf6�{
�h��&�w��a'�Y�T-^z�O��x�-��6S�����s{nkK8���L:QTT��	f�Q���/]=�s���o�3N�X�����X&�����G,��!��<Th:�aj�\6!���b������&�/�bv����7�RښkamBA�|6i�)n�\*�~v��z�+WM�P���U��E�a�Ѵ�d=�3GFG���\�������?�Ǜ�@���ZQ&��`���/��FBI��s�l8�b��b��Jv�X��:���)�:na:Oم3k���Mz]�jL�/XP*%�����<x�A���X�U6<<��Q/J4���R���D�>�U���@�����uy"��D5^*������J��L`�UpM<n��łY��N�(������D2�Kgӣ��5G���I�ⓣ����v�,��}6e��.6��T����OQ��H%��7��_�b���n�f������SB'͔mC�1��<��8�w ���!���syڬg*���q@m~�f�BN��>�d��A.7���-�l�z��#�c�T�������d�XΩ���6�@D��7<2�o��z<���_1Wd[69��V��HӵJ�X���N���
E1��y����^����p�90J�*��e�����J[Kg2��:�fP���|����k�u6�ud0j��NG��%�q��B!91�/�?v��d��ML&p� .�gy���ݠ3��C��I�*�f;q��F�;4�AC�f���������V���X�J�ץ�Y3�8e$8���K�-���Hf�U�b��q��se�gbt�7��hj8���O=��?���c?�ez�W���T�R��F򶩣���V�6s�n��4��+<a��u�Y�{.�Gptllt4�D�zCss��E ��Ȼ\^B}e��� e���d�Vjp�|���P"��%0#�9��b��_��〙7#hkkc X	����d�D�o���@4f���>�護�·���J_U��_�((��ް�ש�[-P���^�̐nC�}���jx�0�1Hy�{���q����e�r���{��!O����c{ޥ\��?|�GN9��K�-Z��?B�n��/��l=84�)��>��/���
}xoP�	�u
�~���!���)�L�*�wth�K_�ڛo��=�|eB�(�	�![bhᬧ5eI�#�c��9��{���M����j?�[3�~,w�X��l\�ŭ�����K.���hk����,�8�*7����?Ȓ*�&�i횵�Lbǎ7\w9<'��SwpXʐ��p��#S�W.��LF�ި���_y��������qӷyϨi��������y��0�z�Q��?���!������+��޶8k�Y�B�̶c��*�O�1��Ύ9�����w�3�=�9�H��j�*p�11��Zmذ�/��,l>~��s}R�B�;�F��4�Ǧ�q���;o�֭�|��{F�G0_G�=~�c9f�@��)U����,ݧ��H.�
�� ��~����!<6j9QJ[ʞ���#�hS(C�*P�u�ɶ�`�֎��Zw8lpaY�����ǫ��.���p�7�qԚ�?�p$:H91#���8������͹袋���!4Bo�㴘����>��`�clc��P,420 Q�4������s8���1���e����1��L	�Ҽi�b�F��D<BXo�P[K]�g�
�6�AY�r���(e����c|r����21������K
cc�y��5ԭ�$��	�6��S�����g���C!���U]��1�S��7P��B��(e�շ�P��CԸ�e�q��J�]�_�|�Y#�^w�ON�N5z*5r��,Vw���M���������5�OY=�\�~s�ɀ����:;;׭;fpp �L�Y�fl|�3�nU�MŰ#���V���j*D�\��Wm�g���c��|s���NoU2�n[-h+��P���C�*��Qe����1�%�[����<�����]�@��s�d���N
��H�2�H��	��S���@u��<�0
�?_��O��ɕ��3e�-���!ĭD��Ҧ��J��g�1h��T��:��g��pem]�_��Ա�큭��ځ���0	f���~�tA�y�\r�Y'?�����F]]]CC�5�Lne9+�����V�3.��o~S���޾���ګ�=���zL��q!���\�:�;���r�u���;����� ����ҿ��h}��IaMm�f8�9�n�yN;�i���FǇFƆ�t�5�34>Y���
�<��u����s���_��,��r��f��w�yEe ���ٯ�FY2J��ыT�i�RQLLa�ᑁ�m����
8�zQ�%<j.��F0P!��˅�N�m�x!4{ݥd�whH�ĩh"O��É�����\��-���;�\y���!<>cX�m&
j��vY1��9+E���Q>��+nh(k*�zl���YC�o���WV����cc�v��?�:�M��������C�"�<A � ��޸m�c��v�%��xJ�曾������~���+�C'�0��R����&]��=/���S��8��HW�ʥl�ՅS��j��l�8GG�b1r���Vo�����7���w��x��9�,ۺu;�=8�MVQO`�����X��d![V��E͠
x�:���������Ԇ���Ϫ.�
&1].�����X����^{�˯��kCn��6~�6�h$B}P<�r�TR�Ԓ'��W�jM�}�k�cV�~�&��S�1Y�dA0��:�l����ZN&���l�Iu;�;>y�C�᠟~���n�	5:KҤ�3����Q&�2k�,�U˾��Zȯ8�¦�5��ށ���F���U0�e35y�w��������t� ��bbbl"tz�dN��eK��p襧��XĀ;��`M�Ř�l()���$�&l�n�~��E���O[���_�+�V����&.�W�����7�m/��^kS�O�u��-���/��qd�D���w�ym�$)��Q��Bcԍ�D��j�%Q�G#ccC���O^�+wm{2���6<9�dUC}#�#C9�����{�����x82<���5KV-s�3:ȵ�ӭ��rS,�H��Q�*�zhn����ۍ�6�&���%8	I�YMyȮVP#4F�v(oզ�}{R�XKK�S�A1Y̑~�z�i��7Fu�N��0�MH���������3K������}���5���`��Vw��M�G�9��_�x�޽��m�
#;��9���(4Z�����7�L2D[�l�k���/)�����!��D�PU�A;��n�.�5멲����H9n��S�� ����Y-Ѷ����|s�j2��CmO,�5��� �%w�j�mm����n�;=�+��4��l�����Z���(��J��r9��w\+����L&r�� ���T���JĨ:�)M���9j����
[�Vo`tP/ʅ5�CݽC;`?��/���'�$���te�h�8��иP���ƒ�fk3e̙�tR�'�ne�zWʔ�7[	��5�/�T�d,�ZͶ�"�2)���ivf���{��9e�J�)���{<u�|�N�j���c�CЌ���vn��7���w�{�u7����'3���ރd!��)�$�RmS'���>���E�����?�'�x�-;0f�����RN�!Mu�^'ф	�A�eKB�ßʐc=<2;��/]7X'a߃�AI������55u�!��e���^�yM��&{g�/�N�'�\�E���2w�y�G����ӥb��Oƫ�N��7�d�z�
�*�?h}az? �G��˅I����M�x�:,T^�lcŔXϸldd����3��g�y��o<�3N=�lY/���܃ٓeE�Rd���V�t�rQ�p924����w��x"u� h�"�G��W�`���z�{Zx����x�6���<o���}�`\/��x饗~��'���3�?o�V��� �����B��egT>f7��h,Zt������<���?����
�m�EF�'!t����29d<)�O>��3���9��������v��_��l$}���͘J%�W�g2�ry�(�t��&L�������ݠ��!ut�ۇ��Mloo������o=���kO:�rI`����@Iڊ�r:Xn�#��(H�Qy��1x �����UW]�ȣ������:j�����5�u���	���pMM�ꫯ�a%�����i�ᮌ�n��%˒���?��[o-��*[X�v��\B�(&��� d����p¡�
߹s�)'����cv~��2�$�D���T>51�+��<�?v�`0?�S)�GԊ'h�Rc[��xa�a!@�,[�J��7��TWW��!G��K�����4��5�����E����eP�`E-X��o0�!��p��˴�5�L�ko�"L�7��*��<�c.].P]B}(�	M��Q�jwSTF�Jq��9眃+�C{����w�|���vdS,�M��E)x QfV�H�.��Д������5vtj��*�4EP�Y����"I*b.R�Cm��:FY�=,wz�b�����5�ވy�F�#��C�{X�-�-����ю1���ީ�(��v�4z���c��:�ʯ�L��Ǖ`90�?h0:�s��s���fQ�����:w�ٺu�ۡA��8/뒔�LZ\^V�tn��y!p�S��C�#A�;���Z�<eQ$�i�����&q@`�ԉ���c��D1=E�d����U}�Hg���n�\���Z�����[���j\-�[��m�ѫי�4��ŋNP�B*��'��_,"j^��r8;�)���~JL)���:���RZ`���x��14��u}�)f-�0/��pp�@�ZG��4\�{������r��IHqώT��hj�!J�nֱD�h�~����7�7:�&$]��H�3J��B���olt�����0��\`p��ӟ���7?�����{z��n��p�
cR������@�������X��,��{���_y����c⨨T��
隲 ���I�r9)>�7�k��=�XH6pB<��!ĀF0N��0�oD9x7���IE����Tg�Һ����}(��сG�F��x�䘡�����?���[B��>V\���!i�A��,Y� �,�ן��_��+_�ʥl���֬���t˟{�����R!X�8��+���H�޽�����UUQI)�zC� ��j�h�h*t�\�$	�t,�X���%1��R�d�8�A��T�-��GFz{�Rx�W\��O��曏Zw#Aex�j�g��j1���E �'��k�l� ��/����ӿ������wS��U��X"I!}��?ֆ�a7��͸�f�4���Gm�N�"WB��u~��O<���?��%�iU�]V'��(�J��[*����!�b^�VS6��ZLSS��B~ұ'�I&v�=�裐<+V,f<����������|_��ᑱ�=��Gp��B �0�$�͜/��LD���0��N<q��n�eÆ��,�T����d@{�����H���yg�>LX<L�z�T.CEZKt�d��g~��;��rg[��B�"�,��u+�
��I$���l�Y�ͤ�Z�P����6m~{���ν���@�i7�'2�,���X�ySL1��D����,)U���c�J!�0Nޫ��-��l4�8�D\��'����?yLe,jZ�	S}��;�ޚ��R�ˊJ���M���ڀ�e�<���u�̈́KC+%�-䲞5 �u����B.�����3�r�����hjj�\D�i���y�������d��q����r9|t�S��@U �?����z⿳�RG��o��5:<�~�zW`���6j4%��Mj*aM)B��b�{��.τw�Oצj[Z/-��x��'&$�-V�~�eC�h�9��D�UT���ґG)�)�:�Օ��Ӌo-^�*�N@��ܖ@����V,3Bx,�i�޽�����|�p*���2ճ�5#S�n�;HZ�������S?g��ikqZ���,�F�>W�%3Xs��ASL�[���9�t�|2Y�۽U5ml��%�����lK�`�������ꫫ3�V{jj|��h<>��h��H�$vՕ8�{����y%,c�ylt��@WmukuC�9i�+dڝ�Q�Q
O���ꝃ{����k�����(j��o^���r4�0���ʏF�CRiX�~�i�)����qM��śv̭2�ʩd��h�&hf�%�(�g
���F)�����#�K*{'�&�����ò?Ip���d9Q�;]�R���	����g�dA��bͥ�^D�<l`B�Y�f�J�a�����fы�X26>˦OR�
�4�U�D_B1���z�u��Sx|��u��U������6�d�J<ext���vܱo}��_m�K�]�w̡������!f�Xz{{1}-���ˎ?�ħ�z���_oo�:\����w8ݔ�2.�sS��s��W^x�����<�� x����c��vh�*G��	���1��}	��f2D⚔j���>|���D[+�*6��˗/��o߾�l>�#�夲,�\���������Xx<��[+�,x� A[3�;�u5��ߪU���ݻ	3a޼y��G|��7�������u�3O��HA+�Ã�f�D-ީ�*�޳/�`L��� �ru�eKqk�@�V^�M"�J���U�o��@��y�ڝa���eb��`Y��o��cǎ��>�nho��5�Y�|R$�Ã���+/�}�݇�w��=�䣙Ӗ��OGȧ��ۇ�<�1��`���\�}({�-�R��]�x1���~饗��g�}��6���꣱(��Ș-v����8�W�x���:܊Z!c�V�ń���0Q�����k�X̼0wK�R����%p*�t��'TEww76,�S��)��j"�[2;�	�njC��G?��_q啗^z)V'�B�VcN�����Ad��ppALnh�{|��Pz���ߟ{�L�2H6�f) 26���$���2q ��rӺ�n���{����H�t������v�:��׍����1L���B���/%�d�8#Jf�w**N���ur�as��
�pϞmO=�T*���������s	9n��Wca�/�z�
Z�r�c{�)�>�,l��+�4�����O>G��c�(U�������z1B�	��1_:rk���$W{�>��۷ooin�?�3�J���W/���t:g5�t��B���lpwV��>7�[o��͆���Kd��A�@$�����zz�VVN]�sI�بC.�v�B2	�z0p477{k|C�'��$�4�-7n��Lx;�!��	F�Ʀ6a]����$�κkN1�E��F,k���J��89J�6�Y�&S��'�
e�[��أ��;�z6�%Am�ŉo�#᥵��`n����+=U�x/�x&K;QGW��s3���Ph�r�<\6��B#]XGn�HJZ?-L�p��o�r2����N��`W�5�`'���O�W>l�H$	6+(P"wuu�e�y\��L�$I��2K�y�msKSl*|��sI��p��FG�`7�t0<��`�!QG�@�"�]:�r�b�[�8�/L�TY̥`�;-�M��~ZZ%
������$�C"��<��֭[�)�Z`�I#�Y5)!kQhG��uFX�����D"�e�2�h*!d�����,������=���o�mQA��P��_��� Hy�t�`��|�����	���[�-�T�F���y'p�������n���o}��?��%��d��z��9��׾~�)���7��$�E܍�{�iЖ��T���xN�p�J4a�Yj^�[� D�뗻�3����j8�� ��5�[e�ǿg 7�}|����H(͇�ܒ�tb�ann3%�a��47�-6�|��0������c��ֆW��r]}}(�<���׿y<	�9b�QG��R����6˗�RL�-.�YO@}r���x�-s�$Q���b1�ͧ�6��d�/��2<~�fTC�D���Րh�	B�̹T�7�-����^��X?�?�����REjtΆ󆆆^y�/;vm��K_����+��t,wC��7y�r��)ԋ�ms����{^{�U��.ZD��,��x\���l��(��D�� �#�G#��b����,�LT+UU��<���a �p�߹}W,օ�~����A�U��������`�d4ӄ˨&�=��xC}m*��F��G����|����m�-�I����z	��������"������F蘸!Uĺ<�U�Xf��j%W0�)6ew�A*C�c G`2���{뭷���;�_��'��MQx���Fʋ��b6�4�%���<p���nɢ�޽����'��مu����Zߦ#�q�լ�g�2�lv��DS!�A.2#�^H
��F�bJk�,-Y�p����Ēsvn}��ͫW�>�������42eE�T�o`�@Zi�qhd�d���R)B5��OX���Il��C0䓱G�ю�a���ԩń����Hq�|v����ȝ'�R��wY-W�t�J�%��b��*��+����C���k�:փ�&�3��J͠s�A�ܞ ��`���'"Uc�T8试�SS��v��g���P�`�]չ��u*���3ӓ��	��BD�a�I�\l���}?.���l����0`�W .`����H(�hB�t�Օ������9]3#���z櫮>a���^y���7}�߾�yX9�|j��QK�X��V*{1_��y���&���6.&&Y*إ�o�5u��ޑ_~�~�7�u�_��.-.��,���4KA��l9_�.�g�X�G���/Q�!����}���j�¨é���M��rerr��[���$;s��aC���L�|7�v(�e������ �>C��*a*	f�,�-�?��;~�_W\���?���L���������8޺���͹L��8V*�-[_LNc�����V!��P�}VX�*B��$/,��v��é]�vV�kˋǞ��0o{C�����t�n)�(+�mg�B
V:ݕͦaR�a��--~�s}ы^�u˅���م��A{�Ƌ��&��&V��*���z��<T�l:��e	���PÞs��.4�d9�GʉkQV/x;����!�����;'g�2"��5��6Y;ᔱ����4u�;
��P�Y�ZidC���|4v`�U��᫮:x�رf��5�9�Ђx�d�V���4��9q�ēO΂�����������)�Ӵ����]�Rf����w����F�7R�ޱ�w��s�f��R��������;}O��68=_SҁѤ�sb�?�������w��Ͼ�٣ccǞ<v���N�[*B�������'&NONOAF�޽k玝���[���oC�~���r�z��쮽���3�Z�C(>�IY�mm��
�(8�=���⃘Y�K�wSLh|��!�1	B	�k �n��!�O�S�~�} ��3��܄l*�M�/����i}`(5��W��߿_v�!�B�M�3�D݄�epLLeTr|�G?�Q�V�������>���8��(/T�>�ɏR�^��7�Ч��a[��H�[�.@PQ������c�����-��m�)v\�+�筻7`MY���^��!�ze��o|c����g>K��[n��?�����뽕����Ao���k�B ���o�ݻC�ɰ�Ny}��p�-#>ih�����-D:�ԘbJ1��hj��E�_	���p(��$���7}���׷�m����-��U��CӠ��	�y�� ,�N�}͵�./��x�߼��X���9aܯ)a=Pɧg&A=x(��@�O���t���T)N��͗N�;J�
�p`h@����i�&��t�m����o~��u��}
۵���s��[�������C�����KK��x�����C]}�՘R�	��'ȰhQ�=��c@�2�K俁(�kRm4�̙�-q+Ƅ����MIɬ�� �'�8I���=c7-̓f��b�'ɳ*������
���,D��/۴)t����?}�߄�^x�N�5���9�PQ�y���t��yT��v�:N=Q�>P�ӹ��$T|��sl>P�w���� �l!*�h��!�<��A��BGGa��������B�x�����/>k��]s�5��R����Ν;-�"��'��[�
j&E�/�=4����*�U�*�8O6S(s�O�_��7o���������X�VG�Ϝ���J)H������@6�E�n������(lٕ�5F�k�!�f��w�����gC%�8����Jy�X4<��"�)��]yj�TR�9,{.P�U�WBH��mw���;�޸o׾�6/�,4[�D�Ȫ��~��l��:0��W@9�s�䏵�܏N�
��hu` �Ig�����=rVi�4n�D����z=�jE���|�zE��]0�,Q�Gz�����m���7��T����Ļ�3��PI�D!K�X���F1D+����d�|���s��L�3$�͕zr����>��B�b"�cf��#��D�B�<�!up{!��Q�B�ΰT��w��w���U�!K_�;��ze��J����w߽o�6\�aH��ɓ'��4k�*39�9XH=�g�\�,�<���ӟNM� <�'���|�ș ��
�)�!GH��2�c��1K`D���_����ڹk��ݏ=���iq68�4_(�\�����R���nx�����}��������G��1�T+��I7\�´��?�b�a1���V ����DPb��ִt9S�{I��w2���#,TB��=�\E���F�U8'� 9"�)��E�Q������;wS3�V�vhhC��E#�`O>����/�ա�=�	��n���C�,*�`snq�+7}��e�B�:P��������)���)�3T
�wI�6Z��v�J�r���7�b���5�@��Q�Lt�Tb=Μ����#*�qZ�����-L�T�:������l��A���#����w����b&�Q�E��0_��W��gw`��p��IN�-mߺiqa&�6�^�v�xfk	Ɩ��錭鄃Y�S:r^�N����J�Lm��J!�R��D�H܂#�{�=�O/}��wݵ�al��t��O��ӟ��/�˗]vY�2 �\)e��
B�L-,Φl�2������'��\.]u�qN�E��ä�S,@G�d3e���뛭nK�R�3�,#��փ�L��`o�;Y�Me�9�@���JQ���@3������?���}�k���Y�F�'�>�`����i��>�O�����~��?�/�����Oޚ�
�o�^kf)��<Z�Q1��m��ė''��#�0Ǌ�cфvڶ�%,q^���Ӷ1L5gx��RǮ�+���7}~��CW^y���j9�섫+K]�=~6���*?|e��68T����V���n}ύ7B0�ݵ}ۦ����GF+�9U����Y\^���Z��7�<���J��5s�Z;T���<�UN�P�ё�v�EMXZ^�����8z���M;/ѩ&���jݎ?P-���[sK�v.[��rl�r��_�:y���^�qCe���/����R�h�ΞX]�65&Q��A]Z*�i��J���9(��8�G�0bR���sz��G�m���F�}H�p�gNO���;���J�y�K��A��4����9�Vn�94�3R��bud��<p�*$˕���T>G�_�L��'���w���R����^�*;B�H)�H�=�Y��-N�됥+���9Ds)#\�^SEG��7��{_��7������߻���l��g&������3��z��6��jf��*S�+�B��[u����X̋_D�����������d��Z�GNM��r	K��A��)�MWEW��Nr8������G���W;v|��?��[���˯zMg&NM��ޱc�R�.>��mXE��vR�r��3IѴSz�2�8.��`�-t����9�i�������6�l�J���}ם��5���d�_�~��(�Sb�p�L�َG`��ե�.Xǡρ����k�`�ƱFmmnv�B�-eæ�"w���N�q��bgd ��+�|��^]S0�x�0��{���f����C�M5���s���������n�A�n4��J�.��
�����u��0�����-7�[�z��^�?���`�@Cz���!�`-p��:Lp���J}z����ԋ���ߒɑ���/�;ʔ:7�48��\�b�+�m�v{�Q0s<��0�1B�|+�t|� ����v�L��W5��iq�$��`҉t&ol��O�E��!���kW�)l�'�7��Bړ��FL+��g=�Y{���fN�5\��:�9T9��f�%*�'na��k���������=％�(�����jܳ�j��X�H�Jb�dF8ו^�ҶH�!���q�l�����Sw^�/Ps3�LRˣl**�J�=�(=jE�(���/�7i'(�G��A�E���Â�d.�O���FkF�V Ё'��=dbv��>g�㋃���J��1axE������H(C�3��n�8v����/��;~N�pO�
�S�Pߗ�ǿ���m�<.9� b�L ��er%ab��'q
��	X�����,����ɷo�;v�Y��|��B�o��ub�(�qd$t�ԩ���}�:����YBf`�~@���`u�����g��Ӹj��q����J��(Y��3IF��v]�E{ ?����`�����QsU�.j]��E�� AH ZX�����޶kW��W������[�����Q	sm߾m<��_}����.9HƔ���_~9�ͱd?0ű��30>�2x�E�II����J6"E�3��G!XhV�tIW9hG��������}o�����
5�u�#�&P� ,������5���V�����[����T��n���=[U�+.r�igY60?�4����*���9�����n|��$7@5x���;1�7���7�Λ�����m�+/.�I�S�x��%�rI�0;�|����(�}�{���/�3����lU-��/����!0n��K�4N��@�E��D��:K�t
�z����Q�El�G}���~���?����6�oV��ŵ��Y�m���;2�3��5rm�u|涢+xG���k	�����?����'/���\6��]I�޲e��+Xw�������T��{u�Ac��B�m�����w���}�s?����ȇZo԰��&!�)T{�8MX�)�k4��ܼ��=�N����6�[�/~���r�����.�j]J7�Hl�Lܺԗ�UmeA�ӽ}�m}���!�iu4��v�m������_��k*#�ٹ�v�I�/|rv��S���Hf��HZwO�k�́� ySf�n�h����������0��L�QX&��T��Y_�oS[��kA��0�2i�`^�^v�p饗�ך7�|������o���� ��4����1i\$E����p-�����v�$-�6��`����q��d�H�&����)F�����5.�c	|���HgE|�A3�5���S<B�N˼���'�V�9����ZD�~�AVl#�`rr2q,����;���\l`�]�/��"�^j�ݵk&��ç�x���-@Ϫ�+�-��53����@��J[;v�P�n�3��j9��4��v4R�B��n��?�vi1��v�ٴ3l˞��䍍㕕���o'�R����	R�}Ϯ�^����������G	��v\��ϴ� =�"�3�����NM��`BA��u��:��<�����yES�b� &S)�|��s���)�=���v.���@�sK���1�L�n��g���l�F�T�F<�`��6Wc��08�YZ���2]�}�`ii���o~R�H8zs�{�`4f���������5�UBFv�i��3��r���(���<�;q�T���(����%�����8!��Wϧ��.S�i"����=�c�`|�\�����������]۷y�����w����$�HB�3{v���[o��M�OQR��+�t
�{�j)�s{�а0l�}Pј�aǇ�P����<�)����O��n�)j���X{�TҐ2_�9���qr�ʙ�B�������+�x�+�[e����qf�X5��r}jeu���v8�����'�����_s�.1������R�V��`����ǐn�x_����זk��v ��2�HIa��QSg��M�c*(AW������j�V+�S�˿���ŗ_��g��F���u�T�2�/Wr�V������j~�s��\/d,�I��b_�ګ)��v\пej��ji�J��֊�R�"]�.Q�H!_����%�j���y+��S�r��֨��@�N���þbk5}p��}��ƿ�>����ox��G�Y��[��]����������Ss�S�|�+Ǫ���|�S��xu�ٶmtx!�,-�R������9��v��(9à٪cL��JH3�T�0�?�+V��t���(00[�N����R����y�W����1��ձ�AӾl�/�˩y�X��o&J3��pyl|�w�}�c�^��+@5��?
�����B9V[G榧R#�0w�̔�;�_�h����D��$�M���\��j����EWk����K���?���������w��R��}��ٙ��}-����MC����mC��ת��Ӫ7V���F�F`�㞷��y�fmǎmF
��9>��˨j��	�3ѵ�r9�F�V���.VT�<�%l�J��������?�ݧ>�O����Ƒэ#{���f�MK7����\�P��<�7Z�0_��VP[^*��B
;
�桭�7_�������zۻn|YS�V*������NF�aB	P���(��}�����*T4
�7��b�*��JY�2�C���l�����o@W����=��/%���6Ugs�F�4��#+1�+����� �ͷ�]́��Z���I��`�a�8̌tl���HOl)Nfc�GQQ�",�0ҋ/��Ki:7m�$���������H���' B�~��9�D��?��\��ً-��邒</��+�o�)��"�[����h(�k���Z�R��1��Z)6.�'u�+p��$�\R�t����Vkp&|�,�"U����^kv�Д�#Ϥ�����3�=�4��#FL�W�Q\��i3h�F�Nc����ߑ!˟3|P�"��4�J� �"�JY<'$��яc���E��	�5W�V�K@�[wˊ&}�lY&-E)�:�l�AVr����o���Q"�%_�g#YE��G-����Nb"��
,��Oyc��əx?E�ۃ4#^5V6iQ��:z��j�f�rͫd]����%%.$ÇGy�s�R/�s������@�"E$��ꭱ|E>�!�h�}����t�%����$_��������g�`pd�50G���_s�5_����W^y�����f�V��\��Bsn���Y"�%���\�֖�V@��>u�`�(Ô޾O��!D�Re�<|g�eg��I��u��ё�l�T ��$�穖���4�����4N���vN��k@�K�L��l�َ�B��C.Cթ�\V�(�#A�[�/Kv�Xi�[��.�������o�ƫ_�����0������@�ٳ���/�}������g&NAڸ��2c��"��rUQ�G�=�U��ǩ���+W��C����%ȍ�\�)*�8?�x0Qq����o�{0��-���卿�;�zի��2�=�C���:��;=��---�{�{wo����n�������B�޶yL��+��f

�x������r�<����*7d�^5#�B���*K!����wOMZ�JR�_��/�c{���`&��� ���H�~X����);j#�co�2.|�]?��?��G	s3�y��G˩k�"�E��\��������^�BK��z���	X/�^ɘ:�Y���atj�e�}�#y����Ts�
&Gר��L��q��3��ݻw���ÇA	۶�En��}��{ϻ�}�]w]~٥�u����OZׄ�7����	�p'�k�4�/��Rہ)/�~U1FGG��k^󚗿��|�;�?;;���J��,Ɔ�#nl%N�V/��?�@C�秧�:�2�x� r��Lm�BI���.���ʤP�aJ�4�Z+�?1󧄃8��ID��Kj��/�����?�a(�t���g�Mrx�.u�F�Qgp��mX����Zi[7����#�H��*�,�. ͞��v���Y�-m��j#���Ky����\&o����a`´53�y��g��:$W<��z]b֡ƥ}]wm��v��4�h��ݵޥ����lSzP<t�ԉ5��+/1�s��!��6��2d�t�p����YU75�8�m�X�xl���L��\�S�7Z��~lp$�xt�+� gs�������$��*mᵥ-��k�iz5,���2-2��c�$\��NTk�a�t��'5`��ԁJ.J~���R"w
-�д�N@U�^TQ�i�F��,Ӣ>$��dm��ӧ-�E4����!��=�]�j9�pia���::�)d3F*��{Q:�ʰ�䠁�N4O�`�SC���|�icW�y�4L�o��y1:�p����P��L���U7�`˖����3?758R�V_X�(aG��vcl�8\ͥB�jsM��:����v@z$�w���F৅[�J�"wmiE�+˫�5��A�.-Y&kg2!�S���������R�Y�foy������ߤ�t�zH�>>=\��߿�>�A������:)��N��r[k�e�\�N���R�Ð�d�*2i���SR�H�T)=���ݖ�ۆ�I�F�ɬ�52��1M��5P��k�����d?��v;v��_�Ҧ�՗^C6�0�Ecæ�J�0"�l޸s���?���~�?{�T�h��F����E���م�4�"��z���s-�B���B�:���M�RL�VHQ65�T3�/k-��j���dPb�L���ڴeߓO~���~�7?��Om۴i�ޙ�9mZi�	*���	S�����8���ǿ�Ϸ��v�"r�-,�� ��ڴ�7�l>����Y����&R_겤c�`~�g�cCH�V�W�p�����������߃L=�w�ę���iLS�6֚����ZMϜ�u�>�Ԩ�A���{�@���=��n�9l���!�k!�jJ��.��C������<�H�K�8��F@4Nr�����>t�-_�2���\���;7�85[,�k����O\p�E�	���q���upփ��W]
�����w���?���Ϻ��y��d�%�K5U��Y��'����]��^֗T�Ra��C����R��n����X.p��
ff��+��z+4�׿���|�+FG����s�]�ˋ�vP�*�]���<"�}rp�z��Qˍ�A�سk�d�sL�2��%uS۴	�XLY��
,��;��\Q�I�$2/%�O˱n�I"�|H������O<!�D����� d�򙢪��<��I�?�&����!�lT�����s��R�2�=�*&���]���?���S���@ j`#J4K|2����N��!*��'[Ĥ���w8�Kq���
>��# �T��[��-#��Jj=�N���J∢���Cr������-�a:s6Og2�L��ݙ(�*giJ��ŭ���tBH����H���-4�uK&S��]��:� ���/�C�"�7�r7��i�{ɳ���
lCm�z�@�!gK>���=�M�;+�����uϯ*�l���j�.a|�j�SF�����J\S!�ŋC�^Z���R��ks9S�K�e/�^I�@M3P�{"�2��+/�НEŖr�R�ݠP[�Q�=K1�,U��*�;E�i5��a��fZ�~q�&���8P��S�,�5��g�)���׆\)�Q� GU	;,��ԓ^(�+.=����k��ၢ�<����U%Rg���W���e�H�0=m-��a���D�Xx����6��-m���b"�Pu6c��ǟ���p��_�cǎ�Ӕ�y����>�9����?�a����9�;���%�$ol"!-$�æ^ +��'Q,�<yrnf���˘�T*�j��{�v���lUZ눢8v��a�u�P&�n�Zo�~������G?��R��'N������~γ�W�_�[�q���,"��&)2��ݦ�'��o�4IV���~�4�[���O>[B�nM��L(1�����~���s��7���4��b<���ۑ����k�Z�����;��G]t�o��oB���_���fe7�����O�g(���[����$4�c��Y�\����(�IQS�N����~��߶u��ܬP5����0�<�t�+�s��9�ȇ���/�۽�o|��eW0+�<���Ƀ�'�
ÈW$F�x��aff�T��P
�s'{�5BT�K.�dbb�������?��? �<x�������R�23�����J>�Hj3�����$ɭ�b䋋�"\B3�%�*$'�+�	C��E��r�s��~�i�/�^��q����,�-�Cbt6[��p�("�/�&�/tʶ�\��JY5B=SCVj����Od�`�ơ`����B�ܡ�uC����V�/���gn~ѴlV7l_1T��Sv��`h���]�l��!R�� [�(�E텪����a�]�w�g��`�e`Rؚnrc� j��������r��TL�=6l����vI�t�6'd*����yQ���V�� � u��xp�!�!�?b�7ƅX��w�/��>�6/���0��]1�q�:�9�E1N]����Y
c�*X��fa&���T�[�(��%2C�0m�P��_Jܰ�Bg��)�iħ�>������*����Ɲۭ{��S�e9��3sr[�շT�̌K�uR��Ie0ZS��@�i���Cč0Ҍ�a՛����wh��˓����� hM�B�d����1U�KU�Xs���v�rv���ѱ�\���_[���|�k�(_ ����\�t��z��;y�~?���Ԕ��~P���W��d	)3�NU+�-elhn���s�?�"��� *��(�QT�E�ƖI�K��t�┞r�`�2B]����쁌n4r#9�����H̣R,ᾭF+�]+��3�a����l�v��+��H�ρia�����i��Iɧ��}]�%�Uxzf�2K����-��6=zڱ��7nھe���g�m�X��˥3x�\����]
uu:�1��q}l�c�_^m�5��Mo���{�k�=��ѣ�*'Nm�0<66{��E�4.�˱�ϟI�f�bUf��TmCu4�x�ӳ�V'��i��k�N��'���Ju�_���?���^����ʞ�.�]�fc��)��%UX��c5�ԩ\c`���g8)�R��>P
>im����X��; �������r�w^p�egΜ��?��H!w��>��_l)���l��?��[�<|���_zݵ4�6���H�{^rK���!3�w�.��z�-�*�aK'y/}Ed=��k���H��憡���СǎM����?��Ν�`x]�g�c��ҩ
���[�7�׷�퓟�$4�׼��v�]�7aKR���;>G$uj�K�;�H��5:�_�`T��	� N��[���{F����Vk�,;�8A��r�k�ӫnڼ[������]7���~�!����I�́�R�?�>����Al�Y�ڃ�B=�֨�r��<�.�uT�?'��6�w�~<��7hW�k�K�4���OB��7�(�������ν�à�
��?:l�XJTwG�Ζ�Y6���ENh�?��n��u��Bϲ��a8s��]3�G���G��dM�1;���ypNG�ے�`g�*��;�s�{�݅�|���O#���(r���%Hi�������|CE�l�Jބl]qW$�������P^�����rF[��=�K�]�D�gY
r[���c/K���M�-�澟�q(V/K}���5��!i�:k���ۢu҃�~�"jL�Ѿ�*	��*�����%x$�ĹT�n%��n�(��bL�,��sK2-��(U��Ʈ��#��X��iL<I�.�5>���qq���9�g$���Ͳ�8'���2�yd�¢(Y�����'P$��'�6����J��&�2'fJ(;� V������Y"�v���U��F$2n��XS�/��
If6�v�����I��T�LB�@B>P��"��t6'EG
5e��VI"HLH�>\��&�:ZA�"k���Rs�^�``�A�xBqnY
��]7L����Ӧ��d+��Q��_�W�9���=�ꫯ���<t�P����������ёƜ��A��+�n�>�8�E�B-���l"�8E�&;e7[� JOǞ�J�q�d~��v[BA���@|KRS�KA,�I���Ǎ���<�L�����&ڃl#a0d�jL�_~���o���U�UBl �H�W0S|$���ِc����2����d%�+�c�WYI�%~ ���-63B�6�L�0ڪbs�3!����R�k�.���۰a�s��-��'	Y���~��w��]�}�kC�Ŝp;�<^N�xG䡱;A���]�'��P����ָX��:�G>�Jb��ڱM0E�|�����������~�?�p�Z�Neч�m�F���_(�k�cڦJ4�7ݝ����;vL��`68�Jh�$%1 ��,)�"Ly�#�	{��b �O�V~���q��]&(-.�yg�}-χ �n(]~���h�࿱ͣI�h� zɽ�[�5k)+�mw����"Im�w�%6��g�ބjg���r=�NavS�b���qʥ���h���h�z�n=�d��y(1�-�H�)�0��T��5F�$c��l]Մe�u�n��R-��z�6�}�&M�C���c��oP���[+�O�2��Md.�G�l@ƆI?T0���F�gZ�G�%��/(��g-�DQ�D��q�J�9�8`��\6��t�;��B����\��'��Je_�BY tS�S�9S�N��'�i����*B7�z�|��pϲ��ir5Mo.-����c�CY���D�(�G���K+����0����r��BVH�EK���G�#���)R�Ƙ3`/K��m�R����Tr�;4��L&Mճ�NƦ��r)cu�nJ�4\&�_a���]8�J�N���E�g���X��HFT��m狹B���ɉi*�Y������9ࡑ���u���jZKQ��� zi;��50���V��U<=�)gS9/�W����O�L׉
��l���UƘ��)��������
����������E�a��]7X�5�A%�_@t�S�"L[?�f���v(B�k�Z�ۨy���Z�4ߜ����bh�t
3YZ	���oۻ�8���n�v��e����� Xf�d��C�t|�Ov���ˇ�$d����]}�s������箻n�����o�\�TtS�����N6a+��e�5��L�)�P�-��"&y���B�AȤ�-�v`�y���٪vyg)̯���v��h�`Ρ����>�=��|��c=���Yy_��Jsyl�4O��y��AL���v�[7�y~���P-�F*UC�6T�:������\.�P'&N�ܹ���^#\-h�F8`�k5�C遒�8����Թ�s�+�H-��!z��(��r)��䂣�`lR�7R����s�L�Q{�G����A1X^��jS�?رm�eZ���ݰ8��iègz�������n���{�'~B���V�?�5L�0Td;m`[H�Q�
�i"m���.E֊%����.:�J��y�f�q��?��� =�ĝ�;���K:�v��kR�!���3�ybb&�ؙ������p���Q���V�K�a�й��Q�,+�F������=���(i��B�?��O�D�� ���O�,����U��'pI S��;�.mu���U�zۼy���(��<O����8@q���P�a���lM��#Hyʷ9m�����juU5nx=����n����ђ��Z�����(�-�M��*��%��w�!p��i�%�<����LL|���/EP����VN�ia�9�n��-*��++uq �1�H���8���ĵ�>����u��slЫg��ɐ��R%eߔ��#mF2�(�q�\[?��иt�
����U�t�����g;J}�T�W����N�y}���Ֆ��8�&d��AB��1ɨ$=��^m�x����NQ̵��?չ�$�6G��!OfL?&o�E�X�<����}jm�s�N�60(��B���W�b*�/��������8.�$���L�R��R.�'O��~��6v�nf�A%��ɟx쨈|�✔��)2���_e�1A&P=�k���O���i9Aכ�"��
N��<�C��Q�궰"Ф	|�3���z=lM���w�X�Ruu�t��?�Y�<xp��8��W���\LDy*)��=z��H��|h�yB���q�n�8��̰�`�I��S%p+B,]�����>�b	3����j�L��^�#,�P�L7ֹ�dVrκ�z%�+��~�L��Jޔ|�B���m۞\:CNM��M�棜#�����r��%�V���K}(����?Z_? kD�Cf��ԧ���72�Q> J����!)J���w�QLo�֭�CC�v� � �_�s��ր2�.?�g�g���]扙Q>ϛ�x��E萢�GZ�n&�d";���H�����ÇC�KP'c�p�r�*S���|�D�#�y���xg�4Y��H=�C���C��T��pva�Q�u�����p=�B�K����ɓ'���;���y�YR_�ÎH���,��K�o�h7��)��*s�,K��E�Ԛ-�8�\��`�:n���΂��q5���5���1�P+�2��̺J�R-��Ź�#G��ך��r<�G��&jM
���E�δۋ��ԥ���|�P`1�v���j\�e�j�M������ÀQ<�-�&�3�4���gHSe���^.�`����j�X'3�TR{9\�--j��ʗ�\��R[B�S�>b�x\�a��i�ZF����P]�{T����V4�E~T?��s��p\B��a�963�|ڎk����NDl��](x5�f�q��iCK�3�R#�.����d[��D�nH80�.�Y��ؑ#����@
�bz�V��EJ���d&45B4��껞��GƓ��A��Й*tvC��q����a��ZF��"�:@��?`\x�>#�o�)��9�B*ݎ�,��V���ڨ-ճ�������6`��T�&ㄙ�'9G�oZ���u�����ժ�'�_�/�l�7�Ry'���:gm�U�R�tnn��jdsf�fQ�Ih,.�
�vہ������)َTĨ�$&C>�#����ƥ�s�KlM�+)t5�;m�
6�q�E�)�hy s��c���-)+�!�O�B���j�UF���1-��ݶ�����+��Ny4k-g��v>708\h6z�\pޞ��3T��������2�\M� m9X�P)��k���J��(�
��z��X���Z��t�:�{��d��v�iO릳Ja�lvWsԉ��G7����k�]2��i�BW�RF��fҶFg��f.Up�ݔ���쩩)U�/{��Ͽ����G�V3���������/~�/�{�>v�?}��������"���1�7==mps�n7���Fl{�P���&DcZS��"Z~������B)��������0�Z)k�N[6?%�`R����o9�$�łU���Ǫ܃Gg\�����X�[�~�Kk��\P���y����l(�J[k�L%��Bs�����^�~�Ã�x��Å�:T$��T��PВT�Ig�Z%+O�~Wx�a,�Eeh~���NoZ�f�E.�� '�m��B�c�+Ns�A!��r)a�L៝�Ņy�΀)��t�UZ���[��&Y�T������~F�`
���MʀpA�&4�Ӡમ�ֳz�k �V{�:���[���8a����^�'*��d��M���r���;[G6c�Bg3�f�?37m	f����W���fJ_�cǎa�Iw:(:�N�"�V;��T$v
TX�]�SN�������Pr���GIļ���&�˵�@��6�O���̶~�T)~������y���sC5nf�U���1�	��.���Zv*��c
:NK".�O���q�iv�SG8JcVN����Z�`��fFL���I�\\9$�!o�1�2$8�t\��\�ݓ�F�#&3#��j��&E8�����L��e�GI�)X�'����P�$�,��x��[Jm4(X���I�l*e�n��:[�����w�#5b�%.	���5߬�7���x����RǊ[�uԳ���7�b�dk��Ǿ�L�!q�I _^P�a��r>��茉*�֕�Gu��H��6�y�g$މ]�F��U]zȆK��rJb�B�I86��HO�\%����	����Hبʁdb�A�	a���r�j uB���nY<9Qo�$�����?������I�&�ك�����۸�In1סɝ�$�B��$���G3�h�6��Ġ���3^��Z�d �Ki�@;�H�6A��6�(�����5����e�X�3�z5�<x��n�a��f�Ĺ��o}�[��{x���0u�9r�������+.��54T�.yk����A��4�gK1ڡ�}��U0���l*I�w���ڞc,%�#��XS����a���N;��,�1z���.=�q�f��k����;�O���h�����g�(q!�c~(I�_��޷� ��a\�"�W�w�a�A\[�05J^�\�+���	aKr����cL]K�1rW�#�b.��83�7���d����_!P������!�������")��b������Mq/()k���Dn�q~Xd(gɺ'S�(з[�<��k���A�M+p֩��Y�;B.�8�r%vtk�~4�$��P*��T��u��4v���T�q�����<�Z��{!5�ڑ&ޝ�膯�<Mw:,F��W�t%����|B�k�I`��:;O�5�FƬ�LH��@$R���̴@+P��NK*����;
�.5�<Â�t�f���L%�}*�RbG�����"���6�Y�ar�QA#�F�@�XD#u����ܠ�l��5DQ�|�@�Xǎ�s=��@��o��<+�TXj�:��q/�^���ANz�y��]�ou����t������>�#)l�*�	֎��Y\ڀ�H���6fy��뵵�j�L@�U,糹
x��䤈�G�T��s.:�$�n�!�n�ф$-V �h�*d��L���"B�b�)�ݧ$-�[�D��[�yS8�(�T��+��ᨭ�K_�s� �:c�&A��#�miq� ,j�h�8�`���ɭ� Q򫐜��$��oj6''1~;�OB'�b�T*a����*�9m�b9�[�\���T)=�"�I��g4:9�F�lK��>A�Ax�*�Bw����v�fH"�S8{ue�R,`���f�����E�ı��=P)po!�U�l����)�g��8��s7��b�����b)C6}���տ��/�Mog�~z`��j����S]�"@R>R���T�U�Z�	k�/\�?��/��(R�D��"(�1�~Vr�}�}�FP�<55�%;�,�Z�f�_YO����*xB3�h%<KYI�D�
+}R�~���Ϻ	�/��f�I�4?�<2ᔳ�TJ� �ҀSg�I
MT�uB������=91Q,�1�^��\+�D��%��c.��%x����w.7ʓ�i�C��E���k��t݅�*��D��^_�����ץN�d����PPXU*J��C�6QVñ��
�_��W�����G�G.��Ĩx�|t�dޱESI���,V�=Ha�R������(��;c�����z���"DŒV�Neu���8�dP5�i�Hf�ر�O���~}fJܞX���F�>s����`�v��%� e�ɞyJ��H��,O�\R�3�r�GlM��r�zT����
����r�Q�jM;R|3ˇ��
��D����gN�7�����*�sSl���r4�rL��و�#d�#��L ��T�/s��G֊����xAL�rDK#�;��GfҒ]���=h�$h��k��|������0����X�)oP�ʕ~ARI�q�{mf�Lۊ�����?!|<���D��p=��:�>;۠T);�#��&;H�w�l٢k&L���jcʷ�X�LI$��=��U��H�
�fg���j:Q)���Z(f��BΡ.d6��l�,�d���]�pKq�H�t��l�A�K4��s��ؗ&��s$J,~%�F��ϒ}ö>����a��޽{�S���'��gNM���wl%�O=)�|��g?�_^��_aX�w�~����|��#�ˬ�R|r:���� �()yv2E�?�>�#1�d2e3v;R���g�3Y�~�,3������P�S�_�"F�J��[ҭQ�	y��wy	b�f;���(�GQ�dG����������sj}�1�Le���C���C�K�4�O��xC�B�Uc{Z|l�w;����%f�ˊ�|���y���Lv"���%R_�������]M)�Ը5�8���Cd��LXZ�	�?��lA���?
7�Zv�v
.�)=ˊ�k��2�<���q<[;�J3�_%ٟA��=�8;��z�7���L_Dç��Ə��L��pU.K8�kkp�������#�ˋ����6�c,��0lg}e�aX�'��jqJ�hv�]�+�T����{b���XƵ���;q�Ćd��QG�w�" l�.���ӳ������R�:_I,�d7�\�'�Q�]C���:�����zT젗�d�0ǫIN
���>���ָ�n�>}:�rۉ�ˬ�/�@�T�)36�	�h�c�Y�@�b��	��x�%�
i`��ꑟ<�*����m�,C��Eͤs�q�)�O���h��T+h�z�>)"�XW���aZ:^�j��T�d���Ʈ2P��(�"�f�.�'��ow��D������vK0:6X��3Y���/8O4���&&�Р�P�T)R���h�q�
�LpX��Xc#,ϐ�����.�u�h�'VƜ(R�o�e`KKKw�Y"��.QT#r���ɏ��
�Q���T�)��1kdtPZ��^�J�*?��T���r�����
�R���"�G��Xh�4;���VH�%������u]º��l�.����̘QL0�P�1�b����"z��7����k��uzme��t[�Av	���}{�c,�3��a��&'~j��q�ƙ�i��vl�NE@#c�~���fg��mo۳w;uj�0W�L9e{�����R�08���A��z������x�c��|&�//"1别0-'���O�����g��W"1�.����rWC��
e��}&Eb��b��@�x��[O��V�w-�x�.bQ���s5�l���J�Ox��?���<�Ou(}��������m��:����t��a�l�)�� a�ڍXT6~������ξ1-Z�_���X�s�]�)cJ����tn�K����Nba����b{5�>l�(_�QV����R)Z"�����b4U���g��*}���뒂0>>~�&�� �%�|]q���~U9W����)}��|���L��1c�҃\8��Q.aN/I�;_"�G���n�gA�Rl���J�)��2��Ï���\���3�t��2<?��X���:u
&��v��Y��@iT��W��o��$���-$�#���˲V^A,���������4I�l6	�+�?������^e;d�֭[7oތi�ο���ܹ�g����艽2F\��$�	���noO/(�$�`���&@%����36��ú��J�xq����دUUXefe(ňW��!,�u<���M�&�	eqSҜ@�j�&���������{ފ�xb��IQ@� z���dV��v6�n�p�_�)"���H��z�[�>�/�E�R(*"�>Q!q}�����1�7��Ʈ&�ڴ�������q��jQ�~��JT���5�������'�Z��!���Q��^D��y�F�Nҕi�
5������@7�7����+�8�(�{��f���Q?��Kd����;c�fgg��8?�T�r�J]�]j�q���ɋ@7ڲe�{qeY�-I��ժ�juxx��:��qN�eL9P�j���2%D6�9R_��Kd�$��_n)}�_���gI��O��5����`��q\_Ucՠ����3�%�Z�+���Jj�x���}6�S���g&�����]�>Ց��F�*$G��ݗ ��f�ɳ�I�7R� v�� �����u���,��|}n�Г*���\�q@��w�g�J�xz���I�l�D	�Vx�L�A\�&���1�9��0`�l��YoP�_"��3�?�s������*P��x���m噎�]
2�R�����Pβ�Cv��+I��W}�h�<Bi��u�|��֛�n+UhR�Bi��/�~� q�*I�M%!20��PXl�\����縺aKU���m�2v�N���<V���2�N�Sc_���u�H#��no�F�i3,W�"ٽ�S�L��$�L���G�/R*aMNN&k,r��:>����j���,-�af*$'9&4l�D��O�t++i
"6����0Vk$c�A�*=T�@���p�u��W#��8a������rz�l8�ϑ�G|ds��@y����S�f�"��fc�լ�K�B>g�F�h���
� �`G��p����G��a�ў�%(�����j��q�2f��>k҄D���(&�r����v_^�F���
����.>!!I���5\q�$�*"�S�|6�X.�l�z$D�dH��fX!Q%�X���>b薯�A��;�	B�P���x C6k��Po�^�YO��6��Ru:?��>h�&o�@z*�w]UZl/*�p�f����2����P>`�)�x�:�#��mۖ�ل�P[������"���,�9}���Ҧk���?^�:S;]���yKssx񌝚�<s���-۶c��;m[=�3��j:t�	�`��ݛƷ>|�?��+�#��n�ݻjȣ�>z��D�떋�={LO�ltz���P�e3&ǀi���P��=���c'v:TΖ爴dK��9�����:��:KE`��a w� �T�gLXM"��=�bp��c��/
i�B��'(��8�֯�3�~���ib%s%Sʯ�rj,� N�r���An��K`D�	lT�O$�&Ĉ��H{,����.���n-�:���>�z�[�V��/�bH��b�I�?��^���Z�VT@�D���Xr�IR.�&1�] ��"Ԯ���	�3�>c��+�I�'����4�1�K�9e:<��Q��#R���a��u�K�d`A��D�a�W*����b_T;�ۦ�M��lK����%�&��#�F���|]�"�F�XWI��G%�n3�f!h����7N��h���%w%98I�N��Z��Ͳ6�ِ�r�����h��&P!�E�ĭ0QJ�-ȅf�/<n۬*�"3�!d'��d�d�����{>��@�LOO���e����4B_�_q�	A�Y��dB�z�U=Z<-�kw����p��8uN�u��v�#�
Y)��>=UZSCȌ��pl^Ѽ�5���w	����7z�����dW�H���ҍhJ%HISg�[WAn�ئP���ЭX��h����)����͠�!G$�e�m��A�4O|������>��q#���E� �8]��u��d%�W�����z�E��:�~b�5��lN�:����qV�M#d��ڵK��/�}Ju��"�����Z��)����Λt��A���^=��ѣ������K^����������iz��_��hN�rg�G�s�I��X��@bx���oɂ����%��+t�8��|�N����O��]DDն����X/�,�M>���-�)\y����~5����_�;끀~U)\OH<+�/3�{_�c�a��p�A�!fq�?�=��c_�����ӈ���ǃ
��4Cټ��:�{����8��H�HW��J���t�1�� o�^�Ʉ��Mlj���'On޲I��(���
��R���LXz��ˇx����b��@>��"�C"���0@��H��=�"�����I������LZ9�$��4e��t&�"i��t�~S*tC+�)��F-�'3�����@�n�N��Q�4fSv,�/�Z_��z�z�<�L��r��ăZ�&s��z���'��K.�L�l��ND������!�͌�P�2��Ù���u�L����(�-�eI��L�|�ΐ���iq�����% �����Y�5FG6������AQ (X�O4���A`�L:I͓�3�5H:�/L���8�\��`��T�$�3�҅mӔprr�T.����0����/}��ϔ.//J�Q@���]0mz�^��3�<4<��y@02�&��0)g�P#㊀�n��.��$��O��۷o�fG�k�>n+ގ�rO�T!�7���v�p��ԬQ6�R� tS���YpG��|�=��L��Է�3���hST4�F5b���LBK c����DrPpb��׻�׍j��i�?��,!�l.M�����0-��;P-7m��+�Ϡ
I�]��Pw���+��S/]G�ဩ�"�~���`�֘�����߰aӉS͎�q|3������AX�����5j��|��$n&����m�N�]L��_�v{���\'��{��#�6U�C� �ľG�Z���f*���c�`�@���e�^�U��>q�ĩ�g*��{��ޛn���믿��GFF.}�������\��~���/�d����ή��{���C�kN�
,Ia����C��f�AɶBmg5.69KHK�e]�a)y��8R�`���@�b�H[��%=�\���%�[ ��#+cP㖹ͱ�]����T��ʄ��t��s�1���č�X&zR����H�xK>$���dO�X���#JR���"��U��+�����R
U�`�0Tɓ�v\�W18�a���Q�[��D�*��]�n6(;US[�����!��m�Z�O t�aJ*1[$���Xx]�K���J���F���$�K����@~8��
K�P�����1Y�m������Ǜͺxs%�I��f�!�[�Q0γ!"A�^ q�3g�����m}m=.�}Z��|����1~\��S^���Y��\I�=��X������&�S�{ލ�h2���G6�%ra�'�D<$:��GJ��TI���N��͐8�덆�@ial&�%�ƌ@~{���Y>p;�h��GU��z5�R")�c�}�Ѥ����"�$�WP�s�7��	d��K��!�$�	��,�m�1�Yq��Y��j;�������wά&��9�wÓZA�rԳ��B"�0���*�$�<y�8f*��K2�Q(�G�)Ƴ�8�{vǷ��5o�3�U$��i��c�먜���p�.�`ZzF��֍�m�?�8<Q���C,-/�R�e�C��x�
F�2��/����0�" �����(>��G\���4��&�Lgpjp1鮉b�\������3;;�����x��|饗��)쑂�m�\*�1��48���P=uꔩS|{���Չ�����̂���O�՛X�]���|��/{��9�qzf�뮓����7���B=��t��Q���ݻ7�;w�uW�A�^E�7�9�e���~�s"[��ݗ���=��t�����A���>�G%2F;]Y�2�b$;�׈D�]�ĦK��Wϋ(q.��� ��� �li��-��Tv��\9�N�v�`��#ab	����L��e�֦�*I���"�u����ң���UԴM]YnP2(��^d�!Z�g6��#|�b?lRAW^�gEf�O�hK!(��8��Y\�*'_���Î�V���r�<s��W�ٿ��(�B�2��+��7O?k~:�������6MG���7�0���Yc �l.��穛!W�!�F�6��Z*
�
�e3Ň�K���0F�U���4��9�/p�5&q1w�w���ju�;�^���:	��뤑ѧ3<��89!EP0YH�T'�E*).*����� 0��3}�Ä����M�81K�F�/���'�0-�"���Q�$aغrèc�R_3%�(���P�˄������.�f�2�\Ɍ=g��)�,��~h�h���\�I#S�mU��X{�8�ko|f{�U�Ւ�܍{Ŧ7SCK �� 7���{C!|�Fn
� ���1�q�\�%�K�-�:;����ֲ̌����oгޝ�������;�9M��sx�E���By�R�Faj�~�%%e�ԧ���p%�+~�MT�`M��e�T�Q��v���`oG�J-�}�`qQ�������QW��2k�t`!�I	�'#I5%��IX����ܢB	l�b3���wx 9�G�_q�뜘�C!�s��˂vt����9Q�&�u�3HI��b0QV>�.jS:���i�Å��ꐓ"����!;ݎ�p8XPl�;ã�M�6�hj�*�X"�z�5��Z��뿰x�⡑�����̆PA���^�}�R/�9�NϔT�`���9����#@�����;�J�J�щ�����Am,֮�N��ˑ]�HBu��e%�/��o<������|���8��ӯ���D���⒪��'�G�����P�E�1w�c��ȕ��u��{O�z��(o�&���!{Jf�J��Q��x?��"��bɻ,��T""M� �(%��"R�cA�A����Vf�I6�r�<�ϷM�\60����t���,���Sޖ�9���RU#1*N�	U�H:�XEx�9M���2.�'�Ǟ����dS�o2#�Z&�m����>��;��t&�M�V!:�&�.ʚ��\J��\:�
C�h��6::���]|X�s��PD	'b[As0��1?�� d]q���	�K��A5O�u�t�\ϟ�)l��\����۫��'H}�7�lF��jڱ��|E,�PN� �;����#���r5J���u]7��q�����zsۚuA���N	B0��p�E��&��H�J+�d��b�����"	.@Pq���V���)�|N0�%sZ����i����c`MP5Zz0a�I&kB���+T%��\�l���Q�f�:��Sթ(��W����c��p���������)�2��he-�����C���M�����p~Coj�a�����{�3�4C��r�OV$W�*���Z�1
]�/'@��?������32s��#�$&����qΜYUUU�8.���6�E)�;0q�$ou)�Gj���K��9�Nn��8�6�LRCbu��n~QӑI��w�,�1y�fƆ�ɡ��:�
��5�,
�IY�Ky�;U�F��bM6b"x����;��	����ؘ�f�jnn�Ec"�Ѕ�֭���J*����;::S�u���m/6^�H;w�t;]򯭭���niial��b�^]M�E��P�Ò�^uMMgg'��Ϝ9�.]�t�֭�l:��[o}��G�-[v�7�t�M�~X�'oXu��g���;vp[B)-�[���4&#{�]�G����dsg}<�O;d�+��!󯢿����d�E4�wFtʖV�a��ʺ�.R^"B~��2&����z�������R?_4�[+T�U�ߦ�h0��B�<�,�ԕٵ�!cN��&�f�e�-[�s{}\�o��쮩���C��e�Ƣ8��K'ůX}�h�'�@L�Kh	��Ǜ�{�q�6�2AL��7��������;��X�$����,�SO�˚i^'<>�r��fz�0�cq�zAe2#���A|9U�LDS�sI.X���r���jn�!������V�%ӄ����lw��95-Q� jK�p��,n�K3�R�L�q��)�a�SWp�L�GO��Y��S%SR���*o�@N}��G�I˚��d����mzMo��	 �'u��-|އ���VTLuD�$��%��n���m���;]�J۝���h|r�HD��&�H���50�*�&6�{-+:܉�,9��BR��xw��)��D����h�4��ڭ����8�.��Nf�b���Џ�U.Lzf��4 ��a,�D2��DPq��L�n�L�R_%�($!%����Ĳeݜ;�p'tI��h�o��uBЧ~bV�J.�vd2�x<��3֮][WW���D�=G�v�����43%C��~���E�)�ut8e��U�S[:�MS�@�Y�9̫���ș�N9 ,"鲸�$<{_�N�2�fLJ"�+65="k�|ii����h8Ii�Шx˘؜D�5�>����%��Xt2�ԖS}���z#���\�j̞��2��m۶^t�_��5%奭�vBfϞ33�Ҿ<t� �����m��eUu� ���tV�9ܓ�D��`Ee��婮�۽g_EEEAaqx�:�������[��(��_V^ɴ�P����G!��??���+�.pU	P�|����G�k���gu���������9|���J�l5������d�nCI����
���8����"^����d�4��0M E�@-�CΊ[i**��r�Ɨ���֗$�U�П�h�4�s�1�6�5��"����i�Q�:mZ�1Zbw�[����bx��qB�xG�I��,�g匼
�cj5J��]�s������q��M�V�lQ��$�p���$�ϭ�*�������m��n���PZZ�&[S�Ί�+ִ�Z�O.��g��9��Ǘcj,�)�8K�z\j�oDbx��xg
�|�Q�������������(=�ڄ��S��cnd��6���Q<���a���y��6C�qҲ���I���XELc��#=�_�:$��E�[6����`]�?M%QWim:�x~�}J��(f�5f�P1В��+g��G/E�-f��Ў͕Ռ�|�����,R^p�w)w��lsHb��L����d$Jy�l��0W�!��t��*&q3�o5�Q0��{l[L]P�t�*Qؚ���9r��gJ2�젧[4S3�
T�Ko�N�i�6�(�ۊQ�N�-��6�������O�� 	{�g%�!�� �9s�,Y8�-��C���!��u�U�˴*Ԓ�G;�w���c���4)���t6�R�6��~�N,j�,�@��a3�C,��~4'��T��66&�ۄ�{��擇l��p�X��@$�tzX�ت	u�o�įG��׭[Ǖ&c�����իW�u�]��;�?Lp<����H/�������Yd,x+^�ȡ�t6)���T�\UU�I��,���!�Ƀj�*p��L2)Z���҃n߾�ƥ�^
-�����_���~�;����̚ݸf͚_zw�Q��,zg��z}b��'mE�<���`���r鄂����c��I)���g��b���(5,���v]42{a|YKޑO���`$���̭1w�12⸗��C��Fc]�o8M@�B$���ؼT��ΤXA�$�O0��f`�
O;=���P�8��D����?��ӫ���jjKJJܾ`<;��F���gE!���n�[S��/�D���דk�1x�5&g��r�e���ŉ1�Y��a�Qy�D={0j>�k�^6�M���|,&4#�bM�3���^�,4�DeʄB�)��<�zsI��t��Dq}ݡ)����r��l[�6�bNM�,6b`�Z�}�0��ai���?���)��$��f*Lܞ���H�ؿ*���ԕ�	duʁGIY2sy6�pQ�`�9+�AE�A�j"�^�8��j�a��j(��gZ��I��NG��2��P(�G��.^_t�� ���C%��T��z���gZ��E���(��"��y�q��aF�D��-+�,�䱅w�n�[x�$�N��ʝ�1;�3)�X�\ibǖ��?X���_JD����w��;��p������E��c�` ���k���h7?����73G�A�j�M~*�QA}}��ػw��=�!�w��U��ҧ��Wݔ�dX��S�G�@��"	FUd3LbD��
��6�C��4V^-�8_AdEAx�#�G1�Sb�0�������N�����%���� m.���f�E8��������~eE%K��@��C��z|��3�LUV�5�j��� �|����.]r���?��>��$�S'@��/,,�
��!l�Pa1�  ��?H���2��0R��Ѷ��&c���5�ŘϢ����={q�SO;o����@��d�Q]]YRR��ՅYڱc�ｷ��oRRRFJmF���������=kށ�^r�r�Y�hj�����c�cT��:� ?^ꋓ�
~����E���`�*��⛌���4*A��n���_$�f���s�9Ȥ.�� z2c1���`o���W���d�4R�/n�AX3{I��
V�Q�.�ƌjb�
���쐀!D�3��'�?��D9$�:�y<��L�FG=^WeUym}�XYB���#�mP!��GGqmA�PSU��L��2�kF��Y���;�q0����Oe N'�[sd��m���D��&D���N� �����6�pM|�J�����+7��ߏ����υ����{���&$�K3%$����H���2`�j$zȆ��":��(ǒs'y�4��cQ9�Ϊ	H�*PEN;�7�f
�������wQw��^*}�5��!n�g�OG�W��;C�i�H��o�������a��m�#�v�F݁ƕ�<
��S>A2���qr��V
4�g-�YҦ��M��v��Ö�iO��j�rͨ�J K)��8?�弜�h��X�oR��w����y�3��X4�|�:
��;/�(�"�L%G갚��v��1.�e�?�_[T�j&?��k���m�vl���H�Y-sa��C~�u<:AN���߀/DgJ/��e@���������b��'���'������g!@��*�����N>S8R$�g��L�&�1>�E��|d�`D�������E����k��}'`�7�xcEY%mmm-�A�b�(��P`��F���(���<���������Pkġ�Q��q+��޽{1�z���SX��W�|����bz�%4O_u��#��_��W_y��~��:b �g��s��r5��)�,��?6�L�D���%R&�|���t�AT����<^3�G��٦Y���cAi�8�2�]��&[0Mg�Q<̛H��R�\�-�<��WL�:צ���`z3����@�<'�T{=>��uNS��a'Q�u�L����/!ed��h�}�v�H5&Xk�A���[)]�琽�\�'�	��o7ʆ��������=�\��.H���G�3�RYY��̈*\?1�OB�ky�ϴU�Ɩ�K|���5����~Bқ��T�D�)�ok�}�V���JhZ*�oKˋ<~��حG*�+�B�|뜃��V*���H���pMis4���t�L�{����Zm��\k*��'����Xd�p���D<���<�Fr:���;�����z�QWW��X-6aQ�,�z�1f�e3����W��`�v��Z�]�`<<���*JZ���ȭ"PI�"{ޔ��IIēAB�ko��"�`���7[d���.�D5e�h����zVu��>�+�=���6ݷ������Ql��.2x{P�Z��9�q��vR6@:�jv�C�/�%�|�p�3D�����Z=�KƓZP�{�\ȔI��b����-dthga����iN�I�%�7Y��8����By��6�e����
#;ś��T�;:�lN�/z`����. ��wN++�9�?�1�ŞR@���� Ӳ:�$$g (����N�z�3g�ʿ��0�*������"����N��� �e��$�=�8����6!ބV.Dj�]�!Y��\Jr�F�'U�'��ܽ���ٴ��GF������d|�ʥ]tѬY�jk�	��b��ww�����PQ�D�%�a&��'&^����Y16�_r�55��#����"��YDI��\ȩF.8i�V��[9����Z�R,:�J��bMl�T�& �'cI
mF&�V�j�F��V���3���c5՞L֒Jg�.�H����-@ G�%�MBj�L���'��}
ߗ�X�{��������U+���܋�^{miaQ��e%Ei%�N��&"�F%�*���ɮ
�������́�!�I���app�H����f���	b�;<2p��k��5T�78 9���[SE)�6Yє������9���5tS��{����W�����h�T|���>���E<�f+)�Y���������<i�����X.+Y�����ъA�i�B�69��t���w]���t���c}R�����߲ET�Ж��홉j���{r�A�SE2��[OtN(�o�2�v�˩dd��#��X	B�k�"��x,M&�{[��4�p�҉d8��)�ƶ�jO&�hr��V�>�7���Y(�,D1�x2�$9C��t'�1�ĺI*��Y���@��ʁE���/+;�l��N�R�0 -G�a����NkѤR(��Y'K��t�<�x�zF�-$�r�,x�fw
*�(<2vqc'^�28|�pr }�^���[68�\6Z�(���f�x`U5b��r`�RV8�&�b�6g(H	�>o �D�I,H:�Us1��zR����$E��۬�"���Ʉh�_h ��(��ᒪ�
����c��73R8wT�V�UL,F�4�3f�'h��2Ar"���=�mj�s�dM
J����T��Lng�"�6^ ����`�@6� N��ps0��s��3~H$O���xq[6w=��!}3���KΙ�DM6(,++c��p	Hyd�H�J#0�/�ɉ��~iM����dM�,_����)`��ķm۹��y��B�,�9v��Dl���X<E ���\�����e�f,�Ke|���Y";dS��ؽ~e�G:�1J�Q���DS�4h#��v�+�sk�~M\�� ��{$3�b��qB�aרa�S������P�x�T�����1��2��@�ӊ[�z�jy)���}K���ld`���l58� L�]4�Ϛ9@8͵2�a�ؾ}�����I���O>��K�����w�2l
��|z3��eb۶m+���s�v=!lX�*>s�ʰ�E�b�]$�if�C��i�qUEy&�'/hy9)�ׁD�&ّfΘ���4�#��6�5g���-�J���}A��jcc���3gN랝�1�&6mڴ~�zܟ���2�$� ۡ��A��D�L���z�mC	h��n�-��n�m!�d\�RUU���A��fR6	���ˡ�n�oi��i��?>��5��:t���i�H��X,fr�̙�JK��0�&��ߤ��������T^E5)\��*�|�2�+�D�g;�(�������"��n!I��N:Ɵho�&-�J�EPT��$�	�Q��^78CJ��X�0환���g)y�3J^�O��
��I*6�F�S��>�&-����)Sd��
C|:�j������.�g۩zgQK~v�4>�3A��X��J�����%����̀�b ^�9�nG2���dUv�����;���+v���.P԰��E�1��)3/���۽N��iSd�j�op���чmڕ�����sK�Ew2���#�$~�]�v�t4�R�������S�AK7�IT������D(X\UY>sVKyy��l�p��0T�p��5>�Y'�����&ht��� &PN&��Nc�h�f$�Y�q�$0��$.��EV�H5Zesv3;�5l���>ۘP��
�,ף��'��aǎ`�T�q+h��p1*�T
[��5�B�y|�'�h�_�E&���?�� Y޳g�!��.~�~PQ�����ŁojkkA�x5�ŋ��-�9���̲ь�ď��ܠ$��r�� �%W$��I���.�2����r{}��AR�
��
�?�PY6���w�E cp�`�'�-!)2��Z�FO�"I�>a�I6hy)5�I�a��A(�zA�H��� �K���*�?��G<FMlV��P��
��>>6J� ���m.78L��m��4V�^�d���Y��=4���tv8p����:�aw@ S�oI�� .|`�6PH*�)���	r�	)C������٬v�5��c�|&Mż[�$�i�(���%�@w�,N�#P�O&q�*+�e�x�!�<t�U�Z�T���E	��ng�L����F5�'��y�
55ͤ,�l���]�l��E��@�C}��];�_���RHV�
{!�&pБ�QL��ٳY�Le� E���؈f���e��T���dC��jkww������<n�f���Z�`��0&���NH���|�,�����XQ{�����q�&���!{��U����Ѿ~��m�$��t璒2�~<��4(�I-'�S�=��os�ʉ/��,d�Y���Iǰ�)��]|�3�ťy�y	��Ȣvw*9�-��-(�=
R6����x5�ۋ�l"��!��\%Ӂ�� ��#6>N���{29��ZY
��G1Q���pQ�#�$�.�	K_6��iR��s��/�ҀD_,Z�x��6��wno�Js���pV�rF������36#�_��2j�36́`�'S�z��=E[�B�!�q-v�6��ϡa�&���%æ�0���a��ၜHE���Nt�*���A��xU�R?+Zy��!�e(�%%|ht�!�p��� _���6�v�Z"1�$�kmm%���(�ܒ%KV�XQ[S�q��J&]N۴Ȯ�텉�hv3���<��$I�R��WYq)�&;�+�5-�Cl��#&ɪFq��bۈu16ߙ���o�.�^ziss�9B�ۦXTX���y׮}��^}�U�rU*EXx��8cݳ�c��(���'�~���߁��d���X�Ż@����^{mq1=��R�E0s
/�י5khk˖-�]��YM�"r���+ĦJ���>�3w��t����W�Z���ۋA2�ƚΛ7�Դ���B��Ȭ���Hr�^�wQ2�� ���c�m���8���Z��WH��+爐w�ne?A�%!,��G9������n��ν��<$#�U��Gq߾#��`�/����Z�͎MLp�w�O�� Z�.�����𡮱��N(�j
��3�*�YV6�R���6TѪwe�����͛��[�F��	�$âϚQʴ$�.��9�B_�)z�����b�P!1�l�2�C�|_����
�d1�#�`���8�������K%�j������'��ɢ�3�,
�y��[���9w�i�sAX�[�J�W���I�l+��'xViee__�I�l��>�7fd`\{��eŦ8|��o����|�.�%&��'�p��G&�j A`��T��4�x��)�j��?�1��;sw�K>ջ��E(yxsyw��|�0�7����Y�>>p����QKnL�����F7�0�0f�Ct�37�,b�8�4�MV�dN�!�������l3�O�Ew�3h�ޤ<��@�`��s	��)��6 �̰c��C�f�������k Dh�;bO��������)���K��![������V1���}ܓ��A9�pS��R��1j�M��>[E�H��T�����I}��ȑ#�<-�m������|,�ݿG�璌�|	�H8�oΎ�����{��!f�y�[o�Ιg��v�J�D=� �t�/h��%<���<TRUY�X�0��7_ۺuk4:
�\YYOn^�����^��V�9S?�FmR^�gsw1�pā��
ӄ���PP�=�ܕ+�J����z�3�����={�͞3����o���??���A�N��c݂�B��w�K�s���d�3�8 ^�.���-Z�_�ƨ��!��у|:}k�ҥ=����?O�%%���r\h �I��Ϟ��*F{1s��Q�g���ME#/(Fc8_�:��A������~�~��c��N�'��?���#�E��0�����3�v��nh�Q���[u;ITBH�Iby�֬�d)��f3�x"������[q�*�3X�K�H�����+���#��-d�o��������*��3�t�<�ܤ��B��k��9:��ް�T�Mʨԫ���!��z��T�f;���H�U-��0s:K
K��&'�ȟ�؜U�D2�E���^Mvj���Ԥ��Pޘޖ���c%W�&��>�N�V�:�Ə�JK˳�r��X:3����Ғm[��
�@a4��,�]�E�}��0Y���<�l��,ͪ���d&IPg J�`�K�g������D�ۺ<^O0KEF�@�! �*+\Z��� \^a�b�邺���M���v�t/X��M�#�{��]�l8���Ɛ������/�|��=�%����-Zĝ0Y�C�)).�cG�'�ׯ��!���:��3��c�O���ς8A$����<ʤRPP>0��S���N0 ]�B����x*�x�n�/���ٓY�5���]��G�ף��v%�o��B!��餬�,��⊬&����r�]�
(eU�
$Z¬|�/�f#2��+�Qi%4?��\��B2n����V�B���*H"' 71.MX�3�#{=�-��	A�"�O�e�)1��-~�T��P)!�L'����\LU3 1NB��X<�A�DU�v���:���������.��k�&ӡ ���1���q)J�Y#��AZ���7�^<����`wP�$���/��A����	��x��X�� ��@&�,T�j��/�e��2�W�@+�/�>�W��%;��7�$#��ر�-[�*��=Ɗ7�^���с�g0����r�iV�����=r�x�'��Rr��f�D#X�3gP2�m�r~ l������W��O�cҚQBj��Me���/��9����}�Yg-_�������V����=�[�|���'-���~�W��I"���ړ/���_��LOZ�?� 7n��c6n�������܌�ѝ����¼{뭷�1�����H������~ʎ��e�%��{��wכ�O^Z�K3�޽�_a'?�
Zŗ�]v��7�L�f�P����

_~饍������^v�%��կ^x�y���pإ�� �(���<#�j�ȷ}Y�Ÿ�ӏU�D��`_����	L$ܼ�� 4wP�5�\������"�dhd�
⭭���}��_����k���.�����~"'6®]�`��qnK�#P��Gp�����8Ibp,Gg9�+j1 U�F��	�Bd��vZ-��,^������.X�����&S�Zl8׊����7A{xtmU!����y����gD
�/1T�h�����h,�AWi�-��e�$�	Q��k��DIZ���d؈�n��d03�V,���d���h�g�gΚ5�8F�I1�χ��� 髫�8��+++s��}��X%	"��&�l����0t��BE��o�[��'��D�/F��,�n߽����Ĥ��L��*�"W�Oqj��KM�mg�xM�5�~�há^1�ԨS�9�!f�9�k�W�O%l��ت7C7���c�1���|2���2ׄQ+4{�\���hb�ӟ��?�h�!N��t(��$������`�Q�o���fa�y-���9<�����b�>,��B�@�h��n��!�M�M�
���`�L�NUUv<�Zjkk��lj���8W��b���|Y��q	CqQ��y�D/�=��ܛӤ����ϖ95�=��˪ �<ᢜ��g���o���1Jh�<n�\L�[���7nē&��������ֺ��������3O?f���fr��Z
��ڌ�9�g
2Ќa>��(PE�`����>�r��ݻw��H)j��/�sJN���J����r�	��-�I�0pR2*��㦂���68�'�� ��������TMM~g��߼�]����{��@1�+���k� 

B��n��$�X�g�z��� s���o����͓A-`R��q���������6224��{��_�z��G�fӣ��`[���"p0��nf�IF�H:N5��|�y�C3Uiv!���ok;�x�uױ�H������f�,M�sw��7l:���/���ݱo޷��L�m���+�ɄEd9[)��D�Ê�{�jQr�d:��$mN����?�)%�"ln�\i͖I*ɴ�v�#�ܡCee���7kf;=��Q(�V�f��;;�-����o	���gl�d}����|�/~~�l�M�������N��g��)F6�����i<�����A"-!r��**�=C����ii������
�����&��56�� �@ƚ��>!*JEe�����$��*�J8\�;��`��P�nhN\tՋ/��?|���.trN���,���e۩j�t:�H$v��R"��H�š	��J��>o���L�lHP��ry�!?�	�c`��%qR�D�a����<�������^�/�aZ��F#�ёq\u���˖�|��w:;�[f͆t�� �}{0�N����tY����'�tRAI	�v�q���8�?f����
x�e�)�0�O=����D��shd籆:����$f���U�̙�N�SQO.�`�v�}``h2.+�ڻo�j-La�q������لSS3��4�-�g�K�7C*����,��/�=dFѳ��) ��B�9ɖ%�M��R�as��)Q��Ļ��SKK�^�Y4��iͤg*�ty����)ˌu)q|o���{�N������̐�-�Y躋a�O��i�yR^h,�k�����0aN�\T�\V���4�2I�3���6��Ut����#����� ��W���kZX��&����Z�蒥����Z�ʦ��B<�C%��\B�E��FA|-�n4����4,��=�bC��U���>_&�b+Q:�ȗ�lt)ϓ�Ggg'���e���'e���Iȑo�� (e���(<����GB6��Iq`�B�ǘ֬YSTXt��)�l}u*V���V�lVq�c��J6��3�<��gb{��-,�;�k��9%���<�0%ME�T�@�a�@�v�%�|�s��6�H$Ɖ�ѿ5�+������,p+����r��e�`�c�Ap�p=��s�tQ�K��*�Q��\�~}yy)�B�� X�����d	hkX�3f�s�٧�z�>���ϳ�J�sE�īD���L前B����-F� �iL���d`ł�~�_�㦽�|��J]��Y�j.��BLL�+���������p,ܿi�&���c�Tci��BLv@�A��gs*��'���b���~��a��0/���Mg^$Nq�#���E�O|�dBx@f��������~��Oc����}��k����;�,L#V��2{6���;X,��&�ྜྷ]]]u�e����@�r2MC9�uѕ�2}�U�`j2[�G�,^���~��*;h��W���4ؼ���3뮺����>�haЖ_{���r�fu�i�lQQR$��l@�R.�W�,anYE31,4�gћ�MN��?1o7mµ���0(�8���3Ϝ{�s��ٿovH����*����Ep�71Ǽ�&�'�kٿd�lF �����	Y�x1N�\|��#�O��0�웛Ac0g�d^L�@NӔ��㒪��O}�S�v�O� [f|��6����x�?MW
����I�C���=Ҕ���U�>�|�)�<�]�+�����,sp9��n�=y��5#��	�M����l3Z��T�nhi
��N��4����&e;��j��T�qm^��1�ݼ?;}�cg��I�̨)�i���!g��)^,�.���� ���e7�k� E��5P ?�O�m�3N�?��B.�r��t|���O�0�gb��D.��`����9�Ӧ��_����|��K���A��P�X�� O�;���@&g2'�i[�l��P�aX��Т/�>�6=H����k4 ���6)l��E|�q�.Y�aw-_���nfwO{[{��jw�<�Tf��Ҙ�rs]RRΗ����e�n��z�wc!O9�pyS�J��16DQ"��&{��t20����I�EܸqݪU��!�1�c�2e��)�Vl���j��\����O��!A��)�M��
��gB	�>.$���11���^�v���`$�|�K_�����w�y'�ܹeޚ}eL��a�)05��ܔ�8e\:v�c�ã�38��o<��3�Uli���l�����r�^v �i�=2��8"��;��|�%w��_۶�\�dvaQ���0��Ñ}B�muaE�]�>�J����qz�J� 䥰����Yp��$l���|���ϸ���RҜ�gC���P���b���i�����5K��@ d�X�x�ɓ�,��k��������~��h���fvک�����%����?XTZ[W�>��}�ȑ���^x�����>�TWU��G#���-�s�q �3V[�jw3�zr��a�02�x�i�Θ5+�%����H&;ΌND5E��F�QܬeN��ȡ������}�I�����o���Q���GCR���Ɠ�թ��T�V�d<-���-G�}	�7XYY�4�t��u(���
���@��e�~�!��;�F�"�ڼ��[`I$NlV(�����
-��_1o>�|�W^y%�!���h�"�þw��pݚ��	��{�vGe���°� �%�UK����Ѯ�J��|���_uhx"Xv~���9;v~��OB;y��g����s���w��VQ���G��OZ������q��?��=--3��D�x\Ұ%������p&�RG`4 q?�ȴP����vYT�@�dY��҄��uXD����pf�l��`��b~���K+*v���+�ĝ�*kp��#�3}��o�����-�V-*).�؜�%�M302^��H�ͧ���m�Y)򃪒�Q��0���'M�v���fX~�;�J�!�sS�x,twrw����xr9;.v{)ӳ�`³���۶mP栣���h�u�g�q�������>��p����S���sTbS2����h�c<.��a'J�Z��@�Ȥn����9a�Wx�)������ ��E �vtv�(U�� (�.�w�����&��'�v̷!5����J k���Z]���W\���C�c���T3̡��%]�Ϲ���f�X9��Ɋc.��L���>��@e���nݺ�[�fE�j�lB.�ey΁1����?��O:����,!����������i�G�Y%�ɍ� .H��*���8��b�S)�SR��HRÀ%Q��m�-�d��0A�am�<k�,����섚��( e��h4�W��1�5��'��GJ�c#s�~����8�ӟ���N�����z�-.�7UQ�t)��#��99��
)�^���]�v���_��T?�5`��Cn-Z���F��	�``tt�(e�xᅗ�.]z�}?y����_8p ����6P���Ɲ1H!��z�p7�	 oq7��������n����Z�pl��me����`B��:ڱY0�����{u�'OZ�����~��?
���bY4WU������^�Ж�g��죎,��JLU�BȊ��+W�<����u�D^܈ 7L��l�Bs��d�֌3��@ر��E��]�v��߿��>}��߾u�{Е'ā���z �m��3�	�/?i&�b��	"bbK#�Ţ�c�L��*�`�F���:�袋��\m�7,��ry@c4[K��r����.�C��ۇ�r������m[[S#�!ʫ�C��G~{�L���MU��F �"l8���7��LX9fr���.���$��(�g	�� �FP�0N����}��_��ZD#IT"̜9�СC�gc������O�	ޒ�81�ܱjF����1�����+���Kl�^z�s��106z�I'}���^�ay�s���n��=�A��dؒ�����{睗^|�w���/�ԄZ���bhB�;>@�$,Ec�?��9��q1����v;�q[I�`�/UPT��FEѮ�^f��K.�����Gb!�u�P!x@*����?n��ח/_���~VS
��Ԥ�l6	��u��%8S�#tf�V^nrۨ�ՓJ	ϟ��Mq�fTj4W��e�d	��(��C"�{(��^��={8��}3xfU˩߿뮂�SO=����<��EH9U�pM��!W9���L��9�\dό���	�p��@�$Z!��c�8He��ųg�IgtFΑd�?�:% �)<_\,���ںj�8�9����'�td�Udv�r�m�D�77
ai��b�x�l�q.�G�|�x�/V4���b�X'���ux�����]����xg�%48���b���K��(h�p�ݻ�ǟ9�����h�M7ݴ`�`����vc5�[h4�n�+ �4�eaye����{�Y��VūbH�G��Ɖ�ڀ��w�={�5�\�jՊ�)�Y&'��?3N�������ÜY3�z�_�����k`��ڭ̬E-�df��&3g6F���{[������޲e���s��F�%"�'���?[�t���lOlnn���7lXc,6��N�U�E\c��b�w�ڃ�ɑ#�X{�p�׍�.8�p_vI�=cM1�իW����}饗D݈�kHX���5G���9������T�j�#�߰a�e�j֬fszE�^#�F�q%C{><>*��~�rWȺ�ş!�.
��66��2�W^y��0���}�ӟ���w���c�@ST�А��(ȑԌJAN��#[i1�L%�Ip[Y�R]�f�[}da	ΕNK��D����'��`S��i�LL2��v��+�����D�ȡV�LqaQ$<���.\��$��w�ۊ�^�~�ߞ|��>r��wODcg�u&3��}ϊL�J"<;�թ�n��R�
�MIa��ឈ�a�v��҅"=,<�������hd���΁6�t��)I�{PU=6�w"B	q^�kh�d�"�,nI�Fl+����A�پ�pr�����ޞ�y ����<I��W�"`Go���Dt#��!�E���v�AQf����H�d����nF��ڹ0jwo��R�u8�$�	2��37TTL�4<�<��A�<���N>y���O<y<gndC]U��D��]k�qI��1X��hqV�������s�):�s��o�����v���>�`o_o�ܹ_��o�ʍ��=)ph w+**9F�J�⸥�e��PW_o�ѾE������~���毾�>����Z<7�M�d�KJJo��rJ4�t{	sB���O�Jq���"�d`l2�#+�2�Q����s��Q�-u"�9rd�W��5�1qz&'�=��E�5�A��_���"V�#���#���<���_���M��b�,CE��a�/H附¤�t�h���z����%%��"�U�m�`GԂO���{��`݃�*mxv�M�d��TH9g���|�[��-̦R���6����!SqfUgW{Ee�7����7_|�m���ko5͜I�E�Θ���"�I�f,J�b볱k�"�g6�!�1�����+�Y�����tz��e]�`��@ą�i5�����E�l����q~(�v1K8�a�=�ؔ�p~((𵤩= A:6��<�����D	�T��X��"}�1]���� �s��A.o���i��)x�W�XQZR:�&T�"O9%`��Rػ���-�=���,�2H��ee��.��O}�bX���-|������іH�._Zz.��}?�։�|�P�� )�p���P~�F��N9e�1�H
3H�<�񦌙��Ԅ��/b�a�466B���;8�������$�����紷www'W�Z�d�_�����r�uRnI}�?��/,u?ƀa0��ַ�?�����ӹht���\ʥ�X�d��[�ly�W�&�K.«I�( ��l�isӡ����֭�0�o�?/���{�7����a^�ʲd� �уT%����Z.���ի�K�(�.5ʷg���0��;��ч1ۛ/8o�������� TTK4�Q 2�;w.6��>��(����/������7[�`�P):� �G�jYɈ2LGXD,�J���t8L��7��~�&�����_,��޻�"���s���\�Y3g��W.G�[`g�"dL8L����G/�⊕+W���[���I8�];���TW��80{�5:�إ-��t��&$�
�S�YA��_q�ҥKkj�tJ�B,��AD^$j[��0	�PSì��Z)�D�H{���8{z;�̙��[o�p玿>� �j��9�g{9�c�b:l31%X�5y�Ԝ	�x�����;w��`I���k��!�t�j�BWEU0u5���4!ƪ��j4fY~�*��/��2l�~��?�#�� �N�n������P9�j
4W�ϊ�ǰ"\c����2��S��r�?n���>�9�����CQ��(^�5p�0ϝ��UR\�σC}���m�}�h�W]u5��w���C���up*�f��S��"spD�d4{֩���ʧq���g� Ɋ��rO� ^�SW|������>С�W *�h���	N�f�hxee%�O?�V���o�_����<���T]^�dj�����jt�ӌ�v)s�_���,P���R�&�1��x�nݺh���n�mን`�}}��O�t�lGGGI1�C`�`e1򶶶�ƚ3g>��O��߽�cF�{TTTPK!��E����+��<^b��r/����I�}(/�S 3� N�6�G�Ģ;;cӒ�K�����m�R�N*+���@fd�C�r�*�x*fKO��(�j���\�QJ�۬�vf�6��4�o���l}\��ă�s#}�q����p�d��/}	/����vvv�mmy����אI��Kg͚���+	]��Jdۄt��34�W>��������d��L�##P g6U��oy���\s��7n����:X��H����L��|>�$�%a���g?�-���$θ4xpL�.��#c�?��@��\y`��D�)C��*���1ku�5x�s�?��#�HT���@�nOs�l�������,Z�[�gτ�b�pƌ:�������7���+����?��]������M��RQP���sϽ��3GIaS8{��^c�쩤�������o��IX�z5����~�����w��M���e%YR+����XIi���ڻw��P?�?��w�o��׿��5(�!}H��J��1p�J����]�h����6���FX����ją߬�����j|�����������|����x�X�H�|�C���T����q�������1�̟��_�x�G���G��ϟ�¨lv9��X�%�@J.���.�%Q��Uv-_���`�\#��QbЙ,�%ӂ��n�T:���~��Ӊg�����?_YIr�C#�%Ed0Ař����s�9�����c����.���M�t���)��e��'"��`d}���r�D4U����wt������s��{\��+���꫃�B�kJֱ�AZ<�l<����ԴC��s����N��ny�ЦSO����tz��q�'ӑX�jî
-Z�~p������?��~�o���E"q�,�d<�	̡��>p!��ff�/v����*iP�����Q��{��|��H~�{P�wS�(��)T�7cTR.閖y�6�L~����Y�f|t���?����+W^��,X���{�6Q>S
<t�=�$�x���xeD �����dd`�(��kW�j��c�,͂�q:6KK��/}�󈄨�������LD�C!��/D�ۺ+*�D|9W\\
��ȿ2��-�w�܎5��|���\x长��}P�/]d�䒉�d,.��sЦ�Z4�������tJ!X�\�;����p<��ȾNP��g]���|�q�윦����*�l�ѱ�����0x�J��`��&�5���m��۠��y�o���+��z��loi���m���s��7sU�(W��Zك�'��
����1eb���C�����{��֮\�����N&�B�|�<J(,���FľX0.~ݱc'ި�����/���K����翀֋�<_,B%me�E\�ɑxI�F@��TIO�P��������F��΅�P�|�?��� e]p�y�V��D�C__/W�,��YW�D1�;�+��9Z�����Kq�?G%p^���0˩ �/b���@2C�'��?���-��d�����g3��#� �ê�`��J�F���:Fs�-�|�_`�ڼJ6:���d�R(n�##�����^z�0耰�d�a#�o���L��(lR4
����x�3�8�(����y��y}>�'��ܹ��΅i)#�MR��0̺u�.����cL�D2!z<���)2'*���+��?�� ��H���\�������|��y��j=1v��i]�p��xt۶�˖-��O��˯CA��j� ��&�����O������'�Z��U�"�ja���1�add�{~��ObQ�23�;':�\pC�Thoe�e��'�0�� ���۷�M׬!H�O<񄙧�g�ƱC��H~��@),+�^�����c���x�ک�'{��w}w���N�u��y�t����O<��w��k���#�,��I���v���7$A�b��eb���.��=��_�Ö��T�]��sQ}>ʆ�r�D���/9묳���1�h<f��b�(�븏;�h�ps��.Lŏ~��T:�_��71���
Q�X'e�n���)#*ѻ(c��^�~=��G~��{��>*)-�����&V�E܄8�
i������^{m�l�~�SH���YE�Q�7���\��XW��+������)P~ TF��lmx}��e��ϘL<kp�R������/8n�馗_~̫����M!ƬXJ�����Tᒩ��Po�������]G6��0}2��7�n��$��?�ob`{��*���W]U�yf��SG��5��[o��N=㌻�������Bz��D*���r�5װp�H��C� ��͛76�B<��ihp�w�ń_r�%�M$�h�Q�S�je3��B�c�B�.�^(F�Q��vd*��T:�ƛo�TV,���׿�5����J%�f����2Ȕ,!+驨�^�"�>,̠��4!�3�Q4F��+W���9iU@���jUI�����E�pKIj�V��:���X�`0@��v��꫰UZZZ�z������_�F�#��M�lԛ�`s��?y��l6�8�]8�l�p���3�t�"##{�D�Ȟ#/ �{d�-�w 20~�]]]���,XPXTqs�E�~��PL�g*�ȿN�6(�SF�6�ntf�	�f�Y��	n�Ǚ"�ށk70�n������#I�{�n����E�f]�dD�9��v�"gC�rS*j3����H.N�`ș
ɢ�+'��|��$BT�)�>�!����R��f�O����2����t�ς����Z����tl޼*2��ғVq��_���0o�#������~����t�I��U�O'|�A/6v���n�UE��u����ڙ��?��նj��%K�8��~����f�(Y��PM��������o{���{�1�:�,[���K/]�h^��m_<nj#D��fāw��2��h��w߽u�V�cT�#[k�"��填ꢅK�ڿ��m۶A�hl��{��_HYX�g��ׯ_�jՊ?��O��Xc�J��,��G0 ػ����H$��. N��^�[hpqJҎF�L+W.��������=W�9+�:��'����f�UW]qe�X9�r箝,��W@%,׷n��\E��;�|�}j����~�����3�8��o����8�#d)AI�9��1`bo��VHD�˾x��ᱡ�ÇʫJ-�3��?oz���o�{��>?LT^,BT�������~p�7^��_�n͆M���O�<�4���vf�S�D���	��$�I�熆�/��~Cl�Ҥ���h�0T$[<� 񋱱��¢@AQ��0N�����=�ƛ�UV���afl}���f@
JB9��ƀK�#��d���6�8��Nl�`�����g���3�������~dw�[���8#9%��j
�)%
��(ee�[���_����J���ll��3��'���G��m�;,�����������1f!����imݾvݦ����:�\.��)K9g(X9��T���;:[����~�{~���}ڹs7䄙�,Ɛ�P�65���jAQ1�㮞N�S]�bŊ�Z�7x(��Թ�rM|^�-1!Q�E���i�c�.������A0Te�S�x� .mC;y�g ��ܼ���2�������D��oix��7@�\����i��0	��!T����== `�#0L��Dx���8��W����� n���E��:���{�l������;�&�	M�F�Yu">QVRTS�}�-uUk�m\�n�}�?�;��PQ�;�N�H�T�S�B8���L&�mv�Gʄ�>2�d��x�u�P���X������q���,�`qUyX�d�545;��bw[wR�Q$H���@?E������x��K/���/�����E�UPX!�p����c�h:ڠ*)��r89����������W^��o�}V�B�J����\H�^���@�Z�'�6G<� I���f0����2Aǚ5��́�C���M͏��ѷ�y���w�]�~��I+U��U\mȆ8�Ȝ�����3��˾RSZ����gΚ���4c��K"[���q��#�,��z���/�r����c��P9�H�p&v�%�<<E�1`D�Hz
��8�.�u��L%��U��?�lO:^�s:.����uP�׮3~�gS��=�lX�gI�����㕰Q������55˖��q��m܉(͠�C�������(i���p�H7�g�[XRbR�Qً���:�##�ۼ��((�`��z+�}�7u�Zø�<v���������1��1qI+/�ܢ0V��$0>.Z�M�q����g�}��9q�MS��7x)�|�k�6�`K�q_���N?��ixP!��<qB8�)����ח^z�g?�6	(��m��cv���&:�V�Z"��q{��ן��$\�x�bZ��$��EV\�Y��#�����+���`����Lcc�Q��(�h#�o0��ǩ#�]�v}����ɧ�����Ut��V���h����ۡ�\vŕ��v[]M5��+Z���f�&7<\ �\�bŏ~r�_~�_�>�5�S3��y��o˼���:��!��8����(���> .#k�
����kv�=�܅��:�<���5�<p�G����k
����D��{0�#�Q+W����{/��"(R�����*��k� �'2�6�l��;.��Rc�iJNe���S�,�KE����s��:/����;w}vPBg���1ɘ���~�r՚Ӗ/_.[)*oӨ���XL��.�/�p��P!7lڴa�ƿ��,zgg�G<�1���F�S���z�|,��v�8�>� �@u����E^B����"ċC��T^��K/͘1jwYiY�쥃X�@�7��A-��e˖����s��������kϿ����C ��1FI�҃�1	3��!���CKk�3{p`��47n�Du�7��s5���!;)&DU�Ғґ�|����]wݍ��?�"ca�)q�������F6���x���������3N;��G=t���|nfLIKf��&�y�~�1OD�]��F��_{���uxVV��G�9vSE�ǎ'���h����A%ۿk/�:�Z���T���:��h�h�
�7(
��g�����+��뮻��Ϟ=��9��|1�ID v���R���eL==����>{��L2�36:N�"���ύ�\�������*��ϝ;g��]I�N�|�֥���G��+��ƆF���۶���?��/~1o.b5gR2 Z��<�Lfb
��YM�D* >777C�tv�p�T���4L׌�:�cI�y0jF1�D�1��Eً{����K�D�Xk�w�_�q����P��pq&��a��af��vH{�� ��mpX�Q�Nxsw��b#��(i��xX'x��q� ����!�^�����=�~����A�q9� �i�+�Ɋ��'u'�����fUJ)�dYU�6��'��s����|��DB�]��=��~r�ʥ���1=S	����w HU_{�2�o/�.�²�����(�^>[�11Q�&Ɩ����φ�Yb7v,(XP)�a��^���������a��/��ffg����?��,�X4�Lȁ@�d2O�2�����s/=���ﳒ��ހ�9	i#O�T9Aլ�M��0�w����5k�����]ʏ��������j=O��q���N��s΁FD(�OMF,@�܈����k�p �Fyݺ��x�	p�A���B�AIg"BG	('
FRI2�j���_s�u0y����xTv������c�z��H�WT�K �M$gL��q���+�
� `y���/0����8U�d5���qC>W�&O|��O?�4�3w�<�@�(�E�1��QT8��6U���[������7�|��w�I��1t�d!}+&D�TV><��ow��+��|��?����ν���>��m�ǎ�x�m���`��U"�8v4�
G����zr��7�H�"Ey9���/>w��w�0���첛}���+�J`X��H�U����
�*=�Ԏ�w]}}4�0��XGtZ�������?i��s�����oq�pղ��]�޻����_��s$,o޼���SO-���R��!iI�K$�=�$E��<Nm`�����n�]崻�?�
���,;���F���}�|���ַ��'�mx��%KG�i����b,*2������bQ��f�(������������{�z��rE�1�D�#�)����v�\��KA�*ܱ�z����Z���&�%����p�s�9]��#G���ܘ��pv�&���r�n�����s�̩����q�J5�>_(1	ȱ�����?'��x1~(��q�sܒ�Z�ɇ��pyr$%y�xˡ�M�]vYɰ�m{vU��+V����mE%%^?�aqDFt7FXL���P�g���5�����[u��+�^]]�p�<����7'��Ɵ7�����s<}a�����{�
���(w��B���p���_�.T�`�j����`\�s�ޯ��GbyF�dvok������n��o�#E&V����7�n��q<��*�J�s*a��Tw�׌���{߽�~����2�}��?��'��P�g�iim��_2l����� �W}��8�v�3/����/�2{I�T�"��&)��fU�jQ���&+Ç�6\���)�1.��;��hD	m~0�����Z��b�8
J&%���V�i�4����ԛ��Ӹkɒ%_r������h*�F�x���s�a"�����	�د�뫮�
&���ihh�����v��2���L��h8�N�A�T9��ʥ�q��h�@\�[�}Iii ڵk$�ϫA�BPK��up���n1[d�Y
���*�vv�c����v���M��B�p�@NN����`�X�lmo��	I�=6	������1j �c�ѥ@�������Ic,v�੎��q��K��t��='uƤ�D��k���c����MiW?�͞>��Sy��>X)|e��C�w��p?�D�ʾeE$�
{�i�����j���PQ��CG��Θ����0�"c��t��T8�I���LJ�I���՟����6n���!"�`b�J-J��V��������N�m�����ضv��)�ﹸq�&Z/\{����(Պ����>������Q��f+4w��7�lٵp-b���Q/G�4�QKq	. �P�5�ڴ���o�=�\��f��qP�6�C~]h����f�;�<��kȴ+LW�c��yj�01k�X��"̲���d�ĉ�ak�z�����N�BM�t�t^+9�\�4��{��^��{cƌ)��O�AH���<

6��몦���?�����V�m]z���p(�H
ljj�Kll3ቭ��isfa4��|u�`�~��\��/.���
PC ѥ�x����?Y��;�s��~���������ȅl-��F��믽��?�����{���⋰ؾ�����s4h��ሀ�Ƅo#*,Q����p�y�̺/�`��ꪄ��*gzp����_��0�O?�t�֭.�i,3�F��4�]P��F�����X<z���W��8u��G��*�~��g3�b4�p�2(�������B&~y9f�֛oB�`\v�X�}���"�,F�&X��9�j��ۻW��R�>��\xr�����6m���;ϛ7��x� ݱcn�L��qO+��Skko��1�'2C�D5>�xfΜ��8 %�Z���n��:mr����SynF���w�2g�y�W\A�l�dQA��U���a���zz��R@ /\����_��[`3A=R�o��(g�d�~����`��/��M�@� c��<q�����6�#C�ڌgp��Ʃ�~����>�ub�hI��~��O����^���P�B��|���[�9�eѢEǎ6c%�s(�d����o{����?oV�l��}L����������8谰����)������ؾcf���z�	�ZM�4	|,
c�K
r�8�D��'����U��q��z뭍����&�=f���~��8�=¾c`x"0�g�yf�ڵ��ߡA����-w�"W?����PU):�Ȁ�s�:^�׏)).i�h+���LS��
���3ZfϞ=����>���8TX��.�a��i?�9��@ 2��cz�tޅ�nXv�'���.�gD�h(���0Y|k��S٭��'b����g6���Va��A'H}�}崂����,��V�RM7n����7~�YB�c����.9�m
�]0)��r�{9�jq{r)�(A[e�S����G���1����Ma<M��q;]\w�eEec���s�'�
�t���ʣGW9r���n۳gtF02�(f$3��{*��P��=���_��CL�[�n˖-8䠏�<��A�|5�s@_�xB�l}�rf�	*gmT>r$5�}�O=��.��1*Ւ!ψ��oYҋ ��#��ʕ�Ǜ������[y�w�׏Ʃ������ax.��kҸv��Uݾ}��Y���QO1���$
�Akak	�+,(|��W^z�%���ŋ1�b���l�)Nh ���2�qѱT&?m~!��0�6|~��W_}��~���1cx�T�b3X)�O{��VU5
Z�χ]0^z�Ug.=��a�H�[�����!ߡ�-6��n;F_5�0�;{1Ys�~H�];�y��iӦ�?�*�uE�B�'�f�z}���բ�B�<o9zpdm���q�W6lصm�C=TRQ�㐦M%�p��m����}x\Nn!���-[@<�����7~��w�e�͛�f 5�����)<䞮x��:Җ#���c�1�-�}��o��uM�<YNDD������¹�X�k"a�4�h$�|ם�]t�EӧDaaN0h��U���`9Al��4�?��8�JG[�<����{;YO��g2Ac�!�����M�\E�%�Ѕ�R]M-�:�c:�v��� ��oAlP��ݎ[��^p:L� /��o>YU��φ��_QV6 o<�a����q~�7������B�v�iXd�utm�����p�9��a| �Yza�x�5��#k�_��׵k?�ǒ3gNQQ���ŖH@+���۳g�]w�8����wN	�~����0�"Q��h#��cep<L��k�_��?�x�oaa�o!��L=���}��m_|�ϯ�t  ��IDATo���@�Xخ.2���i��:ڎZL�D�d�T���JF���p��~���T�;��
�D4Bn�)S��o:�|��/��҃>8jt݈ʲm�wP-\�0|rǮ�f���lGw����JJ�ϛ�Ϳ�������#��:�F��Av{�m]=� ����}{��z+�_P���w�y���T�X8�V�������i'�ͦ5�����C.T���Lf�S6��z�o�?��[o�����T__����oB�`�'�&,�7�|sǭ�P����p����0�����o�;F�D�`(7/�ҳ<n�پ}�@�>o�1�/K�t�O;m>�{t�X�<�s��	&������_̝?���o�5mF ؽ�������C�� H�p�V��C�E8 �>����}.z�F�l��cvG��	^;Y
+Y�O��4�"�����]'H}<�]8o���>XaLt���g����л���T̙!�tmE��&!'��M�d�H{����P	p&c	2���S><w�D�ݯ�&rJ�X�$���٨5���L"ĸq�;v����Ι3G@��@���er[BIplV2X���3�������|���!	.��K.�$K�j1F=���ibˡvu���L�>��ߟ}��񢶶��w�շ(X�@�0�שsj	�_8���Byaq����^�-[���[n��q���x0S���`R� =����h��EZj���O�|;#\�d	�:�z��(�	f�2ͼ��3*�y�H%��Sd���H��:��+>����o��U ��h�0̾,@�@x'��.{����cx.���`F�7d�T�:e��
��W?��C�*6�	�6Z��&P�X�I$�x�\�`A���/��b�Z�!l7E��/��������c�\�b>t�h�{I0���#]�!�5L\,�^������ce��@�㇜(�(���v��#�<�w�Np:��0Ԍ2�*I_��t���3��B+&���E�g�ޱ}�g�1���nw�mT
ǅ���ʟ Ax	�j���ݦO#�U%�]��������r�ԩS+�W�D�W1ѭ**�ݻw�����-Cc�n vr�;M0�P���s�9m��@�����A�@"8��ݼy3�˩�0�k�m�w�h+�����c@~L�1�9r��A�7��'M���^��.^<S��H�G� lI���I�,�"�a����a%��_h5[ME�(�"W��	,Vdl�I�^����l���Ǟ|�0vdO�öm�F$�C����_L
�s�H"����9}�0���ǫV�s��X���Z)�\��ߏӊ5��	>��`3T�_����'L���|���-@���eX|�
��3�|��|X�j��6��/���P�����1��X��	7�pCum�w` �4[GzN�$�0�<���!���7n����O�c�D������}a�� ��˯�z���3=[�b"\ց��q `�g�uִIW�X�j���1uX�^n)"�)��yڴi�}n9f�<t&�	�d�3s{�?��=b�#���^{m��O���a�^��̙3���\s���ˡ�N�2�]�L?EM3��Z� ta!;������)j��ŋ@���s�$�7��,�	'[�?�:�B����q�@1`�����q䔤�����_�W�d�������h�qj�-���W1��#!"�(�ץT4FJw,�e�D���H0���ݹ�oU����;r����kg̞�u'd���|ۀ���w���1��ȑ��|��� �k�^Of0���I��!eI}&v{��\����7a�<��S�v�������.�,��Q��H�V�&���/�;�V}���Os���0��!S8��`��aM�O�E� �8 Jp
%$"���o��������k�N+o9��>��1���\��-��J(#� |l��i����cy��`�썐31����[͘nJ�P+o��S63���Wd�a�hb+Ԭ�<~�T[�Y�䣻�l�:c��NQ�e�����AQ>?�;��2�R�.S����$�'9��q4�.��-+�o;"�^��;o���)(�H�����w'Sќ\g�@��h�j�A����m:��5���ն��O[����*om>�\[�ݗ+��_����^��cu��D���X��ٳ��t��F�!R��ttv3��P�ñ�ߗO��c���0�5al]8���3O|��'T�PQh�HAA�Eɳc7�^�-;{DK\�����.�*�s/��֖79���[�h�"������B�R}���d�Y��|���`��/���P����B}�b��1�X�d��ST%?e2%֬�z}��VN�W\N�@�����G謉Q�����de���N��|��G �,\hs��f#�����f'8�'�IoܸRsҤIL�А0l
�F�MMpgBC2H3��Ԕ��0:�y.��S��?��OO<��$DYY)u ��V�PX�O5Q9ydD�Dۤ��}����㽷^ټ��ŋO�2����v���cm>o�&Q�*��0=P�?����=u��̜�Ԋ?�0���n��ww�Ŭ���䚒d�y��������&�F� u'y`��;{���#+'�]X�S�Q�lb�ݔ�WA �R����fT�G���x�;��z���7������jvhyv�`%��h�l0:.���=�M�+�>c�;�z��W�{�i-*.�z�rJ��&�nb}�`ggGx*կ�?���o�";0�l��z��zp���y�?�<�xk�q�tUJ�ĩSmoo�l�����s������K�� ��7l!��1)�`]J����������㒥g�����UBÛD����Ըa��.��j�H� Px�i;�i��A�)�g�]0��Q�`8I�j��_~�Q9|8�4������p��ꑣ�y��(`GP���[�o� %TM��[�����3M�=9.v,�u"	�� +>�� Vq�"8��IJV�������c����X2|�{�����u*t.ȧ��'8ρP\������?�����'c��U�d��X\!��CG�Y��ݺ�{0��@X��=��}���o���y��.w�����?�(X̒�*�֬Yݭ��6���}8k�t�Q�����;�������'��1�~�8����1�;,8��#T&t�U?(ȪDȾ`닒(,��?X6��/ٸq3�l�.�Lo(MT�0��r3=!4	�#1��wM�\}���>��8���`7���*΅�Y޳�x���eL4֮`(T��L�6=���a'��Ɛ+�.B����Q4&�� ��>�)��Ɣ�^/Y,oL00_�g��O��?�e�nvF�����h���c�L�E�1�s�.~���}�>\��=,�8F��'q�ah���ϑ'.�lO/a��R_�v�������s�@��x�1j���8}�����~���8���@S���P#����PU4�2y�bT-�b�-�j.5~a�}��G���Q�HE1�LQڦ�@�6�'K�h�%��a��.�)�WU-�n����t�3θ�i0S	"�3,������ظ�Rm,f�a�u�7j�I4n�UJ}���Pa���8:v�Z��L8)���M �p(B��+	��,���ƀ?}��GӧO/�QQ\��Y����a�r�˝;wb��D�{��;v�)����������f���������R�U@|�m22@/�N~�"a�xM�l�ܽ��ۿ�0�Լ�a�JՈ*<���� Or�v<,k�((���&O������7PS"�}P�e���`��w�w8D�q�B���A��)��C�t�IW��KɄ>iHJ)#|`�x�$<
V;u����}���W<5~%ut���Q�=ƃ�d���v�V=z�+�-Z���矇z��7O�8�����fV.��ƨ�m���c�@���_o߾�������"ð)+/�2IfݲHQ¹)~���;�4]tQ��yy{�y�=�Xp�[^5k��wf�~��O���x���!ﯸ�	'�������Sf{<��$��L�G1l���ZEZ�v-��a/l6;(�TP���r;���v����1���=g�J�f�7RRbO0�L�w�;�:��(=̴�;�Wx���Ղ�r�,l]�K���ډ�R, �#���)��`A�}�w�~��ݍ{��nX*�aBQ��jiYyWO��]{��'��U*7&�zU��<g�͎�K*:{�0�hBm>ܲw�~hm%��^o,�+)r{r���#:]`R99�a�J�,Y�?�&�� �o��@ �Nop�qj?��yy,�����T2"!����3�+��EM5�I��C��m0�)C�pg0M����6m:����r���&Z�b���c�ץgR	��?��5aI;J�Z�"��6>gT�dƟs�X����[��4��<Sny�'�B��[�l�����'?�	�kc�@�:�w��m�� ?**.~ᅗ^|�E��[^�Q�pX{������=�}�P���0]`��4��Ԅ�H�RIiAOoG(�%�x��/���?^��G~��X`#��ް��&sL�l�$�����\^6�Z��}��S��u��,�N�ɘ*ǅ�f^�$��DJڷ�����3�b���Ύ���=��UN����:Ү�����k�+"I�#f�pe�0p�K/����/���?:����Z��j���Z$��袆���!V���z�PK��RD;[�ǎk�q�������~h�眳�c�d-j���j��JÒ0�rA,6�egN)�� �J�M�	��F�[f����}���~���n�7���_\������,:�Xط�;Cl%���������} Բ�2%>��cX��c
�0l����z5�W��!�&(�R%��:ڹa.V�wxMun����7@r8��؂��c^_~��&PҸ�4&��@ s9(n1�5�\#ܖ+��1�7��B��}��'�>�/���mj�E��P�/Mtp�'B� 4]�����c� GG�b��m�W<�P]�ĥK�L�����gN$�{�H�~�d���f��-� K@��*ʫh�?�AF^<M$cn�+�cs� M������r��={q*!��@7E�,j(�.ـ�h�"SO#g���OD�&�%�aqJ�O�"��A����q��{�;�X.���Xy�H��s?���B4����==�T�崺�9}0�|�>���nW͙����}���G�,�1e������a���E�`�n��RT���M�QL#O�,Z����y��W^���~v�W����.��/))�vl&~�� �A�!����\z�/��y��{��4l
�(p9���kJF�I5Ս�۶m���J��vm�����Z_QAid@�T-���b!��&�����t͘>��w���/�/_�h�93f=F�d�$g�0 1N�f��#�̱9��Иu�G�6���|����-��֓+����c�(�)���B�<��6wx����k1��hWU�ܳg�B�R��&�џ-�5U��j�x��=	����	���>�n%w�R�u��q'Nć��_���vZ���nܳ��?�r�"��D���P���`΂�LR�4���4�k��A4����A�ܧ g�l1��c_a�����r�-���Z�����z�o�|������-	�[�Z��h�q���b0��,�9$�@��&�j2A0O���x*�6Q�p�M7]{��N� ��	�#'
455�7�Nץ�]���$��X�z�ӊ�w�Ȍ�3��TR˪���Q��R" �$��D	�Ǔy�dC2)@��\s��ų��P�%%RUepY0��^��
��re4@�+-��O����`ٰа?�G��e��.S�]�B;ȧ~/�U�d��JN2����c/ͥXo��<���)�6�]�A��l0�K���n0n���K/��{U*�����H�[EW:n�E�������ϝ�g�%��[�n��I��~z0H�4���jy'�!��X(MHVX��g�\�(�6�ZsRՉ�X��(?/jA��9����9é�T����%Q^/
I���>dVW�[�������{ӧ�1`"��	紤�K
Z%�W?5��?1qT�ܤd�Ef?'����#��9�;��N?yT|��P\9��s�8�%��� H�f�(�f �ã�`ҭ^�+���k�{{�j.:��D��2��^��v�<¨�p� �����.���](>�e����}��Ƽ�H,|���X-<#��@�N�
�_y�|�fT�Y��.������Z�ɥY8�p@�L��0����_̝�ؓ����q�e�]|�������M�7㉹9y��b2���I3"L���Q�}��TWW�q�J��FCT��c%GR�������p Cz����@8eo6{k����u�;b�EW0�衇�G8A�5��8�X[N��Y�ߑh���\-�u���(���,8�8n\Q����#�z�̦O���O�������2��Ι3'�b`�$/,,`iJvW"ΎC�ݣ:C�qƌ&�y�ʕ�\0w�i�����A�CfphId�1(*.=�/NG+��� p�3Cl}����U���T�I�s�B�3��!�-~~@,m�Φ��iw�{����\0ߠ�:4A"L�BnN,�a��:���**��(R���m9���^oh�gO�:����=v���!Sۨ"�d���B�[�n-#r@��={�>y��O_�xe	�	� 揼����7�E�?]T��5�O,&لb�:.n����3����B��2ҳHKДX��Hpظ��UW]%F:C��hhh����o�F�&!q��Ȼ!UC���d,�k3ر��$�2��\�Ǳ ���i�2�(I[w�0q�dds�O��W׬Y��Ob�C|�c`���0���{+_SS���h03�$I{��])"������R�&�?x�l4Q�"SY\���EEP\d�� ycѰ�d��,c���#���_~�����?��{���V��+ItXH�;�LW�E����!or\�qckR�P4�u�����h��}4Xђ�ฤtS	��O?�1m���#�U$b����=�H��^���q;�K��e�Fj�HssG B
눚�ŋ7��I��I��}���x≪��ܼ���m�D�/IiD�����;n�L��JJkF�b �w�����Ծd�\35;�9l�T"��Q�T<FN)��������������x߅.�p�y�T�G��F���h���Y3�\��o���}��WS/:PǓ�9N�W����\�H���Xn��1��h��ֻ�qT�Z�vzuE��5k�m�$b=Yٽc'������6���LD\T��Q	fv���unmN5~��I;����Ău1z��6`�A�`���G�r(
l�j�ȑ�e�M�M���mٲ�[^^�G`F��U2uR�X$�q�U��LDj�D���L���n3�"�.���)���_�fU�v��[o��G,X�����JCCu$�&R���|<����8'j�z�����Ξ����*�@Ϙ�ѣF������GB� (�*��!_�jT�~�ݜ"?��NP2jTU�H�5�Ƣ�`¹HD#��2���!��@:8�vn�x�yg��7��1k.�b���2r��ji�F�n��dLh*��p*4��9�l5ɑ��٧c��}�k��v� ��r	؞�.=qY��Ud�l �%�)��^��Ap)�z��H(�_
G�����7P��;�>}����1c&N���$+��j�:\��M|#*A����90����w����\X\�0�h��Լ9�m.WO{�K/�@y'.�����c$�Ƒ#��	�򣥒E��/�_�G�� ؓ�bq�SF�I4RZBM���z��}�;：�5 �;����	g*�Hk	�.Ȁ=veS�����M#b���NĂ�ti.�l�����C�,�g8E��� :�N D��PO��>�Je�������HF#�#G:��6�5�( ,Q��'��QX��$|�!�C���
U���i�C�y �P���f�f)g@���ׁ���HI���\�Y�d���DZ�����ܻ�Cל��~�S&d&��yX�~"o����u�U1���� e���v���b^OE�2��<}~�,h������%�9rZ �X1�ߓG(e9��q��K"�4�.op�2s�Wfj�����gq�_E�E��6n����?��SN�GJw"�)<���]>���é��P�+�З���އ�Y�	�9� ��؉S*++��;@y��ʭ�	ñ7F=i�H��_s�5�cf�t{��ס���°�!���-[v睷O�8v��mL* `�◄偛�>/?��w����7g��D�8�N�{[\��ʅ��UR2m���c�)�.���ĥ$g���*xЙg.��o���3κ��K�ʇKo�"nȹ��v�yg����]�?��3�T�c��)>��";v,��أ�B ���q���5��yj(@Y�n��@cQQ���N��g�T;��6m��f$�̙3�aα`'*�+\���`�:�Z?���x�3{���k�9������'!������&E��)E��;�D��y��0��/��NgR�GUoܸg��[��z��0��1����%zх����6�u�]R��J���>��G��A3/�-+���䇖<J�:��F6#�|�1c��~���uԇp��P0�����=@���gaǍ�9l{G+���I��\������|��7�n����E�^�	ͫs�0|�8	BS�i$�w"������e�J�W\q�7��r�'M���z�� b�_2~�x�yǎ]XX�h_�}װ��4�U�|߾}x�����D��/׮���O1/h�؛m���a�@
Q��\��#	s��,�O�� �T(�������̞����]�� +�S&�"�� ����əF�ԳI,���{�?[�r�NV���U�D����oK��I�-�@�T5a���%R�4E-�RR�j6�6��� 9�&٠q(�f���! �������%��4gs`M�|�MUȥl�!�<h���Ғ��r]��#dq��mIh@:+$��d�-:���,���u<M?*���@8ye�L�:%2<��1a�/*:X�@	����l>����,��x̐�<)ᖏ�r}Ȭ��h�B��f�"u��2�"��%�r� ��i�Z�������T"���b�.;!���7����,O��&�V����Mh��K0<�P�L)՚d���Mᡊ)�渜`�z�a8N�EJ�:��]N3����s�{o��g?�5�z���Y-���~�I%a��V�Z�f���/�9m��Ѱ��F�Z�4�ȤdRP�w�.�J�wB�Y�n]}Mݨ����ʊ��X"�n۱�o�__5���KGCauxS
��C���������[��c���S�X������������N�6���	c8v�:�8�ӧ���W���O{<�	��d��MUN��ԕUtm�^�.Ь�����Td�4[ML9��lN!v�E2ʰD�8���D44	�l&Wmm�ǫ���+/���[e��%%E�]`�vvt8��*."p�ƽ��y�@(s<7�(���h<�����B}g���ϵg�}��1�߻*��1Z�A��5�v��;�*HG,/׃��#Z��q۲U���`胥�>|8d�.�%�袔#���}�9���4�P�?�*;a,�����a��Gq�qcf8l�X�f�Ȥ�+!�	l��T#��%�	�09c��/�,ϏD��?��0g.�39n��Ç��~#������[¡��]�p:�d��o\����'�k�@OWw�$??����"�m$�%��ٓ��$ɱL�錂-3o��Ʉ*8	~$�8)6Cr�%�6������7�����gW\q����v����?r�0p�44om-�+ٹ�������[SD�~��y����ہ�P=�0�b����C�4�<Dt� ����Kᧄhp�A��S�qX��H>�֏E��b4�T
����ҋk>��nZ�dɰa��9z�l��o����V���g,L*u5�Aꗘ[\T��ц��Ӧ(���]_}�&�P_3���r_�TO�TG7'%5��'���*�)�Zl���P8L�c��w��FS��c�P� ��80w��Y3g�8�ܹ��L0H��������O�����8�E� U�N$����'T%�3�p��ߖ�,�xX\�"�YR������_}�b�)ɐ��F+��'�&g���CU�9�A�m�V�xv$�=�cI.\	,�z�]كdE�c���ə*|����������r�^�����=7^?K,���	���>X�����	�����d�}q���8��n5��t�HO���
��a�w���Ie:Rs��A������"��_�)�~\�C�GHB������Y���S}0����-���V�}�4*eP�4�����B \�QTH:/mq��H7Rγ�$�$ƣ��#Ki�LI+ ����k��n̜9spbq����5@U$�-��U������Λ7��B���v7�VTZ�sXTZJX�8�v=��ׯ�ԗ�+B�v�����Ϗ*#w��E�J��$�h:,�m
�%�e�mk"[M��'8M�I>2
;9�âX�ٳg�����W�^�ZҭB)�m�sɫ���Ɵ�L�5��DbT�At���!�ZD�s�(*S,-�|(JN6T�]X����7���'I鱔0��z�P��<8�?BQ���\���-�����n�uq�m�6xPA5��C���[�n�޾N'�v�b5pO�bq,*++ىB�R��N��\���Tu���r�
oB��r�cM���;＼�
��%-�&�7v������<�������	���s���z:S��(������Z��x��/�ے�������ːu��1D��wҤI�w���˗_��K��bR� ��~�#a�8�^* QQ�_��I� 	X�dk��TQ#��j�,HKz5�?�5Q]�y��T8K�-f�!B�zn3Vc	X�{�w�ʕ���oˆ�(�����$2���88tj�����C~������b�9m^���n���xa	����1|P;�Uc�K& �z�<����b�-Z4~��� ��pN 7�!l�Q��b�L_c^^Q�Ћ��20��'�2����>�F׉%��5����k§.����H� �GcIK����mR�6���j��Db��- �-��#7�Hv����as��y����e��ƣ�1�EIf�p����X.��r���S�.>Nlkk�f� `c�o�.LUϖʖ�|�T��"�#��SҠ&S[4NN���a��Trjᐈ70��Y��c���.t�ɃE�C3>���'K}��^)S�I�U� ��XU ��~�����)%=�F���J�`t`	���RzA`S
�^"�C��-qKvH%9�Q��MF���I�i��x��0�,�O%�3�B�$��i��K
�x���[��j�{��	-�!Q!�H�����2��D�v)N#OEr,�,..Y��ٻw�o���|���a�%��m-�])�	z�YVMm==�H($�����S��Z���OZ���]���啔EÔ9!-�ڻD���-bC� �����x,�i��,�d���q�l>_զ�7e�|����$5��8H#$.����2�[� �RF���ʱx$D�϶�������᥅_��I�p{�I�r����n0��a�F؂��&f @e��Ja��o,VRXU����@P8��$�R�H����f�?���p�rc#?��yy����ɓ!fV�X5���޼y�U�.���$�m3&�Ol:t�@s,�[���݇�����{6����Yŧx�$on>�g���d�I1>��D�P�vP�b$�^��-'�'�E��k�Z�F�1��
Ǟ}��q��n�M�=������p֙�����/�����`��YƎ���M��]��8����j���Ś"Z�G8�0@�*�>���&�^�F����a�H�D4Q����{��9+�}�ݷ^y������ͷ�%�ِ�q�ڵ�h7�����1�ڏ����b���OP%F����=U�;���$�;J>?�,ȯ���O�4جf������� �`ISb���p��#܄��)��jr��[�^w�53f̸��_�؜v;5�*f�Z�����BJQǅ1cj]nwSS#�dDi��m��T�����a���)x������35]�Y�T����D<:@H�P�.GqGW��l�U�J��q�ɤ��@QY�#G@�UU�8� �������eW.�:erk[+q�T��0��&M�ka'�� 1�N��id�����|�I�2qT�y�-�S^�?R����'c ��RZ�LG���&烈O�qJJi[���@�2<Ɔ��=Jn=���I�|>Eg$6lӦ��I�V�X��Im��5O^�x"[R�Y`C�o<܇R����	��l���Il���(.�k��j� ��9��E��x�����z.[�8��	����[_:ѫ/e��t1�da��")�b+�ây���v֙I��zS�Ufa��@8P��~}�:[����Ҝ��tϡ�	�\���M��K�����L%U���i����t2���I��O&�B� �i�f�O��0V�)�YI����S����ӦS���}��m*]���Y���opRbJG����Z�����7���|���M&��v��l�]�%e�~^ޒ����*�MҠ6�^�h)�يs�6W��>E�B^,x�[�vױ���[�1C�p/(I[x�D�I���Ll���E.jo?u���ٔ�9s渱c�}�YL�����Ё�)Gt��N9ĺU���*>���
�'��X:<�Z�|9ưs�Nn����௿�zyy9��={�pW\Ix89���E�+�i�&��3#Nb��֭۵k{��c�,KG�_�����6|��lR��/��}*٧d��6��f\_ '<w�ԩx4%ʈ�!�<�bvpڴi� !���644|�6ȍ�qO�Lq�X$ʮ/��TR?8J�F�J��A�?�7�F�]��>->����<��Z�K/�4q�Ħ�&9�`�ǎ.m��3�<s�7_�u�]5�UӧO 4Fn��0"uA��N�|f���ʋ�ʴ�cGL!�I���OZ�h|�������)���x�p�6n��t���n�ml����Jn��H����.Z����?��O�^{-c:刋��&!�B�G<��/���@�G��@$	��	?s6$6"�w�v��Ѡ�o�������8'L�0�t��uk1����n0��{)��B�+)��n�6�O��"�/��׿-��Q�(X8�c��yH�45(�T G^,cR�Ah�KJ��l����@(���2`��ӡ&�m�u(�ı�N�#�����A����9,	f�'�h�"�i��.�$��tB_;=�9��.�q2d�����3�{)ԕݞe)8�:�g����b�6b�\��e�̼0	�K�C$S<9��ܳ�H�B�b�k�������:.���P�2H�|b��$�ag,{t4�9��'!WON:C����J����d�P%�DcW�`�� I��d��C��&�$��B*C���(�'�@Л��tS��T��b(��`(����/ם���z�mm�����I�.�d�Sn�$��ɩmA(
"��_UUu�����n�?~��1U۶m�D�0n&����p��_a��!�Mv���\�W2 #�'d���.BA�;|����t)��7FC���%c����t`ƑX��c�>C���vڅ��I��W���5R��y��Ezh�)��TK���FMNJ�ZU4J�ı
��f��44������a�SR,,��،�͹�M�q��V��=�!�7�����j��-G����P�� 2��ۢ������#��,� >�Ł���M�1㣏>��ك?)"1���N���X����T�%7���q2W~�bwȖ-[X��p ������n�sӦ����N�`��8�'$F�T1�LT�'�� .�;���X����U�G[�qI���a��WD6lX)t�d<�P_�cǎ���.8�n3�6��
&#ԐM�n���7(�σ=%���~���q
f$�<y0���������B2|��P�;���0���睷߸�'?kڿ��)��]S���ۯ^Ⱋ�P(0������#+N�h��D���q�͂c��譊�O�ANb�,&�dP*�#����f���;*.h'�w�����7>��s5��M�Mn�"�����FB�1�5R2��_܈QM�4Km6
�r1o�:~��x4r�pW��zrT�U�t�5��b�P�����cR�P�-
V��F��"uSS��3�ei���\�:��_�︸0�ɩ�0V�dE�g��C���>fK�ٜ�aq΂���ߖ�Zh {$N�iP�Qr�Yp�$��%�L�����c��.���>���vS͏�طo�o��6��aFL�������l3W��f���{�������d3o���-��'���fU���t����״T�WN^.Y�r$�0q�'�r�i*�֙T�}�C��8y/��������u�<N��s�8����`��|+FG��=�s^���Me��9�����L2 ��]Xi�%^붔���Vv�H�]na�j��@=g��0E�����Pɍ"Yg���=(��R�jcp��é���v�Z�]I�^�8�x�d��F	�V���|���hf6����H#ı�=�:[�J������m��B����IN��mڷ����t[�F��x^$���\|N��#���U�����^F6p_L�+�@!X��HW|Ȣ⎰%��}�ݏ<�pmm�~H�xN.�E�И����1MΓǐ�XhQx�O�0�	�g�Z��fϞ���j3>��� �\�d	����/����`�x�ǟC�̚�����b��]��'W�p�̑��$ǨQ�8g�AȀd�z���z�1_��q��Y]�%�'��&o6E(�FUx˨�p�h0S�L�ɑ�����(�<(hCo��-��L�^�ك$V�wLf-ӓ��O�1N���*��eGw���L����nia�?�;�(&�
(j��.�ӌ-((�N3]�X�X�2�}^<;�YMV1GY����n�W�EL��&�}�`L�-����P�<Xؐ��kk�m�����J>STZ�棏@����з8���K(j#,+)��W"<rW'�� �h�3x��<S���=l[��S&��9��}>v��۵*����h���g�q��LU�أ�v���V��j�O�dKY&~6��R@�bH���=��V��yW7IC�|Ӽ[NACgf��l&#��t��z��~�Q��GC��Tn!��ظ�u��ч���h0�'�$L�<��3���x�<-8�;vl�a�;�|�0qj9�{o�}��'wE�$Ǜ�I�(����9C�`�(r\}����9Y��� e��A���8-�f�Vg`�FW�����+�>��+#S0�[MN�c��R�(u�Ç���>"�z��d'�}��d3�����K�l�/9MHL?����a�󥑒}>����Y�V��RdSnn>��E=��dB�Z�}��yT��f��$�-@�����5�e����-F£�%��H1K�B�jB5�F�6b	'$:fh���1r���?��,F���	�3������pė��e��SD�n���V7�m�)����j�R+����s�"��+T�洚R���%XZ��K� ��B�R�[	�S��a���������+RϠJC
�%a�d�sb�"R\J��T%�8��d��p�x��!�H���*���޾�d*�P>фzBn9p������A�a�F���B��HP��D�6"	>�E WZ�:������x4a��)n��R幜���Z4)�cI�A��bj�@��qY;�D�pT�H���8[BI�>0H���U�`Đ��(��ltaOONe������Z8~�o����?l�k���x��:�MĉH��q�m��6oQS�p� �����h����w��0��#-ԝ9���O�ʡ��/p�W��nٸi��2�d����H)J��d�U�O�7�وn=�����{`���ڛ��4���e��Dn��al�����rs�S�L��>�hɧ��ɂTdM�w�Q�$�����2��}-�����/>��&��DP2X]��N�B(*.0{ܰp����E��1�5�ɄM�?x�3��py��'��`���H,s�Y�xMAcL�f�mDr���ҩ"��ќJٻ�T����oHܽ�XGQnQ"���v�KN�[þ��a_�=7������	�@����)�T�����y$5��ٞ(R���EX@�IE!F�%#��d �����m�B�!9�`���AUn(���h4��t�����NQ�S�۝�,T�a�5�������Z�����,h;����a�GB	�X3f�&�	5�Hy�VuÖ�����������Pm�^S�`4�rQ���N-ࡌr�)KtJ���;��N��3+�H���AER����h�������3Ϩ=j��%twp��E��ZMf�� aC�x'&����P�V0ۢ�MX���u�]�w�UʒF;�O�g�g۠lI��F΄�Zƒ��G��3@��,
����?-]�t��)���u�V�^%Ȩ�{��Q�bP�t��!�8��Y~+�p
'�jZ�I�n�������~��գ ��x�"��:�Jd�Y}��>G:�3G�ػ���r���p-�8��Ij��{,�c픤Cn7��[*"&��
s�'
[Vq��x٥L�=�'�J����S�+%��,Ty҅2�k���k���y$��[�"���У�4"Q��]xk1�{���!�h���f�mR4="�#�a5��D�ozg�pGD�HeJ?x_��VΪ��O/�W@��"={��6]�
�OL�-x>zj�����x�E`�I��� nhh�i.am���ރ	��C���׭[w��2�5X�ѣG����
���}��qt�>qmڴ���z#{������j|w˖-�]1cZ�ѣ�QQQA@V��,x�����1S�N]�r��c����F�WɆ��q677/8m����?���袥���Q7��T�M�<�PIi�#Sz"DS3��KNq�{O%�,�Î	R=�`P�h�͎_&A2���eleۅ�<�mݤ����Ԓ8gjz�b�N�I͗�;����*&�us:�,��Mt""q��� ߡ��L${����@M��6XU(I'����YW:IKTO�����!3�}� -v�����#��iB{3Z9�@8?���s�G�*//�H?�����n��R�-~�1{I�S��5l+׀p��s�%R�M���D�D3W��3��,�����.��:[>�Y�ħ�^����R__�l�a��{0s�d���<8.}�_�S���ٳ��2pt��j=v��~��5��dx�ќ�cG��ޞ4�
���]�^S��f_����}�R��#�|u��'�~}�4=Y�Y:�Ĵ�l
��c,�O��#sK=��.48q}T��M�P��ZO}��)��Ք���FC�Ϋ���Ky٘FY��,�+^�2�U�T�jI>aMDr��������?~�a�F#q�-K����F�Š���O�)I����b(��ă�(&E([��(%rt*g�y)B,2�$�����D��6�nM�s�t�e�ĨM�go4Q"��)��+i��u&s|f�����l5f�LF��6�4Y�1Y�V���Q*���q�N!�^'��Z�Eq_���86O�bT�d�G�yhbp9I��xzgg��}���!��L�RP��G�狼���mɒ%��]�F���(�� ��K�8�F�����b8mm�'M��~�z������ر�q�5��f���fΜYSS�6�����kܑR��陼L��_}�Us󑺺:W�kͧ���/Z5�n�Pɜ��ߗ�!a۱cۡC�ӴiS��z����f*N�g{�فG��AuMW��!EE�LY��'H%�#�5������%%%Pe(?.��o�X�;j*��K}�83��H�d���'e��W4�vTҐ�
:}+ݽM�u��2��	z�U@t��V�|��y�5I�z����-0&��	:�\l���j����bq����N���Ir��Ǐ8w�K&6T�,�YQDL���x��A�K��I�!<��T��$ ���r������9�_�ny��q%�8�eM�:��b�̜9�+P�P(T��w�ǣz>xZ�g�s��IS�����qg�{e�K�������1���7M{�|��T*�_B���NT-�L���-3dQ"�-��E�}�n�>�/�f͚���	�D`v3�2��,�9��08`IHY�RF�g�W=�5�@�Xc:+T�
�\�+�=�lM3����V9y�x�KT�`C���:U�)�W����l�/��y��?�݃�6wJ�+�����堾�b&�!
h��	�I��	*�(r,_���7L�cC>uE��:,o�)�2�@����!��޵�~�� �6������Lc=����R�Y�����.Z�R���9�}4��,���5(�S�����e�.rƀ���ǞL&]�+�t���N��ӹ�P_�&Сix'��*���	�0��򃽔���K't�� kB�ьguuuA<���Ecǎ�0ae���x����o��++�G����T�6�nux�q㊆Q���`�����������$���c�t�RH�ǃ�5jTSSS[[��I���s�a;*@�"_�T3f���O���X���1���b��h�����͛ÑԒ�g�����t�� ��ΩSI���Q�D%KJ$m������L�qidIVpx$5͗'�_c���Rt�ȑ6�lV6`��Ț�A`��|�%ѭ#���_��=%�)��)D�����A�l+'и��L���=F�wb���<,Z��|���Dʛ]M'�@a��0�E� �F�\�����I1�>!�C]��%��8"�Nץx�l��<��%��lTH"�5P�@\�|���c.(�=v�g4���^�/6�A��H�f��QZ�C�$Y��Xa��Yd3U}��n�z��.v�W[_ӆ�reg�)��9�:g9Y���mJ��C>�yCCJTfP�f���v�-�^�bNy�^��,�?�ĩ�3������r�pV��0�p���L�8Yg�C�>��xS�]�2ym���K�7�cFp�ʞ�����T�7��R��¶�)�6)#�$�ч����=�N	��z �>LyȨ�S�����4�Ϫb�Ec1	E�=l�u]%��)�N�a�2e+����!g����I�|Z'�b�t��xRD�"`s��l,e623�F�v,K%LZ\%�A�p-e{�O��O*9���I�h7�3�$?�j�iX������s2��D�_��i6'�F�H4��Q��?��8���1/%N�	��Z�:%�nIU��'��u���P0�Ld�|�.��c��ޒ��u���N�1<0m��i��#�e*}X�L "u�0}n,KrKJ9� �$�c"��v�`_k�(�c��j��LĊ�
#���;g͚��}�������+/_r�0�|������%�~MVG��o۱LVx�]s��ٸa�����:jTd��@�����#G�5�4������ĥ��S)Ý��u0S��+��@7z��?~��ۑU#9�-�DBx�t�Ǐ{�p�� Y�3[�/e�nWY��v����ܖ^HbH�@�H*H�2�2##�>*�|3(`��GAF��DfF�OS@B	IHo���O?�}���������|��'�{�>�^�zW_�eA�g2	��BL^,��۱�����/���k9�b����@uK7��y��R�Y�hpy�F i��3�n|$@�p%_z�%86NCVY�J��a�{��	�jT�ACPM��<~�:҈�5��4�B������Hh
������;'�/Ĭ��:�[f���&��At�m��
�Iry����p��Z��e���t�NP����~��u�p;���ǋ�p	e��Z�"ވ�y�KO�F|ӦM�T
��S�,���Ό���5���_��a(�y`��D����^�x¥�Ƥ(��ʥ�,�eH���2`>$<(�����v�M�|��v}]��H9�=����}/夅nh�c�ݵ�jTVB��X5M)]�E
��}����1���9s�m;(OLM�ɤ4��̫����`H�׵�����K���I40��Sn縷��{~��GZ�C�o��D-<�0�R�����P���-��ZtS��Y��*��,VEt��v��7�a�E�Q�A�7ږ��JM�{�FՒ$��@�<У��k�-d.�L���霻e����ď޵4RJ���G!�|~B�5�M��h���-#er�A�^*ThڍXipT�M��wI&^�s��APY���+�� ���8-� �t,wv`���ǅFt��K������XN`d��3�0��Hj���$���+8�2gv�޽�V�Z�bŻ�rj�9�}��g�}�W�h�qgS`9^~�啫V�q�Ōm޼���n��f�.��rxj�l�,�W8�	���9��s��q35~���ӟ~��^0�-dj*� ��`��dʒ_/�>{�ҥK���)���/�O�Y2�&Q����S1�cV0�H]A�C#Tؾ���
q�'�F�W��¸�
)>�t�ޣ�GP��i�#(D���Y~ذ����4��Ü��4D7��2!A�5�Ĕ�St����h�|�9�1�7a@��9՗�[�w]�͸�&�ʡs)rT�E[��'W�qĹW_����菍��E6M�$D���[�����#
�;��5o��/��[���2!S�.|�e�ݭ�E|H|�Ŗ`������a��W���M�W\/Q"N�n��ay�:�Q�u���8���G�I��e���i����Z�C��^����r���[�D&�4b�S��8��ʟ}zdb����o��bWf̘O��s�6�lX�ܨ28<���o𼊴��G�yϋ��E�ⶄ:Bh?(�	���e;OQ�ꮣ$��Yu>��_-F)�)?!֢�j��Jjp�8Я�p�u��u�ݻ�R	�
��܊�9O��K��W��M�ӫV.�T*V�_4�Ϳ�1�ς���:���]r����,�e*n� ��4ʅ<x�b�:)b�slA��4��i�4	�\��tѩ�AG�Lċ�J�� ���y�Ly�� �%���E�q�qK˦�|>-�p$�l.xq��y���]�(����;�H�R"��28tԥa��ܕa���� �6,�\�Wub"7>>�/h>}k��a�dƅ�n�ϱ�K�&������e��g�u>�)���OK�k�eA��1�ō
,�R��>˖�	���瞅Ά
��
9��7�?OY�����G���~�o׮]7n����Ӑ F�|����۷o���P�������v�Z�>4k֬u�����_�YgRɖm����D����켅xք��HIčj%�J2N��/B�����h�o7N���yۮ��1_#����?����Қ����]�<::H5��Q*�/�%�
���&�s8B��a1s����*����x`�$���ĎQ����H�������֢r�J�-N�yIʤ���s��X��}����L��h}�fE|}�,*��e�[�#��9�}=�ކ?F�R����8y��Gw]�8���8��1V,�H;��%h��������}l��jD1:0�\n/�D�=q!|�������ZlPzXg���쪐KЄd���c�#��#�����7�\�|9�ݺi�X�8eb�vww�u0��ݻUS4�N��!�;��`�����H��GX��^`T�2�D�:������t<�����K�>~�������MNWuS>6�"ʚ�Y��0s��������L���	�
�>D���-d��RA��fH(Or�*!?$I/�܁�הS�v̇����o_;�ҍ���E��]U������)8t���3g�P��� �����qwT]y���^[��E-L�KF�\,G�N��U�p��X��&���+������3��R���O�C�ʝH`Z_|*����#hn�,�&R�aDǜ~�S^�|8�S�k\Y��$���bhr���������2�"�!!GÔ�5�zP-ŁS[q�:�S�����{���! ��!ߛ^�\?I�N�}K7A�.�a7���M�lg�@��8q�����=p� �]�p.K��\m�o� C��r�-�^z�����[ϚE�%����S$���'�<���O:�$��W@�۷�����\�5P 	�J���&drj_<<��X`%<�������`��E����
cc4*Ի袋�͛�Db}=�45Υ�ҷD=���(�i"\j���ɪK�&wC������9�/�� �9��D�`�֠��RU-�`Pg]%��z�g��U�V�}���cbƈ����+_�0F��k����  �`#�o�><|���s�L��B�S�.MVm�])�r]�wy�c�P��	�J��N8Z�~�����T�~ǆP��w��T.�ҔR�/<L���rX�4�f [�ۿs����jI�Z�����s�FB F�� �7(IR�:c�Pʣ���wR"C(
k5�j5�+��
a-��R���5��1m�
V�A<���{<�鬠B�S^�?K��D� sE?#~��dѦE�MiQ���eI�@�Z����6:<\��K�G*���V�8q��y_�sG{K_�FFl*�'�9(����9���ݳd�T<�O�6��P�#�(�
����4>;��p�QE5|E��r����8��a>w�566q�\ Rٓ3_��;��ԃ�@O$��Ӈ'��Zm��.i� �,�[$+�V+�"�Q QY/��UB�1 � �?!�!�qZ��4�llE�:�P�PI�-D��,/D,м ?M.�K��D(P��'qD1I�e|�ɸ�hl47:21�%˯���䎕l�oRy}�m�Kָ�����*�|Q���UbpA���˕�]݄J[��p,㈋#|N�W������Ƭ�In�ܵDh�Ը������Pt� ��,%�NS�W�����Bpӈ�D��iIuEXS�@.7����Z�d��iZ��S�I<DskN����폍��b�B����I�)�$��[
�LA�3���ahh �c�Rhj��E(��r�6,��V*zr\[F������������x���G����/���]�����P�ǎ������?��^_������|.*a�0��_(P�2�Qp3�*8/P�R�g�Ai=�	�R<��}}=�ͭ\1����p]�� ��v5_ß�3;.��{���e��&��B1'��e�Q�%�"�m�I
ϐ4%xf�AJ�i�v(�$�!I��=s���`�k�%�c�N:ڇ�)Ĕ�>Z��{��Lȡ��L�'�a֟#�)���^Pbht+I�ep�����h`��*gs����Y�,��jWN�iii�:��cl.#��@�@��~�:��ݡ*�ʂ�qGFFp��R٠�	�c[�����Z=�GJ}"�A�'n4=l'�$�|������
����K�l@"��z�!�$mO&�x{L�q�O찆�:2�� Z�%n�.\8�
LL�KV!���g��كE���6n�(v �3�BY:��JP��e�`������VɆL���d���K��.���(�i�M<�&OH�O�/A�7��}��;�b���3��W��k�Y�9�F�&�VN�W_}5$�֭۰J��C�t���:_y��������pt�J��ݳA�������>�ƲU
G��6/�x��=d!b���P����bH���7?<����E^t3y�՟-�����i��(A|nE	�����Aꉙ"Z|�O?�S���ėUE���~�+��G2�/���\-Z?��]��p�aJpZ𯘒����Z�ͥR;??>&廔�*:
�l,>�&WQI�C�-�7���b*���eU����� �'�O�g�uB"�;�oI%����$�f�����'�<I!��'�ɭ)K�rɆ��H���U�d*12��[��T�PD�2�[�ڲ�|�T��]�-Ӎ�����C�$uA	���ˆ��,�"��]GKb�
c,\�~�O<������/h�T/a�o��O9o��]y����{!���ى�L�����]
W������QK)����5-S������/j,=�p���eZ9N͙6ԑ2�=-a9�x`�3C��617�cq���VV��`�N9�F$o�P�Q�R�6���D%�J!���f=W]3� ʯ�zJ�u�g�ջ���6<�iӛU7X����<�홱�ˬ��pd�ޏC��f�0�KղX�d+�����yX_O)�jQ Ci�DކO�[$ddX����8��g����EB��x�K��Qˌ���ޢ���#x 0��h{a�Y>,19��v}�O�kY��X~Zʌ �p�`����~Zߟ���æ��K��T�8� �9�F��������qpp0?��*gv�w���9�7�lѫ���k�V��:?�����F���Z[)j3sc�[�CQ�r���5wYICU� ��R�^��E����lD���i( 6>�3����|\X��{�<���6ʂQrG��FX2�3�2B�Ti��P��qY*��ʼ����V�tù�Q���"^��{\Рs�Γ(-B��5��O[#�U)QT`t��¸)C~���B�	YSOV<ny>ɩ����/9������.��3���V�ZP�%RT�q�҃��S|>W�ۿ�w�y��Ehrg�L߂'D��&u�ڌK�������x�u��`C�p�1�(��;�h~<lAh}-?��@��wg��Jb���R�� ��� �\tu͔�{�>H��Gѓ�3y����zͰ�?��ijjH�HĘ�,,�O�@�Aa_������=ۮ@��E�[r����ͤ��j����/�75�ؽ��w}n�M7�z���Dz���/�=.8����b����R���۱���J���
�)U�"��8m��Yv��q�<��p(�{��p��_���J�K_�bkk3+9���ĕ�
&K�؆Y*&�S�����C� a�D�Ǭ�L��q��2gnFթ�a|X�x��i��h1� $-���2�"jP�`N�Q�x�*���Rxʱ%��gK�(��`��ےd$N���5)=����5�Hw@ �G�r1=�����e�}�P�q��q_K'*��-%�D�d�E����1e��4��pi�'���/:%F2�Tqe-R�L@��'��9�(��=�	�
T��o���B�v��#�X,��l��:��pd`k��Ν���c-10�E��F0L\0���36*oEM�����ȜR=b�D�[Ty��������G`Z������)?	ek�����<��_��w��ͺhn�ʚ*M��jÝ�?:/4��wy�T�D��U��}��������l�u=�xh�U��h}�srGP֖6�Z�q�]�0���^}��r�0/`S�Mu�z6NY��y��Ҧ>7M�[TZ���)�F��t]�4��H(�����$���v�D#�ka�C��-���b��\�,��4���pmR@�b>/���p�)FO(�R"ԏ�V|}Y6��F�o�@�EYB:Dry�%�n͇�`��]�'��k�F2fq>����ɽ��y^'�����bynY\4�̠.q?�YŲ$����Ҟ�A#,\�v�qa��\@9�9��7 a�)G��$s`8rW�����A�m���+Q�{n4W*I�ɾ�8�6i�1�TP�!��g�x|d�R\V$=��^,����c������+!�׭[���Ss2����������O�P<����!%�lii�A#�8�Đ�������)A��^��k�����s4�uǎm0Ò��t.-b�*Q;E�*-�0j5ՓxRO�Zծ��Ӓ������t�O���"(�[������ŹR�f�:X?�N�}t����n"y(Z����É\���Ǵ�������R�ĩp�O��t�d�U)>��J�����Rq��wO	:�9p����/!��Y^ǲ%�k�&b��C��38�w�(Z0*�`�\�0���	W���,F"~����˖m۲j����\���-?������]�a��GHQ�8�X�D����(˩�f�b�.���ݑ�(qS�x����/��pM4����W��`0��N�����ij�f�g��@�b��v��XnG[H��s$#���=,_��b�!����F쐌6r�n{�:�`'+q�x�!#@R�Ұ�āQ+W��R+!�ZF��a�Ď�",����*��4k���b��#�?j�]���G�?J�(�D��ڦ�Y�U�Gw��k��+b9q�"�^�;�5+A��"�@����dM�^'�T�a�.���h~�f��*Tsͳɤ����Pk��IR��09��[
Dt���w
{�հ;�Pk��'���Fݠ�x��H&0yS�n�i�KC��x�>���t`yaA��6���3�Lg�q���7XVR�OT���RE�,�ʪc���J�O�X�:b!a�C�\w�wuu��M��;L���oղZ~$�����ȘT��n�Z$�*s���@gP��A�*��C�������h 5����=�g%MnJ���OMzI���h;�ۃ�Ų���o����,_��ۛtG;z�_�cg�}�F«�s�κ��;��\�H�L2�/�9<�����9+w'���3�H&3�ܖ���NtԖ%j���C��\�aÆK���e;%+��j�I(lԅV���2��0w���R,���r�ڍ�3R��*^I�PZ�"^��4Kuj8��r�a��ZF$��o0����}G����b�|aB��b��zcS������4j�]���\���Ď჌��B郿1n6s��q� X�M!L��	��e��J���qdԤ��rE�^����.S	@>�a��vz�u-�i�}tZ�ٓ���/P��nq�g_ۺ�m��	�ׇy�4��`���A��&S~T� b�^X�,ݼ��+��$:�E
��NS����fm���D�q)��ŋ����{j��~Md��D�k}׭��G�}������t���ٳǴ|P��9s�9"e��/XU����Ç��]�vÆ�=zv��o�:�3#���l�+��cs���(������T�rZdl���P_�
�i����M3�t��ԏ���+��I �A�S��5qr���hqy�h�Is�W^?ŝ<�ᴈ��##�/P��S6��)S�\�y�l��~%@����Ie��3u^-y)�U�8N�p�~lj�F#d�8�J��~@Ii0eЭ��F��l`"P!:�����Vi�!ч���ʛ��s��E}�����C�J&=�ե��XB�,;|)8 ��r'<溺,�Cg����aբ�M��bI-i�/g@�TC��*v�����Z?�NA:G���,��4$�U.a��76H��x�8��7�|�E]�Zr���ǿ��~��eAV8[��СC�ׯ���={v}�UR�	:��sݺu6�H�R
�M_��� >s�yg}�S�:��^���j�c6�:�@����W�ɞ�!�t	ϓ�G{���콰�H����,�f�t_�X�N�-X͍+�P�ܰY���@�Ї���TZ_x��'���j�]��1��gf3]�&9�����>w@�A�1J�B����.�n�LX��n/N> SpDJ(5쇩U���V4PČ���!�ZZ	��\���/p���<Y K�.�5k�[oq��BB���կ��*�N?��Bc�v =b�oV��Eā(��drz7��J�D_�: �9s�������>�O�Oy%\�c���]K�mӂh*Yo�>!c1�'F��	� �����r����F&Ee�p/Z0oά�ёC������'�R��h�K��"I�����~�W�Y�TFLqs�EP-I�1Rc�MwrHLsR�����v]�?�t�o6�I�������<mrG���a��tNRZ?�g�]�Aw2R�N}PRU�Xp���r*$$(eF\b��*��2��X�O�<Ʞt� j��ܦ^;Z�d<�e�i;eQ��Jg�''u�EE���8x�0���]�:	>�.�}i��He�Ɇ3i�ΎV���/���.�u�N�Y��IcIr�6��gI�Wc���ER#�:,��_��t�s�t�D���B��E�$�C�S}ĩIn�2���Q	YF�3���"qb4ת>k��J#�4��	����H )��F�V��8RJ����}�!� ��@�T�W��;���^�fێ�_��ח�__{ݺ3 [�ׄ����b�
��y���r�m۶c.jm�{��a.� ��;w�ē'�xBcC������:*�T OdT\�3>�������KJ��M���x(A-D��U���3��4���I$�-��c�YJ�H6G�G��2s#�-��u�q��X0@L9V�T��l�ЍT�^�P�C@�>~���d��#�m��̎�r#��]B�.��x��F3��xX���L]I�
_�Σ"
�6�#c�jjj���=Ww�S)��R�Z��e]OM��hJFݐy`��D��1+ZX�%c_b1K�y`p���Dѥ�t��C}�r��7�|�Y��W^yeF[עE��ipZ��N;R�W��h����J��r��î�t�h}a3q8U!����$8E,�G��Rt���������6�;���UZ_nF컠�BE3��78�;�N�R*!�1�3�؞�F��d�^d C	S�e�J�HZ<4tDҽ؆�BI������J)Ŭ�6�*��-��$���j��"(��2$րh5A�f4G�v��D�����yt��[&����'�ūF��q9C���F����p �:	�J�&[��y��)�>�cP�$T�HWA���E���ˊ��H�b�S�K|o��

�Ʉ/��D^��I˓d"�x��cj6��A��n���b�I��E����x�FL&###��E�����C�2��}�T֤21����Q8�z�9���0J4RI�� <D���@(۟�>s���&cк��g{v�X���~�s��M��#�66d՜:�mk�����(��!ޚd�@�:�)�N]��Ҕ���.�0)� ���x�ȑ#�0�C�Ν?��;�|��_�q��]v�g>��|�y޼y��z�c�=��SO�����e˖�n��g?�J�g�v�hOC5 @hHA��芽�,����5kN����G�I����:e#��'��hܕ)�"��!ְ��T��yh����A)�
iv|k�Wţ?sZ�Z�j��LB�.��FH$��)f����B��HP�Հ	����F�4�]8�Qe��34j�`����q+�J�CM���BayqJm��\����ʠ>R_��O��$��q�2��F��l�gL�Ø@Y�"ǎs
>����U�9#�+ŧ�0��ݱq����5�[J�e���/*>�~���Q�T��	��+��K�R���|Є6?�r��o;E��v�`�H�YAE�������T���2Y���صo��4Z��B�3���x��ht�g;e�kw�ٷ��,����lKW[CsC��Y�{;EmF]'	��r�4�Ǚ�l&}��RI�����w��*c��R���M!���l���slld������p衁�#�bn"�d�[���DhR�:266�Lɟ���D*=:>!���4�C��+����� ���\k�&�T"IU:9�H��W̗&;bZ]��2�65��3��8���ic��V8XL�}�JlS��j�D*}e+?0���)��� x,n'��h9�$�i���xEBL�:�j�S�u�W݁��9s�POv��W��F�Xe���I76B��T�_v�j܊����e�5 ��G'*���hTv��ÉOŴL&U����q��G�w���<f�K��>U��*�Y
��7-_@�,{N]]���^�mj7U��.��.%}Ǝ��hii��8�����7e/��&��DbLq�uxH��T�'��C`���LxTp@�bM��]�`����HiIR�2d;��CX�t|:g���J�25�zՊ�IיI�X,AvQ��l���E�ݝ4����ΩھU������x1me�����.'����I�:����<L���cT9ۜi�\\©�
����8���3����ٵ���nȃ*���#����N���s��ϕ�fW�@��yG�hz�R���i8}̴�jx��q�e��SO����w�s�-��Y������:u��֖�|����;�n��7�/��z�D�400���������-y���5��w����%D�{6m����tmVgG�R���5k�>�����az���d��Ͽ��k�����yv9Mm��s۰]�P�	�m5����Q��"�W��N����@��?A]̗l�|#��t5ќb��S�������H	�_�����U3��W�u��\,���������q�-�#����Pp>9�~�AQ�s�43�<h����R�M��x�jx݉�,�x<�J%2�G5����@��°�h���Ēq����
5�9���&3�#�M]������\ F��S��H�N5_�����'J���Y�t�es8��r�skh�	���٦��(f
�B�KZ�LK�D�gˆAw��lc6���ϔJŮ�������f3�.��s[{SCc��[𼩥�q�}���ŗ���x �D��qk4���d<{#^��I��u(4�N%��,��Nm1\x��ZRmstd�Ue�����ēС�}
��w'2��;� �)��|��з`�o�s��8E����s]���{��s�����"�]iT-4\��=�����0�,Z ����~�b�
h���Pv�a�� �bŊr�9p��C�ߝ=�{�֭�2��@u���e�����`�>3WTw��2 �"��~����XE"���a�����8�41A��Ǝ�\�v��:�ڒgmoo�M�c2UL��f�L��1XcR�M��S��(��<D�Ys<|�}���J�c|A��>ʶ�]p?�����G I�͝;���ƹb?��ă�GY�rG��VC��g��ü)��K=�]�tT�Gʌ5�&iQ
�Y	RW�Bu:�Q\�P�P�+�R ��3�n��Z
�#�S�6/�Ґ��X7�^Ө�_���a�B�T�����ɯK���|a�G������K�	U������T�T��Nʅ4�w��ʆ���(�w�Z�ӱѠ
Z�Nf�v���c�p��$�c���q�$r(?�5��}K�j4㉫��jɒ%_���>�]#g�[�=�|��;＃�p x��g2�i9��s�ʵkq͉q�O���o����h���N�d �p�>��Ԍ׏>�Sv�UW\|��=��EXy�yWõ�F��f��=�������z4?h���	&��8�5��{8\⪊�/h�qO����"��l����mC���Z�*�U��C*��Щ� �_
jqB.`P]�'�C"خW�p� �*K�؃VC�4E�7U�h+�P�/8�eQy�&~���c!����� ��s��eϞ=��ҥK��]�v-^�D����Y{�$� �K�9J�!x�A��'�{J�ha��ǅb8�jIX�S�:��a��z@M�ƽ��$�-)�q�� ťkP�i}������7n�½�⋷�z��� �	�����ۇ#�ߖ���j�:�3��E*]�l������Z~�42t�����ܞ�WN�R�:L{�JDe�S%+&[���2ñ�#�{K'�H��٘�ܱs'�zH%Y��4a��a`S���X� ���44�	��N-�LX����׎\�!?�(��Ã	
�%%z�� e,X E�ˏ�|0-����x�޽{��0E�y��T��f&#ޗ��&k�)*_1���`��P 0x�ȑ#����������W��2YxK� ����poS�����ki�[�jE
��V� ���bH�m�-�� �3c��ӧ	��0�M$0��bN�,c�(����lrtt�1Cx�2�*z�p��G�;f<Y����\g{�m)�3������K9�RQ\!L>�9��J�m=R%�	`XN�|B��B���x24:"Wo<�+Wu����an��iҨ��(RyQ��͉qB��A�5�Z��ϙ5'x?���c�|�U�I��t�>a�\�a�qt"�34<:6>�sv�>�L��p
�Ѫ\��Nрډ�*�D��+�3-�NvuwOL�`g���42��? qL�<�sD�y1��x�A�@���p��<y�*��|�?�z�O/� ��Ƒ�=���k֬���/�
9vFf������/��Zx�y��.�I3����c3��0�a�o���|9aET!��ŉ���E���y睫V�{B曅r����/����LG`.k��g��U"B�M��"ߊ퍰��3}Pr�T*MW�i�bPYt�R���踌�d��O�>I��"h���-�q��`�还%�-|�+�b!G64A6x�]q�R6� ߔ4*ڈQ|���'��W�j���U�#F	Y�U�&#��Se+�iS�H�e�&_����V,��gK���b �ٞjLL���B��(�KzN�1��V9�Jk@��c17b����AE6v�칶A��'B�;F߱�b�3R�9�2� ! �	c�g�yf��w�cx%���yЧhW\��H ��\Z;�k'�S-��Q�%4:<���Uݘx\*;,v��ۀ<#lo3��E�D�w��
S�ʣ�M�����s3,��9�c��d�1U���y9S~I��a�8;w��ܱcN��AȘ,Ղ���~�V��c(�Qi�-B�ٍ��03�V�%�3���_���ׄև��D�]y�BGUf(ֽ��`ٳ�>����=|&h5ȗ\�� �|f)m
)B]^���ܞ������d.y0d]]v��� >�jժN8A]�l	��8��ݲe���F ^��ǆ���r����"!
��K�`J�AΛ7��:ȅ� =)ȟNa+�:XG���5�8	0\/^�.E�%T�ٌ��wdU�<����ga�|��7��S-�J���xB׫�A��zZ����~K<P�	��)ڐGa�H����Z�����Iw� ڄ��
�:Z8�Idw�T׍)`�{�2�+��i��+�d"I�]��DWe�]GA�u3	V�B�\�M&M����ImÖ��AO��,w%���T-[��$c��W!�Ě�g�>�P�A�/�!�VK��a!y<�Z���!4�'Cy���A��y��LyR]a����C��L+����m۶D"%��ַ�~��w��駟~���?��O�y�1��k���k��)x饗�yz���O���MP(l>��%&r/�ڵ'��_{�6\�5Cp�g��x(�j��TQ�DQߪP),Ü*���G��A3��a?�6�����S��Q[��\�A{��ٙ�c|j$����!
֗:5�j����
�_����0���Tj\�C�)G�6d�Ei��׬@J���;�8N>J�����SZ _ 7�%�(h��Җ��ůu>k�J�!.�*����#EU:�~�.%�7j!��;�do��Ɨ�'�Źs�pc&�}qM��(�X�#�̱r�� ^�vc�Fp�.n����QY'�$X��RK,8ڦ+�����i�"%$�>+*�s��!���h^3X�pI�6����zꓟ��%KT�H�<0F��)�� ���2L���Y��,#*ղ1e�� 6����(e1|����ͤ	��nd�02�O������v�Z-�ܑ`���Z'�ttՅ^8gΜg�}v���8흳�J�Gd����B�r-iSo����t��a�W�0�U(��nr��r�衳�:�+�hiiR?��V_�������w�]w�������%����.ȣ\F[��E�X���U�Mt��%�=���_�g����%H���m���h�Z��'����̆&�4�b�`:���;�u�V�Tgw�ѣG)zVWOI�jE���KM�|�� ��N`^��.��D�Ę�H��.�S��N�-V�B�X*V@�x*�J�I�U.T�9:�cV6[��S�|�p��gL�K{���E��������>M.�u�M�c�}{���s̈́G���X�]��`��~<��P��[*Ud���xN���r�[)���1�)l_� ��I��A"�����)�#�;�f��y뢅�GFr��=>��E�k;"t�6=�I(�t��["�ŷfk�򯷟J�qv��Q��*t���I���ے��J��$���00�_M,�X�.� ��IS���mohh*Wu�W>W��lǅ�mk���MZ[�/_�c��T"�i�&j�����_����<��/�rl�0�����q���\�fM�p��^}<����ݣ��V����S�A����Ȳ�.��RȁJ���;�Ak�
�*�-���P�E�/��7r�#T0��U'�ҥ^��Y��R���]�J��ģ���<��4J��o�@��"�6U]�!�ڰ�-A�dTB@?�պ�|�,i�M��I��8�V���3�ܘ���ӤѼ.�Lep��E�9�jӔ��e�S	�ji($GP���̘�.S1t�rop�2�2��5�&i�q�>��T�[�������ir��CT��ё	�2+����ʌ�阡�$<�Q�/�?�	���ql�9<#@,ķ*Œ'�����,ݠ[�j��`bӰ�0������%qa��޽;�O;�aq:�;���EUe�l*�wɷJC#~F���KQ^���"f��64��坪����Iq�<�1�\���!�.@�@U�?T�G�|��K%h7)c|�R>M`��\���^���ףӪ�ӿ�>��={.��bx����s�P�^8��?)o��o�t�W%\�$���/�����&�<�'����n��k5-���reN�H`���q�V�X���g��я~�M2=���3�Ra�G41&��@b��-��vÄ���C-[�ޑ�F�s�����7�����z�~���կ~�۔`�������fL��H��������<�lT�A��F	�7�޻o�Ӈ>�!s�L媼��1���{-ݫw�q����'�x���$�/��0/d
�	�%���5�:_�hQ�)ȧj��)��z���Rqx�
��Z��/_~�M7��Ay��Bss�#�c}�p�3�<�cg{��;e
���K��t���3)IxG�u��T�K�21k��2@�������^�r��g+i����'6���9.����0��p� u#�}�w-Z��$gAn7g.9�Ja[-D5�󔗲�eؚ���Q"m`�e����~�a%jDO�o�0��ZCϱ���J�_� �5�U���8�0�'r#0)fvup^`BƁ���g�
��P���Ep���\�
�N�ڬf� W����<���\���W_�X�z��%�#��P�3�����u�uׁ��:z�
Z[�	�K@T�B��t�q/��P���NN�i��7���"2�e/޿�v¨<a��"c�'"
`X��g(�s$�*��)���i�τ;�� �,��<�"&dCЙey� ;x/N}����X���D�r�%�'����p�l%v�iq����<*l��9�@y�	�bԤ�;�K���:>�����}T%^Et�R�0(�R�C1�0T`� 0v�]��aV����ڽ�x_-M4btt�j,*A���Ȉ�����5���7�����(N���m� !gl��3J7`�&�$��E�O:�R>����Q��C���dK!hj�Cl��8X+���ጳ$蒂8���O0n��Q�+�v��đK�u�H&�Ԩ���6�L�J���wa�q�&+�
�2L���w��n8��^��g�U�	Q� �2y�������.��(�o���"�
,���
�ja�j�Fk翹W�Z��w������T�+r��Q,��o��֛7�đ)um|<��Tw����8�O^w�G?����o��)�:Iե����2K�J3I��u�҃,�/�<�b��
�|��`r,Qg��q�
$m�)a�it��B��Qʧ@��fX	�y�嗯_�����G�x2fɈ����r��>A�Й�~����*!+R;fRb�Bm�ձ�e�I�b	8��g�\��ZV�y���_��s<�����Y���	����P�_��=�~��o���f��]!W�VJ��Nh=<�z�EAY~JFB���6X�S�M�Pa�gOf��LX�V"<I4RPqx|<_(�v��O^w���|��t:����:B��{�m���c�r��-�%'��-�kK��jK眈t�.5nP���x����	`K�`<h6�[�L27:���	��@W�v!�K�7��->���gK�1\DM�]��wن�}��_����Ι	R<|��呒��țIBk����b�OW׬�G����M�Az̙M�s�ly��\�-��y�f�aPf�X�����r!sg��m/�����3W\s͚U+�/>�̾ݻ5�}�s)���Ty���x�����n�V�ζ-x�ua�S��0\��&OD���p�Y�ߋT�����J����;Q�( ���`�
6�T��(��kٺ��S�H*>=�ey+�h��	��`0yF�������t�f�	J��X���>�1
�8���t6O��(����T�NH�'$���Ut�I$�f+��u��R���Q��`T�ٜ�e?�u�Ay�򧖞I}��\�o�㎫���P�����O�$[�s���C[8>5L��>��v��~X֙�^��}^%B�o�D�E���n��|�`jVCC��8�Z�
�۶7�S�ђ�aq.?a)���c=�b��K�0�~1�HA �>��3i�|}H�R0}ш�����8��h����ybs�5V/g�G%�K,O�^eciJ��~Cc#��
�ԃ�����W �X^����*hP�YFf���=HC=[���Y�X��!��$׭ѧR[��b�4K.I��}��}Ǟy���x�-PKu�M�X\�QBVT�-S���~`�o���֏~�g�}��۾};~T�)����Ԣ��t_s�^X�-���{zz�6�c�=�+J=��acɘp	 ̞=�U0�8ハ<��7��t�}�A�Ϟ=����l�{�qQ�S�8(��A�m���>bw��"�9s��޻��$F#��!w�2_�'��5�� 8��u�<���>��{����E��w�Ԡ����5i��A�C(���´��O� h�X0�W8�eKO��|����{q�x�=�}d�0:2N�<Z���?ƺS���G���9���~�w���������Bʒp5����t1h����q��Q*V�B�1�e��4.{�4g|��a*U��۾��{ҩ��Sݖ�K�m
�i]&��C]q�>��D�f~w�Կ��4�
[��&{���i��f�r�����c�u���q`Lamsg��!|2'�c��e�L����5sl��/��O�/�q�2�9 N����?^y�P˖-�kܣO���K':�L�C�N��`���u[X��-#����o.����.����#��۶m��O�x����'�|�� �lp���z�`�BH�9}%NQph}i^�2���c�dc=u�dRIuL|. ����Վ�T���.�IZ?��Z��r�
tI������rx���3��T�i7�p�}S� W��9R|� �<��3�
��*(�0�$\�!=���{�ڂ�K2Ȏ�o	F���g�Hb�aP���D(ՍD=}up��'ꇽ���nM!��*�U��m�vE	47 7�T�֊M�,L�����R�q A wCU���8"�
7>i��uʎ�N싻��N�/[��h�ʁ8 ն��UAͿi��p�eT�s�� ��W�b�����0	�䎢�Z*���~6i,X���N�C{R�&�ɋ��8�<���M�{<��]���A;�_i���� "ִ�~�����s�}�k_{�פȢ��!�2�U�[�$a���$�l�=Xu��X1?^�	ʦX�NJ�����!��'������zG�L���H>b�-���a�ץK�B���Xˏ���w�<�$2"#�2-W8�Qĥm�&(��x.�
#	�S��J_O�v�k��f��L��S����ͷI@"P�س;v�V�Z�����/~�u�3h(8e�,�%TD0�W�M�^�8�]�
CUd̆ˀH��t�xZ6�Χ>u����
�O�X�@�>�I�.�8����������ϯ�55���;6\|�=�����/cU�3Z%J��FޘC֘�aH"H��an�}}���	�)NLPQ�fe|��h���=؋�k�^t�Ew��FT�G�x��Q�O�/�8�#OX������s���}�y?��6���sF{s._!f3MNČ'q�gM�	����x���&�us���k�,aO�P�Y,��!��Y,Q&��b��;w�馛>��ۗ,]�.�������l��� ���z�����5\��=��/�h������5�E��@�t��"m�U�������~�D=@vd���Ι��o�<2E�T&�{��>�E,���ŵ�o��+�����o��[e�s��X���ݻo�������|�7��iӦ' W�Qb���f(��Ne��g�|�j�R53�9�RC&^��=r0�����v��=;vnM�c�X_�(�IB�T�Խ��ڀw�[�/��G�_}=Ga��Fο������k��8`�12I�a�勸�5W_��_�b�=���2K�����&r��'&���s��������eFC��8o� ľa0u�U8c����І�����]�N�X2)�i`/�[[v�����o}�on�s�I�G�&bq�.��p�[�n���B�484Z*W�z]6ˁ������Z������6K �����T����"N�Dc0)�F�,@2�=r�
��%�]ݸ��˖����{�4�W�9�������F�q��1~؝�j�b�r�tի��W��'���+�vIj
�OZ^aqI�\���	I���1�c��u=�S�v�J�ķ��t}��m��9+A�������̙����R(���.8VO�h�Us�i��f���ўc�\��s։'�R_�����v���$3���k�>�>eL�=}�T���r�RO� �Y�(�;���(A�}ز^�Zb�,��Vb��t1r~a޼0����xA��.�X%���W�K6��Y<)8n7��ke��qbv)���U��͛��s�=���O������8N�����y�4�0�;��w���&����syx?��3�8�o��g��P�;E#���z�����J���2{���n�p�u0#z�!������K( �o	���kӐ�q��uA�3�}�P8��/�����;�y���F���C�:���ۺu+��u�]{�~�[߂wE�0]���3x�iN���	Y�8R�.hHT6L�m�-��k�y��s��ܬ��j% #�E�X��(ܠ��Πxԯ�/���ˋ����/��7���W�����L)�!va���|hp@IҰ�6�L*�Sq�'b������}�]w����?������x>/��u�r6(H�$���+���Z��?��#��������l˖-�2�F=r�7g�l,��T:�q����eb&y#^-�.�vѨ�iF�Js�E�b��ܷ��O�a7n\�d�f�(�i���揎�F�0R=��]{k��SN9������:�����'�e�a�����0R�I�L��1Z O�����Fp_4����+�dCu�;�'މGh�q�&dSp ?��,�5͠�5>6!�L�,'�bKw � ��̙�����������8p�������g�C(b���ynǠ�
!��fj�1�ƭ���/�#uݐ��SvJ)+ظhSG���$��x��>���eҴڗ^z	7��k����L�ol������8��
8��=��W� .�#����a�gR���l��n	���@���	Z2���K6�y�1+v���>�Hg�i�83�֬]��o���~�����{��mi&'�>��ti�F�k]��dRp�!_P,Cf��}n�We=a���o�288��Dx.x	���V�+d`.G^�����l���7l����O�{�2w#c5��t��s�~c��=N�rB�9JO��� �@�Ba�N_Q���D��R75Q��X���c���+,)��I�HSRW{������7��_|���&IK�*ē�:|wN7�P����+�4YE�`��,�%��+�0��5@)�p��9�����
G�!���	�lW1�e G(/����������#�;F3)�n���I�W�����H��4��8�hA���I9T0r��!8| %<���;�xft͚Ř*�_��M��e��r��q�d�`;KT��{�ݻ���w �^�������Їcq�'#[z�\���_�z!����-d�Fgg���(lj�2� ���G}�g����$ܝ�����Ng�0�������y�8ϸk���w���� KG��:����^�)G=]����FΙ3�����aK��Ս�-��&|�BA v$��q�nV�_(nY�<t��j(6(Hξ����.��+�-[2i)�Q���b�	�I4<̀�c�񸕫S7 �����S?��O���G��@��c� m�%h��M��EERb������)���ҸF}]K&�8Rr6��~������hn�B���QzL

3�.��O�Q+6�G6.�~��h._���я_��.y�����'?ٻ�ܹ���C��A����>����D�5G(�~}��L@N��.��^�T�1U.�U��}L���_�f�m��z�g64��!⹜�x�.�a75�	E��1�8)U�7�~K�]�������>�?����1<:1o�l��
T]��.!1��*"<�o�,�s��NL�K'�njkm�fR&2a�z���'Oj��d"�i��ο[~�4AN#0^�����K�|rvi.v��c��A�aS}��W���W^�s"�lh�y��Q��u<Q�:+ S���O����r9��4���38ȡ9��R�Y�N.�/���l��`���ly��`�{����n�[e�A;.:aɮ]�zz�!��l��75S���-�=��s�9��o���_�
�A[[Y�U��)Ѫ�](���4QU�����[d� �)�?�KQ}hSS[-�],�чv)֭;�ӟ���E������N�'y��|�;w�����O\u�y|���������rE�8v��1�8�=C���m]=G�K�cO��^Cc]6K���[qJ,�T�I3x�ܟb�F�N&��� ¨)�͋{Z�Z���K��9�ҥ���&��g�}����%�R�m�˦�7n|벏b��ſ���>���ޢ{F��m�(WJp7�9�4�Kd�;^���g,��F�ZTA�[Zz�����~<�>r�W�=�;�`&&Jo��ֹg�����TߺeK+�V\���:�������?r��?�~�{�֭�T�Xt`���я����m�r�l&�r��K�?0<�c���C\+�z�l�J!�zJ��J�>Rv�X�	��G*�4-�Z�Hc�X�BV51S�i|��T+�S/(�\\�2�T�1m�}*�n�W�i�Z_ls�礤�t9yDW����3۷o�<��F��!���ǿ=��O>�o߾SO=�s��i`]�Ng�-t-��� ��;;�2 	��E^�Dˈj1	���������Ң�M�����hi��-Ll(o����?��O��_�u����#�����h�R')<�s�=�H�ur���wv��&���=T��� �͍��T�)q!�~k۶���O_��O<�?���𧻺��,@�pվX��M�Ha��e\�N��;�/_n�A�,��Q<���δ�cx���b����-Z1�$a��w�4`�o���.�e?uxh �/���n����<���R����
�g��Oջ}�7�p�����|��n�G��H`C�թ�#��X�N�#K�'ӛ�o���v����ڄ5�S��:o�������sg56��p�����ћ%�ÃpV� �vCK1|����Ǥ������_��UW]e�j���a�ᠭ��R����C�H�G����a�'x��]�U�,���~�m��XЀ�E�q�4ʙM��*Mj����%Z(=E����k�qc��C�B]t�_��;l�E$W��]���w7͒�%����$ qfAjX�����'����~u��o��?�ӎ�o/\��N�JzG)��rě+�}Cn����̥�0Enb�z{{�D�4��றk:��뮻n�yB���ܾ������?ɇ)O����Y;욫��T���{Ϟ=�fvQ�c�B���
Z nR�Zi}7�K�"��~�~;�[�wvv�vO�!�����R��Ù`������.mp�9s�;:�u��֭{������ohH�DRR��"ϙ$.B��j�w����ҖT���0�d��HA	E�l�י�p!vK��-m�+W�\��#]3g�+ڸ �&e�zؾ�e˖�垲z�)�W��G�y���k���[��"��i���7ds��<����M ��%r0�Fi/�s���$s������l�{��]��$��}T����H4;��o�^��?�뿾������{�b��9�!,cP~����	�Ϯ��0X��N2�+�ѪYCxG���*l"�N�HC����o)��R�Q
'���{�В�!�)\�g��V	BKŒ�����1�.������2����s�QLR �!ʸE3�����kl
����A�̀��ؼy3N���w�����S(���Z�f��Q<vt���8v�v<�*ƶl�>[r�) �G/����Kc�r�vә ���q!C&���j��+�;��-_���s��ϸ�֛�=��{�?��?�nyw��sv�X	��ȱ� �?�R�=��K/�������勃�M�1�}��5�\r6�}ER��c�g���{	;�����n��oV�Z�u>����#'��8Wf8SZ*�O���R��u�p��/}邏�.%���Z�L0�xC����'8mR+�2��*|B���=Sr"�2>�3��[������~���?��w��AL���|p��Pq�o�&�rt�e�ҵ<���n�޽簭��G��;�5�%���P~���M�y��?��Bt�#]!#:_����MEi�^�0z�G��<a_W���g��5k�Ͻ������ڹcS#�8��=T�&���jT�v!ON3�J[kg�P��7�y��h���W]���|��EBe$;z{i6.،}� ���|��R�`��Ƀ��5�`O.>y�=��;e��w��=;����?>x�0,�
TU��А��U(���{�Ǌcc�b�s�ļ�KiY:$)Di��#T-�G�sE�2�X��lpoG��X�X�ᢶ
�e\4���	�.��1p�(�kh���>��x��S��'��+�jYI�R-ʙ�HC��;zp,#'��QH?��Gȸ��Ϥ	�(�]���֯_�9x��u��8�b��[%�R�q�X<����J'i��ǁMom��6��oo�������?���]m�M�%(6a�حV��GPf� Zn��y�S`����x����
�z�m�}��k�R>;:������In�I�����_��W�8�.����~���o������--1C?p�h2���L���Ii*�D�T�}ۡ����3�kG%�T�'13;��߰}���Lz�9�?{�!66>�e�f|xּ��b])7��z�܆�Y��.�zƟ_~m�	�?y�-�\�����߶s\�D2եǒ1#6��C�9I�xO���RT�z�cO�[2��`5wQb���
����k��
<���H$�k��A�tC=�k��C�Ěi�o��z�kB�Z+�/�_}c�O]��;� ���_��?���xa�������Y`v��Lg���Jax� ju8G�AU�*!�g�A��5�u��T��T��b�j\d�e���z��>wX�e���l��Ș����� h��L�[$*���R����jW�6����ң��M!}̲⚊����@`�k��d��ֆ�a3
w��8<Էtٲ[?�i����ׄ��� HO e�+����Q����|�͟����uuAK�@�L]tŒ�5�Q}M{�����9k�d,�� ��s�=_|��?�
�d����#���le�.����_���?~��v�j�|C��D���+�!�R͠�S#m�)��Y��$�=�pjV�:yժ^}������^b�2S�q�$L*㤠�qh����[n֤�/��"��҆��K+~�Z_i�dĔ��ǽ{�B����:'�x�@/��
������>��0P͟G�{^�B����fww7�V����7�p�7���n��?v����������᱉s i�C"�9u�FE���q�J�6�����{�IU�m�gz����FY`i6�.v�%�`��XcO^�k�FMTb�&��j���bz슊�E@�R��l���>����9K������p�9s�s����]ZV|޹�s����wך5-�>"o��[zR�7��|/��by��

������y�^�~l��*��R��p$���~1�.�4+ģ��%[���$��BD�w"�Rq���������׿���5�dB�P�"���$��a�R�Nd+�a��7	Yj���������:k��	�����Lݯ��� e�	��뵵Jľ߯�xRO/ƌw�w��n=��c�=�ag� VE$�؈�� ���PA�CW.ơ���s�g����^Pӫ�U�RP��hH0|0\���SV` �w���qP[�H[k3$ѩ��M����?����������O���Ǝ��V�yZ���(�u��&]N���zյ�����V�� �_��MT���`ɏZFm�|�����>�o~��n��8��x
�5J���=KK��::ۉ� {6)+��bM ��_$\�L�{il���R��<蠉��ře�6nlI�;D�%wM�0t��G½��ч����t\*95Lh�ѽ�����O>�d0�7y���$��V��h�/�q	N�� ��%g�寙^d�B�1�&8ЧX�����7�P+ֈtp �⣏Y'����8��EM�#F�|��g����Ν�hѢ=��J?#�i&-C�QMgˁBzdi�!qH�QC�@�O�����~()�u�Q��	���^
AY�,�7|�h0~j��L=�$#o�9����i�O甂Dǰ˰��l__�:�ؚ1p��V���"P$r
�����|y��H?+EJ!���t��ګ�\�=��?nl��/��f�2��K�s_l����cN��+j���	ݍ+�uy�~�(0��)E�535��Hح�З��!#�ey%�g̘14a>�Y>��3�?�8�b�JJToq����i�z⫼9�u,��ώ��##��I8�����ܰգ���޶L� �6�9�pec�6m����Ё����?ӟ@'A^?��CPF��Z��5�"��h�'���7�q��_|���ٱ��ޞ>LVi���[�[����8�l�j�#L��r�~NfqF1t�8���ĥ�����`4�~�7�t饗~�{���j�T�I�4Fu8�9	����޴a3�Ɯo��y�Տ��+@E"1Pފ�a��֎�b�;�P�h?��T�vZ�P-�!��haq��{�,I�*<8���̿v�ѣG��_�s�Q��z뫯���H2�Z��M�%^BJfUWK�V��n���\{��Θ�6�6m��,�X�J��$X[��O,�vy�&?H�V�Y�[�lQ�&ȷB�`���[Z����YG���?����_~��IQa탡t0b��}6����a�D#��vnS�hl0�������!�h��l�`l&��#�ǟ�_ =��]�@UMC�Ij>�<[}
ᔔt{4I$�x�Һ��k�����O�����?��������<Lo7��l�k{�<.�� �YX�`��v���ц$��.^�� I���s�IS}�1��Tz��R5���Z OM�H��n��ի�O�<aΜsfwz�`�<p���:��t�%���25l�F����8j¹���z\rɥ#G�¯�-- �?�G��T�W*����R���`���*C.�WD5�B"����#�㮓N<�'?�ɟ�"q�5�*�[��?�����V���/4��xL �,~GZ���5S�H�w"mw:��pA�7Jh�ŕW_3a�<hV��+V`��U׌\���hA���5��Fb����Op�Nom�(K*�ъ�`3�g��<�+�geu1�Cw���q�c*~	;w�}*�8�X$<Ck��\�p��V�l�X7��-��/�nu�����yzk�{<��PRV���E[���O�(f�[�v5��`�o�{��YR\r�ɧ�zҩw���/~�^��gl��D2%!�!_�AqIWwO&��&u?-�#NJ9F�!��"�G�8$
;�j&I�:-���V#���*��[�T�;�����=d�f:S�akͭr}�����2��c'��[�>u�D^�x&vf��ش�Y.%g2��RA�����;����������'���;4k���H��9����N�w�܊'�����:~,G��J��q�Pb2����0^��K�.��s�B�������4�~;�F��UW]9�)h���e�X$�$-0�&�2���D3R������$&�ˢ��� FL��W_�f;��9R(���r4T��D����>���{@�'O���{5x�Q���̚��k�(���eh�(~��c�@;�;=*�x(�2�"1�'��˗/�g�}y����_��_.]&KȖ�U�;[�FБG�;z�� �+��*�/b��z�եPH��D�k�H��P뻫���1=��0c��\8��A����؄ݸǔ=���~��;������.7���w3��v�},j��.����T��z���e���/��,O'��`@(z���4Ø�]P$�F8����K�doO@��0��7A2.��E�s��?���^�0�@Y0�$���&����_���#k�?���<x�5�Y�	�P?f,�:���{%�`Hi�����v��SUU�|n�#���b�5������~��'���y��;o��7�<�͉ �x���H�mYI��*��~��p�	c�d�Vtvu2|}K�SXi"�U�thhaQ	���
�:��;:�w��z���5-x�ʕ+�8���x���=;��>�B��c� vp�[�ֶf`��j�BO��}@�d���v����-���L�cG� $���%	���t�ܜ��i)�.A	��w��{>���>��/o����6���;��
�-��׏���=�]v1M�K'���)�oo��-�����N>�0�A{V�X.�M������h�r�.RV*�N�̴nޫ��H�Q�)p���f�M7�~�}��ʏ���+V�(�*D�>�TR�Y�?/[)�T8aE�J+�.zHmG"oB�U��}'v���o'Nt8%Cd�u��؈�)�+=��6b�u����1� �cj�EڬǸ1�	���w�;�;��0ޅ�M�=��%3{��Q��6��v.6��RZ��o|�PG-6DS>��C5��0Ǫ�PKM��a�i��!;�>pp#H���x�aٱ!�����x=�n�;�_���y۶��.���s�ќ�	u)��,(,�:M�M[:�v��.,(m�Z��W����{�׌�m�.'_,���|,���{X,��P�&���a>���>�ʯ��Y�f=��C ��| J�QFȇe;i���j5���������&�j;%v7e2C���Ziiqyy).X�p!��7�x�%C�����r�X�]tя�c�//3hd�U�_Y�V�ڲ94·cQ�l����ֲ.8�HY`GG��D")�w�%���B��nKժ]}�l%�u̸�W�|�7�=s��w/���᷹C)[GW����˧o�1c�%U<�J�0�H4��!EHkՐ��o�ܜ�:W]�x~MU�r���*hnm9r�@(��d����߼a���8R���%�t\�Ҥ���A80���m����?x��>Z�<}�d�;c"� �>wE��/��[מu�Yn��,�F$B@1-�S4)(�-�1P��̫��@�*��$��n�*/MF�ʋÑ���ah�2��:--!A�u{1\��Ր�o�󑣏}��c�y�B0��O��E�@<nl+e<}�	�]p�^��c�
g�D�V�#���>H?&b��"i���0��MDc�e� ƌ�=��N0)X#G��H[m])�����+�[ZV|���z�<��wކ�k��I���d�GR	WJ�J��B�h4&�o��X����j��
S����6�v	N����A�0�6K�r(�R�|Pb-��&jLVR�tt��c�`^ZZ�`�?�^Htx�[��.�p4�=����M%y� �ۑ�?_v�a����cIl�����W^w�m�f�Z���u���}]X"�1t��MB�b�A�gH��n|h�����d���@�?����e�$�TU]����s�^s�PA���
O�ן�0��$��@Z�]c��6�pR�>�;�.�8��?<�_��%zC���{/�U���=L��I�ш�HG�����,�<�����^�����;����z����^k8��������~�m\P[틹�{��7S��Y`���>�xb{��j*���R����?�,A���kkj�є"$t{�d�e
qSꩺ�]m�y^o<�Q�w�����p��z�
���'M���}�W�f��p	D:顴$�ؒ.���u� (�z˄J��.�>���TeE��Lwv�p ]�H�X����W^2��?@#?]WF<��%��,V{L�rW�������ӆp�Ғ"�fA�U����y-�T4<��wJ��$Î6��t#�_��T�g�ús4���(��������+`�Q[�e��QG�CԤ̓�H�_�j���p��bP�h��B�9LuK�ٚ��Ӡ�|�T�$�2S2�ƌ��/9y��g�y��Qp���m�Ŗf^�`�+�Y �V��F��(})�n�[x� f$�Ov��c�]�P!�)��5t;��KA�D�2���3�<��c��Χ�zj������S�<��s��>.w(Ir����4g���Х"��I�$$�@�6�K��>��
`�fH\k�62���hY-.�pb4��_X�����[O<�Ļ�d,�mQ26nlk�����}�I'����Z7����	��
��}��D(�.X��@�.q�E���&bB]-��.�����ߟ�������
���ڇ-f�|	G���T/4�ӎ�ʔ�vN:;{�ϰa����E��b���$�Ut�v8#n{&�5~�@\!��0��1n�8�px���^{�';���_{�%�\XX��
�h-���"��g�}��G2N7$�H�~I��)���FxS��I;}�tp/�3v� '�ܨ�+ܪ�IX�hF�6	��b�[[[��s�=���N{p��X�eb����^��i�lIb�P��ǟ|��ٳ��nڴ��9�ġc&uA4�1!�ngy4�-���g:��!`y]b�Ç�իǏ_^Qq��Wϙ3�3΀���F��LcZ;b��Ј��sc���s�&��t�a� ��V�����bln��h�^lI&��a"%ӂhw1�|�æ<>�h!	��&��|��9s&4���7�<�*�r�-c�3&O�M664
}0��:�]ml��.��n�C���Ƴ?AfA���b1������	�2��dN��a�`�'L��"ǃ>x�=��1�3M��w��&b�M!ӊi���P��1A�?�a^7n��6�J���e 0'Z F��M�ÇO�20	�;�)���}y�uk�Ac[��ڵ�H�e��e�m2��[d�+�RK��C�(' e��R��şobh��!��ϫ�x�@�\��7C��/�0�6��sc[R`���]��#ɒ%K�n��o�q���Rl*Cdbd�O0���/!������u���E��~bb�S ��X��Xac~����4�FL.�@:���K�b��qǏf̘	�
��������ڸ�.�34��9Xˀ��M����dUz(�Lv2�8$d�nP�Z~�ζ[#<��D�`(�tɇ���7�>����e���������=��7\�}	�1�1ԓz�gQ�/��� RxJCCC_P`���r�4�2:��~B~B[E#��g�(M>d�DW4"�Z�[����g�={�>�<�����j����	�l� rv̡{��<�l��M�}���L�0�L !
�(zE��a�0w����XC�!W=���eh�jX��bﭬ���HK������q=��_��ȦІ<��N��t�Z�H���oϚ5ˮ����٭6p�;̯U!(L_���	�W(UXf��Ek�A�1���IVZ��&Y@��e޼y`��������[��/��W���@�����ɒ$ÞHY[[���A���J�{�Cv�1��-*�W�Xq���
�)���x���v"z%�1����`�y�c�m��Px����^	`��/���/�zhŊ�.�k2�����,G���/(���vt��� �K<���AX��)4�0�v���6)?�b�X���Σ��CQa>��@�pK,	4ָ.�~���Ǎ���K�<K���y���x��v-3]P\�ΣVF�ᥰ����v'�pX~�XI��UTMj�p�%#�!��,EƥXLV�����=�
�ܐN��_���
lm���D��XD]SIb��9REr(�]�@K��
������qn���LH�E��!�e��O(*hwA�/Cg�I+/���Z�%[mh[J��뛤C)���)2�k�֌Oy|��r=��9F6���F���G*��<_��M���Og��̞��D�k���L\h�\R������֟�j}ICٳ�/�����b�<�0�\�(�\>��H~S����f5��@����p����g����N���{�}�qǙE�q��
�R0.���2k@����.I~3fds�>�QqR�%����"+`�aKh���)Y�D�z*h(�^ܣf +Cj�ϟ�8y�q�����x������L�Sj�d�)�4|����L\�t��O����ڵ��Bs�}/�ab�ݸ�Z8C)m
���&ae:2=)xֺ�W��V�4\w��?l{��G76�a�@j��јؖ��$��WH�¹c��&��c�]0�Tq�W��h�1:C�A��ޗ(o�X-��7�%�]��w�����x�'�&�VM
?��ÿ��ﺝ���	���LՊ�{��0h�}!� �b��`�(, �WI�P4�jP���]hNlJ�&-X�4l@�7p:z�A�מPU���`�2�F'�E�	�8��'[%�O�Г�1ATM1�ɮ�2L��PV�Ӊ%GFK� x�O�=,{� %���\x��e�ĉ߹�SN9���'�\�r:ޓ�
fO$Bq���q�'�|�	���B��ŋ��I��<���ڻ����/�A����#R�c�R�䄯���a��COpR-7�x��>����Jc��.��!�����~��+/��86cZ�pwӞ�h����?餓=�PC-=XE4z�J�cd� n%��$ڠ�{A\Tj̏h	>���zl���$� ~�k������{/�NH�,�4��j�jc�HNM>fS�5��/����7�d���8�'J��e���~?�%c�4�vDz���'��YP�bf�-��_.�0	{.�' ��Tj(
ܐc+�7��H��i��Q���{����r�!w���/�&a���~��2�f�i�!u�um ��*g�*..R� }��bD��=I��� �V(,=p,&M�Bpj���V�i���9fW�+9��n��b��|�
^?nǯ��@EEyZr4����Үb��nsJ���Y[3|ݺ��b���覠���z��eN���Xk���"�.z�)
Z��jKuklcA�`�� b�.^���؉{�j*i�f|����<w�k2"��n�����z|h�YTJL���烿�� %¾%̋�����d~͑c)-2z�`o�ĺi��kBe���3�������$&$�Sgw вE\3yƀ�M�(ҙ�~F�bL�:�R <Τȴ��-H�X��*�hn7^o'�m|~����&�Jq#�ȉ��~��y�Ǐ���k�y���v�3�<s�%����������x7�(I�;-�����H&�`���L������^A�qS��b��H��.��id�1�y	����B&O�,��+6~�_�Nj�p�7�:�C�z꩏?^	=�����a��9����h8�ֶ��]�/A���o֘aA�oD�$AㆨȝJ	�RU/�[�?�`x��X41��sWg+���j���d��^xa���++/��?8�����>���?_�{��l�%g�y�aP@9䐂�gkW�k�eE���.�O���g���$v��d����d�E����\�x1�N���,��V�1�@i�6L.{���ȬÎ���������.ڷ�^g,��	���;t������cO!�Z�b9U���?C韞�#�T��=}O��� R�'�RB�1s�b�tR$�/ځxDo�QG��2
(̔)S��>�Φ��A�_q�^x�!����@$i��S�4-U<ɐ)C�F��� ��ZV�)��Ŗl��He��r�¢"�w�h2���LR��)l��o;lj��!�u&�;G���!�_ڑ��0_�y��,�VQ4=L&F2���Jp�fTo[�.;欜���۱+h�'���'�*��q/��g"s�]��c(��!�OL�F�2�v6�4ٸTA�:��=�i�͘�E��r2N���8l�!i܃BXu<�^:�,ؐ�D��G�ㄱ:��� U	*��i#����fB�LPi���%F�9D�A�'�0M~@��R���G�pMt	h(G��5��I��L��j���W�\��K��*c�:��V�ؘ�s`�δ ��v�o���a�q�Y�.��͢�A�S'�8��Qg��]eF	�'�N�85\��3�Q�č^�t;15���=.'�|��ןz�38�P3�@��k�Ĕ��%$�{cꍬ�K=P��ճ`4g/N#��Axt��PiÕ�i��3�G��9�QV,.�W_}U��]z�~��믿�{��s̱N�����YJ&�1�Z�j������oZ�ЬY.������]S^�7�U,Q�/2 Vp�{�	����+y�wp�ĉ��?�쳿��o��/^8�	�{�W^���;�f�j�XƌW�W���"��I�&�q��o���t����T���{��i�J�%��}�rNe��i�FW�8����y�ޜ6mڵ�^w�9��|�Ϳ��o��c�A!��#�8���=Z�7b:HYϦB�X��q��!>sHI�;�:$�jJ���t�D}��|�d��FF��\�)�U�p��ꫯ��w�������?�{�}�z���$ܴ���.��94�C�N��8JҌB��Q%%X���HUҨ\IVQ,�m�{���ᖤ6>�Yl��'��9�'*����8>��~����:9��f"�ɥ,Y}�>>G�3<:��3kNp*��J?Â�B`T.u�����IQ�m[�&���JJa����-�}*����S<'�!��0���2�:_��%B$�=�l�����Ku#�*��F���:�R��������J``z"� !��@c>��`���Kc/n�f�㘀�Z�hjPWW���O=%t��&LE���Z>p��fi*���HV��^唴��nɀA��m�C��EvN=����6C��t���,X�0��,�f�� ���J'�Ѱ�aK��[���vUVT�ڰP�k��++:m�D�W����ɸHf=�lU�6��vfL	�;
���V��f��8��3t��������k�*H������~,.����Y���ʲ����]�b�H0!���7锵��˟Wh 8C$<��t&\��)ʎ�G�C���*�i=�5�~�l�QZ�B�\Z����N����w0:0��L���*洱q�ɧ��%��\�~SS�&�) N���"�;Bp��� ��3�ψ0i0��Yf��k�7�Q
Le�}��#�-[�r�G���Ç�,--W�`���BU�JV�õ�4cƌ3�<��O���oD?g͚5i�$�nh���!X���⊼nѺ�E��)����ͼ��Mpb���ɓ����È]� a�.���d�j=�w ЦԐ�������+�8�G�8����.Aϭ�<�C��������--����)	�55�D!K2BU3��L�8�)T;�jNM�� `r�z�>�`b��)bVRe��T��P4�u�5לv�i��rZ���{����Ղk����A`=t&�b� Q��&)��2�s#���{Y�UW����pcJ�h9<�,��P��S+�s9̤�!�I�b&�3�������e����X��F�o��Ś�J&�	����3�Z�U�<a���$��7�t�F8�PA�q|�,�9����?ش��P�Kъ�d\/֤pHYCl���8M��Y[ErO$��?���4�W�����v&C��r���BY����[@����*yt��J�|}
Q�6�ij#���/ �������ǁ��vZ�_A0�|}PUR
��]}fT��[����a�� ��̜LA2Q��'�$@��Nw\ffO455Y�e2����P'D'"Z�������Y��D�S}��e�����]��@H�NQk��
�b�n�gՈ�k�B5dDDP@�/).����p�;���)��R�a�^���'�|�M�J�࠸��Gh�ee�5�$)'� �PM�_0������[��b�K�q�H��]�#G�/�Z���2����ǲ;�����G2֔���˗o�܌v*+%m$O���Dd$��.\�H�VD���@nt�������n��2C))��x�cH�䒊�Θ5��iB�0e�K�.��q�7�m/_�s$�6�8S�'#1@�2�hU��B��PH�;ȅ�p�w��%����_�ޓW�^MP��Ѣph�Bޚ�
CATG���0S3����#����{����ݸi�����
�Vi4�j�ͽC�����y���'��x
6�N,!��kb^0���菆���e�ˠ%Z_��0# ;7.^���O>�o}��G�~���r,]�!��hݡ�n]U]�0Zkr)�#�;2eӭV�F;�uz���a�h��!/&4)!O��B"=���V�Ar��yb��c>�|g���0�~�_������t�a~��&cd�|�����Y	�ԓzݺ<C���d1}͔ڴ��p���T��X�'�$Va��)I�T�)��t��T:��z| "�{��FzT\\���	�niF�Q����Q�3'e�������;�r���HGG&㥰0/�&�.lT���J��l7C94��@�$��>�z��^�[Q?�d�¸�M@��8QY)�7Rx��į��}N�A6�OdM�l0��	��b�1�L�İ0T
�R��5��)��H�2n�r�;��Z %�6�1-�:@�bɄ���4$���/��zK�EFܲy��8���_8�X-�S(��A_�5���a����E0�!�!���N�@V-��VYU��ڊ���c�d�^O�Tq�ki�`
K�BN���mm��Z�V23���`�S��%��im��P�Ǎ��ɉ'2����߷(V��@�1hx.ƐzժU�3��RD��ڼ�����Ã1��SXP�����ֵe� �G#I���Y�4$���`/�KO6�i�(�T��G.C�G�E��\����4�E��x�E�0��褳̢H�D�e�C��0�U��ŋ>$�P"2���r��vhskW�<��+,��K����b��0��v��0� %|���y�#F�1M���M�ǌ�>��3C�����,�+O>=V�%��m�؂Wk�4��]ӄ��Ze�5k"�$w�"Sz�i�g�+F�;�!A`D$�HU�N�M�E��ơ`_?�dX]����˛U��hLּ��;�=��"oCC��WX�p!��Z���1	ׇ��3R�68u)��|�i�%��G��3�VnL�`%���L���V��E��ű?i9	P.��e�_�c{�=E~Әa���l�<�΄%�$`
4r�>���At�$I��@[⣲ i�
�!�x�[GcGf�>�s��"����e��h�k��~Mb�p�q���F�8_d?�%N��6�3
��V���x���M�⨯���n0�Y�--�Z6�zq$@ܙ�ui�*�-J���B �Kb
6k��X�}�3ۓ)�4�3L/&�R8�4��+�(�J���"4�Џ�a����E*�����e�D��c���DŰ\\R����%;]Vp�xb�\��5pM2l
�
^��=���W�+6���%���y\�3�^����ԍ�:�,�&��`-���n�F)���+�/�A�|���@]�ہ��$���&�81-�]���V�W-�+�����ߗN_C=�6Ek����)� ��y�`&��K��zz�i�Ǎ}}Atx��hH ������'R�������X`LCe\:eG��e �D+ג%K0�{��\#0�:��I�L`���V;te<=�qH,�nrCS��<���p��Šy������Ep#-�t�p�ϸ�6mK|1*��D�}0�O�9s&Ǚ� ��_dWxe�F�����
|�ԼވE�K?&���˗�;�K�p�-5�)uh���.F&)J`����"��6n)S�pF60�x���lRTJs4��=�Pܲx�b6ŕɱ��ŀ�]~bԡE╥r�br�c=Kjq�P3�1��Sw���j�=;�>�9Y|����OW}��d[�0�>>�#�ʅ���@S�%��3����Ͱd|��4��h��WE�esr�p8�$�e:̔�T*SK�6mr���T�HE6OI�,�k�Џ�}�<1+3o?8b��l�x�`us\��k)��Dor>�;�F\�	~��S(?�
�����IA�	�IiIq{G��G�.K�C<Sġ��E��UmU���yA�8���#�I��C$.��2 ��?����h�䞕�h-g(2�`C�)t�L�_"��hc6gw��P��`���vkǥ�a���ik�L����➾~�+�L�ʖ}2�NAHW����A��˘鄟��0�>KfB�l@�Ip@��a��^mx.�fRQP�Y[Z���{S��	�"3�����c�@�����+e�V���G��G�1t��� ��	=\�]ej���y=Fu-�AB��ñ�
���c�;:�.'�oX-uZSx 4]2�"���`(�y�����F��!2K��Ä�	ňQ(�uv2�ť�~��8_ZZ�>����c1������tź����^�R@��ϗ=�n�<��a����;9}V+t��۫�/�)-�c�j����s�5�!��
ǲ�d`L�cԡ3[ɥp�#GԡM��p�'�̞�)�����#��`8�%BRJ�jst��1��.���n���Pk�n,�F�5�����iG0�)��,�1������Б(q��^��L�0	��A ��Гի�R.��A�n0`��ٙ�U�F+�Ci��4�@�'��Ol�	1O�	S?a�5[�b{e{���y��1����ݵ�s�L�%7V����?r#�9|���;��L7�)=��rt��HG,Y=�IX9�-�:zn��F4[%�i]4��B�D�T��\�d�Q������Lk%J��R���k��A�|"A0�C#[0��gZ��i�z� m f���e˘(� 2G� ��$I��Az�����#�}��g�B`haF���[R�[�B�B�7�gh*�-�d&G�O!ͥgQ��9)��E�)K��I�3ݷ����5�8cQt8j�r��%8%c>��0()ӦRUZ�e�gɬSZU�5[���ٕ�aN�!�����c��O��XE�)q����]�V�T�O4�)8���F����6�44���/SC���ue�aR��M 	h�f<)0?�����ڄ��P.'{���0�un�{��(-�[��H�_m�p�L�ь��>2��a|	��k*�th�gi]Cc9�����I-X��0h�U�4�`�m�Y�b��s3:��A������r���˦MJ�VUW�/��/�V =�4V�en��xDF{���7%��J�x.�ڡk��O2c-2�x��i5�E����c����,^9�HV�'�$Ԩ-�f�<h�6Em23}f�	~�����˪v��,�x;�ǲ�)om�o����O o�a�:�X��PM��o*EF���-Ǎ�D��_��I��$d~�ڛ6��#��nr}���I��ns}�'�o�M3����b�u�l����62���)���ib4�����TF��f���Wk嗚4[c�9M>F6�Y%��z��"�'��L��YI�$��14ƞ��$��[��z�:A'R:���jn}�� ���Y,6�W�l;o����'p���<��~2S\04��qQ(=���:�lP�,����!:;��6A��-*�l83,i�W����!���`��V1\�Z�i5��à�7�x��l�UM**��̤H��X$�1�_�I�h{O ��{
�}}B�놁��7�E�b~�id���	<�����<�'A�W�\)��0m���'4������kqMu�0�&�3��!î�[�=�L����F��AY�Q��tC�]"��I��_�!7�����1J��=��i�#����g�x��͛�`�SO�)��$>d6�>�Y��&D�K)Qs�␢xă�$d���weq$1ȁ@7eY���߉�J��ԩS1,7nĐb��Z QA2��������%%Ie��pxXU�YV�'�:$���vxPtV�֝��W���Ht[2�V���lٴ�il&���Wۃ��aÆ��:L4]:�1�<c·3.��/�	�)P�,�F�ڋ��$KJ2SQ`锹�%!�9��AS��r��A�gh'�^�D�� ��Rx�zzz֘Y� �7�h
rJ�w�Fɪ8B�a,-7#�&M��s*�,3�:�8|_I��7�-�d����J�I��s�囿����ԠHG�y��o��y����v�_{�?�aJm�����|kwl�{M@�;��V&5���T͹���꥞dٔqr�xz��}4��uu~����ą�@*7��Q��J����$���nd%H��x%7��OC��	���r��C���5$L}3N�L�0���4j��,�XG!�{�A�c����¤/�"���f�u���a��n��W:��<UUek�n6���VC��8�WóMI�0��Y���cr3Ch*g�#�����f��p
���e�K� �J�3pL2G.���O,��`�X,�p .F���7k�B
O�g���d6;��{�A�i�č ִ�e ���z�����ի��o�lc�FwA�
 y��-4�k���RY_�nf����q��&�4g��d�?\�+�����0�觙o�n�J���C�+=�4�p�)�p3j�!7I9������ކϐ'z��DA��t�*w"�Mu��Z�/���M�lb�͋������q�n/�1��e�9>Cߥ�����'h����x/S 
pM�`�����G���'��0J�e��m�_�Y#^.���n�:|ţ15�)3`�t��e�/_N�mt���銆rS���q?|f�,��1�"ΪU��o'c&���	(Rn� �0I��3�٬�^mX�^�"]���0�9k�@h�H�h�����<��T���@�KA�ʏd
(T�of�#S~�w���΄�jV�CH�C��na��1��p�Z�-R���C����Q8�;dF[�>Ym�����L��=�������|�m;X�}��0������Ue��ͨ~����$S  �7�+SP���)��hN4�f4�*@���F���F�N#-���fU�=�)%�4]h4�Q{0�	h�"u�vEF��i\<a�X��h$���
��������8���#��nQ�)	u�%��
5b�(3����5��ܚԜ�O��@mB����ɺȉ%��餸`dkaT��^sB�IO@1���m���X2�8E���oP��E�>LFkG�VqQikk3-/��a�)��FW�*���0�L�%SG!?f�>3�
�$�e8L�� tbXW��G�|^?xlD罨��t9������Q֥Y'4��H$�G�c�^Yv,"F*�L�tL�0��0 ��ș]B ��x���
A�+,.�u:$ ��X-�|�%f��7(�vI�����>#*�T:�Z��J<(;���p��nD*˭� N�6�vu���:rd���lmmok�
�t���H�� "/��v,���ZCm1Cn���X$���7��x��^L�<.'$xAh
���F�S��0�7����)�$��<�M���)�+���/��a���0z2�jw,)/þ¼;ܮ�`���U*y����,��� '�C�XHk׮5�=Q3��O&�P,��N�P�f>��f�?]�tH.�q�Rd'}�i��1S�R���
{���i�Hk.:c�8�t?Q&�eq�LbŔ��a����֓��s)�� �5�;��$&t�X=�D�Q�X�MEs�i[�����;�������ܘOٱ�˓� ��,�ך���
 �ï���f�`��I�0�8+L�3�'�!2=���(oFF�ȴ��e\P�����tJ^
T�!���*ǿ����V��V��5����6k>����>�[3�|)#��АL���Ɏ�v�JfH��XQQ~8S��Z�%AU	��.�w���A
���&p���)��xZ��y�"����!I'f�-�͈Ht�W���ȣP�
.m�hj��%{G�!�G,����dr(n��S����Bљ9s&��M�6���eTژDw�T-@2M�7�G���W��)#�{����j�<F�.$��<�a���bI:8�Բ͌&�T�S�L�gA i����T��7�]q�ԩĚ�5�:9������Z�	)A��g4��'���/&"
=/�Bh�a�V����h��fn�N�npv�u�`ъ��m�M��|NA�UD
暒[u�����ѣG��+V0($��9�`8��ə�+ڼV��9�K��z��1��п�8&)p�.N�b.p~����IIE%�\�f�|<�%-2Ql��'Ƙ�<���Թ�{@Y;9"o���,O�Z+"
��23M��Q�&۸q�59�T��� (LCԀ���x4!=`AG>�xz�ZJՈk�YF�����M��M��jkk��1���EU;�5��E�TΑ��s���F�r�E���\�:�U!NӚ�H��k[���At����1�y8�`#�R)Q�/�l��C�̮�h�t���$/�ɋǔ�9�r}�C�u�,�^ߥ�)�6ָ�&�Rڎ����D�X�R�6�U�Rh�bx�]�]��������1�]Zwv.��w~���?��T�d��GFL�����_�?3���fX}N/��]�)����s��2M^]��#T����e~��eJJ�,���z�)+)��w��U�I�Kr9�f���Lh�!j�����F�eX[[���`�j
�ӧO;�xC����J�pTVf$-KD-�>diq�s�X���X����/~���U][�p��xܩ�[������#4��v�aQ�+�t0��Hh��a�������m߰���l�ɢ|_Ӻ��qn\�F��p
r\1���t�;����P2z"���h�j��<�@��i�6�`X��:[i?���/۟�'b�E���=����J@j{{$�k�І|a(��G]��޴q���H&b���腈)Ib�m��v��t<���K~h�שu�z�h0Á[���?�m�$q>�m�a��#�e�z^<��������X\�aq'���!S�e"�$���j5M�ⱈ���|u$�y>D�+�ErM�,���Kum���i�|��H,��,�(,(� ��Hx��F���l�TQVRVRDQuS����?8v�f�
R��8���"��S���U�'���*�<���f����.r��j��0C����NW:���G����,�auz����7y��.Y��M[6��;��1,K���dl�'��K ��֮_SSS#��t"�4�:��ر�[[ڙ.ȄIJ*��$�ZB�Q 
Pi5N$%�2�B4�)B���A�$D!'�����ROS�%�u��;ڻ��;ѱa5)��ބ���m,��,X��9`��� �?%�J�!1}}��s�l�9E�r���m����$�w��g��*�m��v��e�J�����TC��#S�>cp	�
�8(.T���.����J8VCC��� =�1w�y%%%�)?H�z(W�B@�#�юĐ������U�$h��'$ $:��RՖH&^�%�|a�7R�e�?�e�I�
zE߳A�a �G�j����HhHőv`��͸��#��)�13�AjX2̪��sԯ#~���ǔ?���WӖC�	�hY�W�����4y�kh`����C*�$�#31G�Ce�ϤY~IY)D�<�D5�� �ل6	B�`t�cn���G���T��an1v��"�������Ps�8ъp妣�FSSSb��UŹ��٘Z
?�qo���?���g��m�g������Z��9�����d��Oo���%�y&!Wby�/��Q��--lu���ڋ�M�$�27n7[��؝c�\�k���=���q6C�J�Lֺդ����s]���|��pn�%yđ�5͸����>��C ��fy���d��������w�K��0sOȐ�#�f2��n��1����tĘ!�8�0r^f"g�MN��f���Y��X��2�{,�����#��͐���[F��Q
a,[D��ꏷd3x٫͛73���1,�ȜO��� �@rYF��g1}7�%���6�,لd�;eJH��(w�����c�0'���t�٨j�8��(�p:��Oe^�Û�%l��=�	����\-�n*��J���G�!���]�深�s5�����h�����܏�Q����.~M���َ�Z�U��f��n�����㼆�L���nҔK>�AV�K@@�>]#9��l���8�+0d�IE�4�U�N>ޘ1c(ܘYjl3�$ �9d�&�d G30�f^�n*�fIJN�� 	�� 	4��M22����A�L]���kLp~r_f�1��򼙱\W[By�ɢ4BP�`d��Û��%��d�3����t��bq	S��򨮮�HہTNٶ�CQz�l]W�r/�|�7X�]���y2i$�̙H*�C��[=e�G��F}�:�z6�RT�y��[�!�:)	��>��T�7��a�ꯔ�l!�WqC��?Kq̲������K��{��?�*��_t�����
_ɑ��Q�-_�Yh���!�������9������<�'�n���߭���t�|bD�6M���ŉ2h� �� ?�zBy�V~N9�6cH�p��gZ�ji5&���|��3���l��!�D��"�|P\+�����6O�����5k�Ђ�{|y^��D$�)Ϸۈ�������?O�zl5Z�6�7>��^����k^A�߰a�A��ձ�݁�oe䯏��#�36���%�!�(�W�4�����q  ��IDAT�GH1�h����ʖ�Jj���������c��~}�t:���	"��֨�W��Mػ�Ꜥ�[i�@0���%�8͸ݾ����΂� �uY7����sc&�A�8w���y�h��!�"�!�\��)K�iΈ�hf:�scJ�:3�w'm~*��؉�G;���G��Q
��sXs �>���c��9��Ox<f��}��fQX���3ẉl9��V�Z�r�J&��ԖM�2Ѽ��e���6O�����\n|%���6#�[3Z�Gf�}�ش�pK�a���cO�~��&L`���2 6{��c���f�˯��ju%t�a`Ѭ%�+�RA9��5�a�@�6�5������o�8�eU�l'��E��g>����s���d�V>-..���e�O�'���Wmc����}�����/���+� -��+�ϟ��O444���Ǟ|�I�xkkk�>��/����5o�q6���{0�N<�l_Ͽ��/E�����ɓ'�5
��~�-��f����.Û:m,,,d~����ԩS)Lx�޼�~q*���료b��I�:?�RJ|I�5:�3$�b�����d�CX>�B�:w�!�����C�p�B��ehx�� ���c�<2�wT4�k0�`g��хn��[쎙�?��̡W���=�RT���vw�T��ݭe!�g��>c��6�>�6�o9 �$�	� FK����N�[�1v����Oc��a�],�	���V�u�?�T*�����7aA�$%V��O���-C�jA������ɚ�뻬��V�A�$[S�˗�x�~�T-5l��^�l���1cv(B`�o�����0��P������9���;f?}�����Z�z��8PO?�tP��n����w,��￟hz���k�ԃ>����cUﳯ��a��v�mh��O]�h���_��'K��Ñ��o��=����Ňzhyy��5k�#���J�I?��On����z�l``y�7�O�~�gbO���{���X��?���w�Y__oɺTIL�����>��P{kk��?��o|c�ܹ��u�]!`cS��?|�7@������^{A�X�b�<���Լ��K�.5��c/�}�=���G�����2�T{[����Y�g�رe��x��P�,o��*��8C��zif$#�vc�7�?��7ږ��N°n;��!	�;;����n�l��yr�"�Yl�U��=r�$lkbqb`K
�M��ɍ��`S�&2�]7���@�����F�?���"dU����[`ؾ��F��g��)�� ����TL 1Ux�EaY��#���b1�.q�%1�&���T2V}Ip���bQ�� �aV�C��wV��a)��V$��4K�ȼ���-���ď�=xbyB`1�7Df]tQr���0]��͛7c/[fG�/��2�bvq��k|��)�o��"��n��;S��MǛI݆tlZŐ���wv!��dQn�!��Ln���'M��6����Lmlk3�<w�s���w�O莏d��r��j�����g?h�ǫR	Ih�b$�F����7|��o]h^��М�����'���+�[���<�C~��G���G{l������ĕ���_~9�5�¥%��[6o�۷�zkEe�o�鿹��{�Z�W�\9b�#gl1Y����{��f�f������>��c����+!৅���<�{{{}��o}�[AfϞ���o~��.�袳�>���C�!~;�����s>���>����}��w��k/�f��y��.]�����=��#詬,ok�0a�o�ۉ�&A:��#O������������_��W�P@:y��w� a@^9����������2i�$%��v��r'����&����:
RO���=���ꠃ���	1��rٓ��5A�V�Z���"�|����c�AjذaP];��X�ڴ�}��{i�K8H�>����x0˾��P��Q,��y���|��n϶e%�)#!s���9�gADn����u��7is*�V��dp�\�h���^�J�0�X��f��ﳏ��lz+�9g�����^������zF�G���k/	V�/mhr'���>؂�4�\�b����3�2}�I��}g)- =P��>��iӦ�F�m޼yO������􂑷x�]s�\^hdSrw}���O�i��CX�.Ff�O��I��7������ � �է�vx�{ު٤ӦZ����kU�����Q��5B���la��]���aM���\�")�xIR@���.h�T^���g��4u���uם�]vYUU��E�&L��'���M����
�,�j�I�)dO<��̙3��?��ߜ3���l�	2ċ/����Z TՏmh��
����#�4}d"�g������kƍ��'N�ȼm|�׿�u�G��){���Į��~���;����v�}��[�d���W]u.3T�Nk<D��������?��<�ȀV�-*��~L�?���9s�r�)��x��{L���g�}.����^{M`�J���� ��[�l���y'z5�so��6d�L"PH8�ͳ�^�n�:	�s�9,jl(�+^���O�;w��^A쿬��~���g�q���Ì����+�̎c��7�x�뮃��¸�6m����V�ˎo��r=^z�%\��L�:�W���B	����g�Ou|�,?7���<]0>�>�R�p垌k�c󫙔H�JlU��jᑂ����]�}��?'ڂ�|:���/`�	o��C�T"�O�Ӆ֨%aI��d�H:��3n��)9��گ���tm8X�A&x�a�;p����I�lL�٢�[�7e�s�p���g����Hw%��]mp(<Ȱ�Ѻ������}����C��| ؎��_�Wn(�9���HtP=�Eƕw	�A���x"�P�����A>�j�~�_@�kjj�<y���`#1���?v���Z|7�F&��}�![�ЀFr����fx�������Yr����?�QWW� RJ����s��)S~�ӟB'���}����|��믿���h������Bvt�܉hL�S0	gj�Ͷ���Y�BaUm�ʏ>M���hM�����֭�g��m����+�6�>4Q65���r�<́5Ņ]�J�<Ϣ%��>n�����=�,�U��;�v�aI��1��7b����B�ǅ^��O���w����,���/�8m�T1�7o|���ha���g�}��Ԍ����KK��ν�'�p���=fL}Ii1�li��������cӧM��QR^���@y�Tl0$-�=�%� 5HpM�s���%�\r�9瀵O�:�bza{P&t�7�+Z�����c���`�i��\^<Jv�u��7Ͼ���2v�y\���6�a��O<~��W�s?��ߝv�I�xw�����1����X"���
s2��G�ӦL�F��K�#���|?��"�G~�[n���/<�<�ikn.+.�:�����W��sB�I�V�\����c�<"���D"�]R�c ����5s��|�a�ü�� ���#�t⬳Ϙs��t��q������[~��:Nk��J���rk�S,�j��d*��������@�9���?��n�A �}y�7����k |��W\q�5�^u߽p!Q,���lDHfM #'�<��BD�a�^�Ǆ|���z��@#WF����gAfmoo'ps`dk���%�#�����mH�"��jQ�Lq���dv@4*��E�ß�H�)�
|e�wwvd�&�_n��E�4)Rj�n���	�5KcGO�.���G��v踂R�9SX~4j8d���l� y�pX_9�$��ѣG���'���������1�f���́��e����T>���-����dނ,����H��K�.���Q�Xm�6�2�b�*�aGa;�{��rf~�_�/_
�F�$�'�*�ؓ�4��%ks�}9f�\�%[xp��3O�L�1y���M�!׿�=ܡ�@���K/ݰaf��c��r��c�}��K�60�{֮]�,_��7�td�G}�ꫯ����B@XO;����׃/��x�~���7mb���;��o�jԩ=��sѢE���5>C��*���Z^��p�AX��=@)<묳 �@:���0��/��~��ǘ֣�:��oƸA�$�����nï��ջ�Ub�y�i��q��{�5m�3�pb��
#s�G��PYp2��∩9��cq������[���xЁ4jԨ�O>=��gA��w�qF�);9�%5���M���O�ś�����
�G��©K�h����{����������b�f
�c����]�͛�'Eˊ������x.'HZ@I��"�Ъo��Vt�����~v��ZTE�Ř���Κ��/�x��Q���\S��5f��5k7�r�	�mm�тA��a�twbR��� ��jt���.��"���z6m\1�E��hlt;��z�)L8�<��@�!Oड)�^�����>^v��<��6�v\y�}�AZ������V[�?�/�hL� I$��� kRt�%U�]ሠ�c��6��iӱM ����w�,��+�X���>F�΢Y���!�45洢�b���C�*��Z���Ęc�tvv>��#�-��D����q�Iwh�����#��,-�h�W� j"#a���E�5f����̯���P�� �K`��6��I���t}Þ6����mS��&?ģ�x4��/)w��m�J�zz���9��幽>ÿ*�_�uw�
N:��g���7�Ñ�{J;n_~~ҋF�F�ӕ,I{�z��U�FU{�a�lI;[�[�W�3���;�x�������n��'x�F(�HC�'��O��/İ���믿��=n�8�:�JX�y���#3�j����} ��P������t�~��`N�{X����e�i���X��vĕD<��ҩuk�>���P����T��v؜9s@1MN�(��邔�02�oH����@��~�Pj��͸� �rEe�if����Tv���<@����;DÑ�W��Gc]��T�_��3}ziaa�����"��7f��[o��g?�ٻo���N9��=��죏;~<z1n�����uwϝ;��{�������C�#�h��~h����V�4��5�,����7`҂�ν�i�:,���bpƏ�	N��?��O�珸��v�Q��#����g��`<�g��<��8� �������;w��c��S��`��������aȺ�zE�46�4?��/��Ts�Ǐ?q�$<+䇷��qd���/���� �׼�����
�=���SXT���W�z̉Ύ�����3�8�|��w@4�hԮ��dٸ\�t,�d,fs:�s<JXYo�ݏ+���c�����f��>��Q*QM�2�Ѐ�֖��}4q���\|��x cS��cQ8�v"�bˊ���s�)ҁdR*�����tpp�ƍ�&����������F�L)�$�7�xS<cƌ�O?=�OM_�\��*G��Ц���<^}���S���B�5k�	���� �a�e�W�ĊB��k���Ǯd�a0lA�qd�b
Vqx���ޱ��)��@n�	g�W)���޾LƄ��wl��VUcH�������~��O<�o]�]�������4�m��ƣ3C����򩯓����5J��BD�!�f'hl�p�o�1�a\հ*>���}��%��;.��Jw�� 1´����֑a�D�Ɏ����K&R￿X���So��կO��~��s���m0$û3d�,
�ho)w`��tl�U�n���Z��gR�b�M�u8ҡ�F,Flm)����L
ɼIɰ�8��H�R���v�77�W7L�f�/�ko�?�>����vC�q#G���{.mL?dd�(j��z*9��G�I�t��p}.�&(��A��e��j}+�Nh� g�XJk��Uz/�kzѢ%�/��~p��GSdY���\s���p�XwwoKk����l�����u�GQm��^�M�$��P��*��JQ@�IT,(M�"R�yH��j*����l�����$!��������8���ܹ���}��Sħ[�p�Ǌs����|dY-U*S~��%K�/]�"���Ι��[o�1��	2�W�X�}�v���b(�Wu�4m*^�u�Vm_	���8�Ǐa�?�D��c�M�6 7�Ml��*O�Ųw���ׯ�`�5h�@���LM����	p���i��� ��={��A��UK0����У%�r�@[�7o���f�]�v�.ܲe˼��v�z���իWC���X/t`ǎǏ;�K���Ѷm[0<���կ_b@݂��n�{��D����|f0��g7�\�w�}�վC�jժ���>���m۶	�KQ\z��������o�>�#�g��l=�bXHJ�*٬eK��W_}��1�5k�3$61�M
��~��(z��'���'`���GD`��qz���E�F1���^~�	�;�W{��9�ᙏ�?�''�,�E~���J�*���`�*���\�إ��𼇏����CB`s��+[�VݺT\������@���r&P��G�1�Y�5�b!K�j�}�F��/\���\>z���C�6l�`��eK��wûGFDB� o�����`��(QV����K�Q|A>�@E���Ab��b�<_(n�����6^�Y�o���˗/���E��&/��������*^���GDFB�1��+W/o֬�.D�ڽg'��9r�d�9|(�X��~@�@%BP���{�`pqA```�G��?�C��/�<-5����b�������[��Tљ�R����b�.�z�j�˅\�IaW�k�de<�4����5.ߪ݃��S��RӺ�w���#���-'/K�0ڌ��M��nv����
#���K9>^��;�yy�ಂ^��-���U������<�m��=�򟞒[ü�1��;4U�A�A��"~�9s&**��hthJ��5��J�TD��@ㄼ�i�Hܗ�Oea��T(��DV+M��7��Wf̘��j�aJ�:u
��ԩ36l��c{ς��_�4l�0�/�i��� iP��>�Ɩ��\s�СC��ư�2Pa��iP�4���k[�jՔ)S��S˔	&�o�ĉ ��t��f��W��m[���8���>`�2�µ=dȐ�{�H�qeĈ�����㖍���	�\�hщ��Z4m6b��;w�m����Ɯ\|b�U����.]�FY�� ;Myy��P����k׮Q��Ν;S�P�/�$^}�Ո�J���n�藵k?�������A�BCC�͛��0����/`��}1Fx4b����x5_??��[�C��5�f�-�s��Dk����������7oʒ�!���/�_~��eE���N�4j�(�O�CϪ[�ޮ]���� �ܙ���Gpo&�/����MNA���Ңxd?d�֭[�MlwX�[�	���*����O>�}0=!Q�A����0����B�0	J*p����u���Ij*f">
��<x0zJ944��; :ᡸ2'3X	�ԩ���%� pf��=�����:zL?�����c6aa�,���
��}{c�ao`�A�@!Kx����w��(�:�|���M�*���:u*��7w�.�Ɵ���ӭk��˖=zt���,�虸�x�賲��VW�:@<��b�;_H��c��u8ǳ ��9o۹sg�*U�.f�;�G���C�E^p@�fΜ	���=?b�|��5ݶ�N���cbc��6c�@Bd|�v�*�txM��3,`JbL�>�_�k�9�1���+�UH��-��"�/��(��SO�(�'DkЉr�V-�.�1�רQCQ���߼y�ҥ��X%Yg]��Me�"5=�ҡ�P��X�4>��w ��i��?0P��'�%]��q*��9J[�,�O�Pp���d���|�;��	)�I� b
Y!�W��6��{����}��ͅ�OV�Y��s-X�Z�B>���K?%/+tu����Lz��+s��Jqq4�#��A7�<y�ܹ�<�W�KL#�j՘{eBC�u@5�D�#�B0kXZ.6�\:t@�t_�f͠q(�����~��g@��1�f|����ٳG��p�B�U�%�DJ���%<�]�f)�T��`իWC���6 ��+�/���n/Y�*T��
<�²��b�"��<b�� Z0@��� �� �<�	�go�K��0X<�{�n�D�E�V��,�4  hsJy�w������;@��w�WZ��=��?Eè�8��*_�d���d�q/pG?���E�ذr� �9p�@�*U�+����Q�3q��	�O�,�
��xq��̌H�h�<���;-on��	m�U����cp��x<7�O����X�gtllt��HO�N�
��m|�/k�χ�_����c��L���&M�0��բ��bb ~ni
L��j��s�W���Ͱ��==a,�:�5v,���Ag�m���i�Ǎm4�8�Õ�ɓ'�m��ɓ'	ի�]�֋�`|����%}Z�6m`�����jb3�g� ��gc�qq�♍1Fk��� u����VČ��J~EWHXl�޽*WY�rec�� �[�=�{�r�@AA�a�t�Ё�K��ɴ��1iYe���T���s߾}�ӧO�	��q�'��'���`�Z���;4�߭[7���),u��\��Y~~~P���9��V���1QtMW^5Z;n�J��5�!gub�6�0bn�O"��ٝ>��"�
����f��D���ַ���-&c~�Z���t�?�(�%?��On dSH�*��y�eVfm�)���=c�A���ep�½{��ի=p��g��L�g6U��!��u�Tc�S�������rә�湫+kU�]0g�ڵ��2o/Oƻl�T��F��͆�7�͆l��S��-x�����ˊHC��.Yq��OV/��w�9���6�ͮ�;x�\L�Y6,��׏H��gU���T(_i�O?cb�5�g^4ժYK&����%�Z�j��h��?u0�����[��[��Я
��[�UkT�L:!AƜ,��-7+S��(�
O�\��0�?�<'3'����2eB
�)7G�fx�e�#�ۂ��X��̹x#ZE�Lo0h���;�ԩCӦM�C���v[q]���#T�7yҧ��9�8j�ș_�ػkד��� w��b��*����?�S)�]�4e��qc�H�1�i/ߔǜ�z�%�T��8�1�N��:11qٚ��խW�Zu��V2���KmZ��'8�I�6�ΞS����tR�*	,�B�Pk6i*S�23�n'�c_.h���ɖ-[%�<NI-_)��]�~��M�;u�5P��I�iQ�\-U�n=�4j�T�rZ �A}ڴiE.�2AJ�L�F�"�,�ph�����V��i���v�<(t]�<��\�p��2�ܙ<�	{*�y)�Ճg^�[yM6�j���y��X�\%�%�~����� qEf��#������T��r���|������_�Ig6��O���Lr!��XKv^6ȭ�dai�X�G��|W�]���䞾~�1�DрJ�	��f.�Pȕis�7�L����'O�FEKېo)�+��x�;/�n�� xB�4���7j̒��C��C�nm�vd�Lf}��L�������+ �W�����r�Ud�\�ւ�����!Pr9jѼō�7�e<볘̦Q�G�5�?��\lL��8��@�r������eg)���`���\஝|sZ�X�b5:���ŗ_s����z�y�5�tX
�b����T�pJ`��G�`p��;@*~B�B�6�|���>�p����޼�my�N�B%�9����MKȕ�s�΀�/�R�\�$�#~Q�+G���:U�Pf<IO~��?�_�f:r�4��lU�&���_h닮��$�%�.f�ޔ��,�Xk6�=|������f���Q��˃�;.� �z���[O�h��r[,���-���AI�>q���F�/�7j�1{�ɓ๱��W��;��x�hAR �JNN��)������汶�jՁ�B����+՞��{��
֫,i��z�yz�ՙ��ݏ�`�?sƨ^���L��	�;~꣏>z��77n�+�9�k׫Ƕ9E�{t�B�p�J����E����3z�۴iS\������M� -�W��eʔ��:9�L����F�F���R���������/4)thZj*y������pS�\�rx4PV>�YO��Xv�.5%�ŋ�;v��a��ʕ+���:�n˖-l�U+\B��(�72Z�h�������={`��9s��A��O�<�dɒ+VL�:u�ƍ@�1c�H�� ��NH�f��O���aaax߳gϲ�	�:%�+�/gY?s(��s�s�رk֬ٶm�wӦM��Ǐ���8!�����B�u�ԩ��ֱc{|������u�&��~2q�~��,�}��s��1��0%q�^={�y[�m�/_����?,��f��m�����EÁqONJ�(�Uɨ*`�˝�f���'!ha{��*W������ҟHM1�v�H	�^"%����K�^�0@T#�b���ъ�a�G��"P�a�s񣀒�������"�0b�h8 ���h�y�<7��V�����#�����[kD���t����lV�]����!�W����A���+���$N̖���(�ïbP�sJ�K~��?��'B>� ()⫯����م�X�tiϞ=�?J&��T7Ol9�s��Mh�J(��!:S��Ç��aÆϞ=��V�5��O%.+v��ˉԍ7��}��s����(9��(���l�^�V�+MV���!-z�*�>��$Sm��J���
*ȭ*�l��;W�|�*$X�����Y��c��W�����jV
�#�tk����*K���I�J�կ&�i,�,@���O9ҍ�Z/(���Q`��B�����0	ԗB8�hCV���e||����b.*�����X�ڹ3��E%C�v�r[3���8
�`3`��>}��75L�A��M��c��x{xzz6lظs��mڴ�O
[K�	�~&�e���*�W���F���ѣG��c��mĒ��oaf�̠n�6k(	=B&�{�njZ��<~���n�t�֭[�	U����K�Y�ڵk-Z�ܲy���/��?Ds~߾}O�<����.]��	&����  �o߾=t��իW�VP=��᤯)�Wœ�@��>}�c����n�D����qO�'e��fA3�7o�^]�jt1���/��/>x E�> �s��ū�nx� B{Ξ5�R�Jׯ_^�|i�׆ k�<@�ӧ���M�孴�����7nܨQ�&�):y�����RH�s���*4��K׮UF�5k��ڵkϜ9�޽���x�7iDxo�?��q��+W�� �5k~�t�uU޾=�������A��ͮ,��`+p-̼d�}� ��ӧ>.?B�i�W|3����I�������rȐ!�b;�;�A`0:��w�WJ�V�xcAHH�o�1e�T5�b >�+J�z�ԩhd���I������`r,�l�'2�Cg�D�]~X�+PpY��d�O�d�L�-���O���6w� �ݜ�lV�]�� ^�5��v�w���f縹+�}��c��>qA>NT�p+��	zE�E/^,|Fz^ښ|Ƀ�#A~ � �;w��b��M�R'������:�W�{ժU�I�1C�1�+>��8u�TΥ[���Ӗ��O<�[�wӳ���;���?��J����x7mjQ��,y���ie||��!FcN�ʕu|�1��U3�v畵�B�3�b����K��ՎNwx)����X����`K�t���9$+u�g����J7�.����H� ���^[��+�^�q����jՒ�M��hIw���Y�2�g�s��40��[�23���|�kQ.:����4-�,�>o�BS��ѣ���{﭂�X�f��_���%-9����y�2,B��|��%�R�?l�0� �3��={6&�A�����5����j$����\�?,��+�;w����Ǐccc�w�z���͛�h���r�X��������0l��N�;�j�
�Q���"��;
�xÆ������cAA^^			��n:4��˗'O�L_�С�ߛo��`���ӧ�PiЂ�}�~=sf�2e�M��n�: ��+��ߟ���4x�`�[���W���J��������T�~}(���P�=_�֠A��B�s��Y�_�A�ޚ5k�o�&�X����ŏ;v�0a���fY�x�u�X�=���P�I4|��{�6dB�U���2X�n�>������0b��% ���~�mt;z�É�{۶n�$���+裝���c���2�y�&�
�t��e�T�j� �ׯ]� a�Z�l�oY҅� t9�I�"8p %%	���6.��x���Ǉ8~�b�ή�{ �ݻ����j���ɓ``x�+V��	5-�ǽT"�1u�r��xϛ7o��w�C@�ƍ{-��޾u��H�pa9�1>�����J/#��J��U˖����y��n���{��&z͠���C)����J�2�����4K ��`�Q�a豽{��g�5kF�6!��r�+R ��B�j�����
�z=��FU�8�
�<r��9�}'p��R圛��d��d�d*H�жm[�a�EV򐹦@�n�����&KE|��E�����������ޘ*4���=Sd=+�0�f~�Ym<�,�%Oa�Y�1����w��wGi�6��3A�x��V�s�CP>v�
Ȏ�xxYO���s�o���s�#d�L� ��^����>��k�3���Z!�[ur��|N��K�����&T@�c@����+<|�z��R�Ƅ/W�ߠ)���~*M�(|�6P��K�#T3O3̊n����^�v-��;�A��7n�����t�N�ٺu��#G��yh����G� �n(`^������Mǎ�0�����͸���/���_���K�d1�%��ϵ˗�m
�^�N���V�� :vh�?��w�p�ر#F8p�:~���J�@�M�4	&xLl,�v��!�k��R�vm:g�E�
�)�8v���'��k={�	�-�f��1d�@��Ֆ-_����>���[H�1���ޝ�2]�ɧ�JG*�g���o�W�1�33#6"z[��V��g��޽{���"/��۷���3f� � #��_�A)Sб��'O6rDS��Y>�8�7g'ӦMC�s4�W�*o�4�2���QQQ����c8p��y���͓?�x`�ppd�z`���^{�p˖-+W���bn
=z�8q�@ l�����ٳ/^����Ǎ��[o};g&&�� Ecfp'D�RϞ>���ӬZ��b��DY:u���ݸq�߫W�cǎ��n���Hq`�;t/qwK�|�t�Rb�h�g�}V�Zu$$��r&�@�V�,f١���������ٺi�[o��t���VV���S,�gd��d�;�8F9s�ݷk7��lٲ��u�������Z����7�^[�xI�n��ݹ��;�x��.�+{�칠�`��ZRƘ�c����jժ\_�s`3?���t��%:�~׎�0�[�l%	�S����OӐ��]����t+M:W��z�?_�B2�݆�B���}�X�䁎��N�O*�dv��&��&����&���={X"2S��$���t��t�O8�z,H�Mpݺ�G|�!NK��?x���C�Οǌ�������E (C ̓6�l�k׶��$�{�_��x�҅]�rrrhߎU�e��1ܴnB�چ���mx��)h@>�D���ϝ���������p�����]�(���`��RW��B#��;@�a�3�e�w��O�Y�n=4r�z��[S���ܸY�v��������.\hױ���7�N.����X1�m����������_�9s��%�|��E0f���d,�@&�+�J�y^��
���C���wY�^�>}�*8W5��`��H�%h������rZ���� l�@�Y���|��WY� ����s�r�XxZ��(d��{��s�!�F����1^�x��,��sI���o�Ë�Zw�'��3�W�h������*�\ŠM��aȐ!�/��&� ��)�'t�$(�yY�5k�ĸcd�W��h���C�_�N�/��X������� ZL�y�{��!-�s���7�|�z߾0�@�l�1�m�LlH��Y����#���-P�ɓ'CZ����ףocʕ�;w�!�(`��n\�yg=��޻wZ������!C Z��s��J�*w-qC�*T�P�F`ɾ}�@�� !�`�YY�x^S�c��ɔ
	��ݺu;�����}�����:u*�� �]�re�*UF���@�\�zl��%�~��1蘳�0�5��g��+�F�mDt�رc�
�J7�	[�l����w�=��E4iҤQ�F����:�ߏ�� k���A�����ׯߜo�lۼv3 �Ab"S����XS���Ǣ�i�y��O���O?���_b`�&LX�b���AV��n�:0Ht 4	4 ��GAXYYY_tZbb"�*�. ������ӥ���}$ء0Ke�KZ	���{��x�֪}'�'��ǽ;5�ֹ��M�T�,BV��@ �,de�ٳ&R�g�
�6��`Tȼ�-�\����ܷ�O!/Oض[{�{�27;���%���B*K띛,���?�����";�A�[���.B&�7��v<(##y QcCBB�:O�<	�%%t��f��<P��ʘ���/t���C��b�c����)(�P�"�9⡄�r��!2��r��Q^� [>08ӛy'��r�7o�?~�J��O���of�1+V����:~�t�)�&Ԩ���]�]t<����g��.�my�����f��	��<��V��.N}��k�lkJ�qJ���3$,w��X�޽��9H�^����UZs�Q*�߻�,�ɺ���fI�8��"�B]a�+��'��!�x�ܕ��,g�k�z֞XO}ɒ%�<�)E�0T�\rn���6^j���+�[�����N#��܊/�[���B���c���[�Fr������(��ii��xYtK�u` l��ݻӢ= �m1+��DZ� ��V&au͙3'))	d��Jɜ�	ЕP�%�Т,�7�xF���E

8~�8�\p��'���-�efB�^�MYp3?�aGn�����4P]�N���,I�aK��-q斯P����u��Kxg�`�$��y�o����k��,:|�]�8xʻ��7x�` 7n���St��w�@PX�W�2�8�����~hݺ���>�4�|L����-^��i_�wp֬Y�2=�I�

7�������Ge#�rŲ�@,���A��3�P�2( 8+#�{yxg<�������a��سy9FO�;w��Ԫ�x�~����^�|���_9ᓏ>�kV�^C鰰$��k���y3Kj:���}�$&FG�C�(պ{�ow����w�;z�'�|X�6eznv�k}��|�W�*U�/^4s�L��y���1Ő�Y�t)�=D����8z�(e���;~�XժUK�'��M���O߹s'��ka�9z����!H,E~A��Z>|��_!?`N<�PR�ҝ�z��1O�T��[�(��)F����w��_̥�'�K=x�ɓ'1�Z
����]#����ܗ^a�/� !��)#����}Zf~^^��Ð��ԋ��U\`�9|8��s�2*���{�	y;�B_����
��#p�"zEA)1Lb�Ya��Jq���א������r����!���TGn��$�t�a�	 V}����4-IARMJ�)��6(�Ç�`���iߡK��3N�����8�רQ�%��ܺukӦM0h<y�/�~�J�o�F���<�T*|E�\P�N6u������p\����]���I�In_��}��8�n۶�2l`�(���ӧ���Cʔ!4ţW�\y��]`����+<\��� ����\���~h�5�7L��VN�Yj���~��Sx#h���jt���Tv]$j��V��t;��Ԯ�6r�ݻ�п+V�|�H��0X��ñs�.P�x_h��z�ܻw�\�0ܠ�����o׮]�^��&�f�>}UJ�E��Q�֭�۷�0c�Oww*L@)k`�	���E�.��r���t���x�)?���]C(�e��`�֩��b1�NaX6k��w���~�`	{�� �,���/Ϭz�R	G����џ�=~?q=���#z#N��,
r�[5o��z���t)������[ܳS�N��(���Yz��gY�\1x�+�Ա�v��iii�[�nů���*���x�/��^o��>r� ^ǟ��K/a"�ffR�Y\�䅈��,!�M��{شBF�	��<�KHx��1�u���T 6`9�˛{Ԋ����8a�!����W^��������T�����e��������C7��`z��b��4��\4�o��6f7tE�.]�;��ǃ�H{�����_��v�P�A�{�2'�b^��2�A|q�;4걢+������-��'��
��|>JNԷ���LH��$�z^�=�F��Wt>�_&� U���DK�Ƀ�<=��0�A:7�n���!��K8t�g��*A���giS�-���M!��p+�|j���*�	�ﳨ?�_�ƍ�鏡L�Aʬ��Gz�%I�pc�S��;n�U����|�A/�����\��w�<�����M{~])�M�(L3��C�ٖ[�2�^�^f`��	̼���+0�_:��6����V�7�䊝L�6e��	М�\�ҙ H���||��@WǏoѢEC����o͚5�XB}ܽ{�o�>U�e��<������I=z����믿N�8�Nd��#0A>:w���Ə�4i�bذ���Ol�s�_��aÆ�<�K�ݻ0/ qbRt��ү]��r�@%}���Z	�l٪��Y�@�0ˀ��>Z�p!4E�>}��qq�o߾)��k��ԇN���h���AK�z���/��WeR��;{@5����}��}���1C\���5�c׳gO�6�1�JJ� ';����5�y�ƔI�@7U��@�x�m�0VN�:U�h�%:pͮ]�2��/w����U�̅�}��ъ�*уV�X!UL�֙3�B���ܹ�EUG�]�re�mbb�̵���f�R@�Ϟ�M�ƍ��mٲ%�/U��i`���0m�4�c4h�TXXX�-��<�2���:��9�6skP�h*��� .ZK��u��m�1�?` ��~ʦ��M�>=&l���΃r$��Z��\�?#3��O?^�`����o�����/Y��Ұa�-�7Xl�yZI:���c�%%%խ_O�	�jT�3��Tv��DDE�X�r����/W*
̦�A��ӤE�U�A��|�2ٳ�4����A>w��[���DÇ^���^�g�}6eʔw�}��w��m2����9+zF�|�A��B�0Y@Y`�8` &r�^��-0 _Hl�=`Rw���ĺ��	�I[����5H� �R![�蔯PA��$efd��tO�4�`-0�1�P2~<��˗1Lx/XD�^�k�������$�p����FW|��@�A��ע�>����+�	�OKk�~�*�,�'��+|u�|d��ɇ:2�"7Wg��X�#�ٮ�{r�>�.� ����|��c���� ~<�nߗ_�M�VO)!;���XR�o�M�+����|oނ�T��1��6g	v*�J���f�$�o�ԓ�cگ�^)��Ď
����&r(=N�c�9��P,UW���H���@���;�x`��K1��o߾|��ﾛG���F�8������T�,���  �5 ; �ba�%<<����s���8�e�O�ey*��UI�6������N�M��3���׵kW��?%%mܸ1м7�X>��l�J9�H�߿r�ʜ9���h%��7|�]��_}�P_z�~�~(p���m�P��S��lZ�n"N ��@>Y��~Ѝ`�gφ�����.]���0u�ؑ�M�T�1P@x�ŋu����hK[�ьx�={6o�ܪY�6m�4h�hٲe�����Z��ZS)�[t~QQ2RY�?�UZl OQuo�	�)'6��y˖lO�e�����ZQ�����}Wp�n|�V������v�ۧ���wq$�lܴ�6;�4(]rr2k'����׮S� \��/V�Q�%%�<|�0�R%�%��۷/�Z���@� OKK�.B0BBBh�F���ϟ���ڹs'���UN�8��c�VK�,,_�<� �ܪuk4 ���q o޼�f"_�x�OoL.�Ţ�h^�u`j|Ŋ��Ȫ��Z�
<�� [Ҹ���p}}k֬)֌���X�l�e�y0H&���uNNM,S�ʅ ��~�	3e�ҥ��c}ذagΜ��:t(>K�5��!\��N1P�&O������c��ɓ�~�qǶm@�'))h3�����!�xӖm�N��	(r��1�
\��2�}6�%^
���<IO?�?�3=��C�a�8q�c%�¥2b�"��640݂��������!::��:�����+��v�wy���]y
�BK�%�
����ޡ�7a?���o���ţ� �7v*�Z9O��W�c��h�3�����11_�\��ўO%��j#-!�Q,i�U��}���X��(����U����]���ƕ�9jw����1<��M��&#��Jf��I߾���)�Kol�N��+�s� 3��:��kg�˟��`r�ڥ�����Q�R��l�I~m��vq?G�G�������۷���:1PO�������8ś��@����C�����C��D���+S-���ч�:��X�!؂�E���M��������y�?�	F�~Fk�:�<�� ���Y�W�p
Ꞽ��͛] ��	�OZ�j��B3B��M0�Ha�o0�1����� Ѓ0)��жo���7i�$
������=�~��x:^���:û����q��-[�� Trsr�+$�}Ȑ!�"��&0:G����W�뮀�o��棏?.6��
#78�-�i����}1�@4¨��>�����4��3^�T���q{f
�<�g9�1���@K��h��\h����0X��T^D����[yzy�����)�۝�v^M��ח�\�)��U�Rř��S��x3σD�
�k�y�<%ƕ���������=|���xY<1�j�M�7�Tk,q����1vի9���x��	�A}�bm���׳g���۰���!�b���ǏS�R���WB����5��C�>������D����J�
�Ӛո�8�&**�>�##6lX���W5a��]��9�˭;�˔-��؏?�*C�=���ݻ7�%oe�`����mȈw�؟�3�1�{��rP�?0��/��x�n]�����)�Z����p���t@�e���g�J8+�'pe�Ƥ���4bG1�3����@�i]�b(9��p~��}�˫�A���j׮�S�P�
BnѺ7F�Wi�_Ƀ�,)E�ͅ7b%��=�D���pK�����������b�Y���x�܇6h��@�L�z�0(>^x��wg�b`�����g&�a�)��w�(�T�V�������5��>7������������r�*��0s+	����B!���Z-�,`̑O8�虞���⥵�񒮾����{w���A���}!��0-EZ��*M�A�/�@����Mh��+̾��V܄�V-�8�_ }J�n��JwՄ��D�r&��he�4z�X؀jV"%00�o(��O�@�PtJ��͡1apÈܸq���ۡ���&��@{��Y�f�܇q ����ʕ��d���J������Lx.���O>9{�L��Ç�R'Լr��ԩSѤ�mۂQAM�0�A��0>�	�L�Yx�\��֨QK��n0�R@kC����v�4���,�B�IDk��nf��޼i�d�:u@�Ν;��52*�R�k�c̆f��)Y��y��tf��ҟx����b9��Al��0YyV�jQ�����KՃhi���)��|f��l�AB+8�_�@�y��@|m>�Dx�ߢ��[�����="�`ƟĻ��<�U⎢��x��#�qE~R�+�'�<�vF��Di�p�]|O��סC��pg�w'�񒣔̘V���4B���5�iӦ�!�m���Z77�Q`H%�`��C��S�B_	��^,�n�F�_�W��c�2L.\H�֮];��Q ?�����cb�B��ݰ��?��AbbHH��5����߉��V���o�Q`�G��z��|�z�ֱh�0�ٳ�.Ġc�`�b�Q�2��l]+�%� �=*�+FXA�i�L,vŌ~�J��R�+��F��}���giK�N_�eZ����7���t��g���Г��j��7:�~���pNcR����)GlذaȔɦ��]��u�������'�{WT	w����ѣ�舝;6F�o���%�6���\fl?�կM�}�H�u��]��իI�SAic[F�:s6�R�""BЛ.�����/�8Vy�=q�dn*���a����k:�'<�������z�Rc������o��UZ���8��R�Y������,u��	����Ʒ�1�	:]�$y��Ka�xz9#q�V-���U���{�W�.�ӵ�)���>�a3��@~��� �ЧPs?��Ppƌb0����'$$PNL�'�=@/�[!7���L�G=r��?f㡰�A5d��PaW��V��rv ����ҥK�v.^$�x��}�X��^� �`6Ԋ60K�������v���s�V�X�V�Z�(���J��} �p��A|ݻw�SD~�;Sn|(��>�h�֭̿�'�&Ň7%a�/ Ӗ�����g�?$����-[��Z�v-���2e
�1��(�0	 W������C�
{����n@�sg�^�t	<��]�`��7�$�G|
�:v���'޽�)F.��z}���q��ߓ���5��s�9�pA����z���i�e������V��áѺR�Bm�@.�����P��^��y�&�	RA��h����D�w����_�ś�)�r��b��L/#W��Uȉ����.�����?���/&�ލlk�3�.���cB�A����9�����CƆª��rGm3LU\s��=�?�;�S�޾};,,����]�t�y�&�6����ʊ���9U�TAk� ��=(n�ꬺ:Y3R�ͳ%z��\���0ti��_F^B��ܭ�MN�hl �TF/.��4&�;��MKMe����T�����ϣ[�����.����ݼx1�Y.�Z���ITe=4E��5���Q!��,���v41Ie�Z)���>B��"j�Jc�[y��f���`Dzyz?y��ﾃXW�\�k׮�?\��^(v��T¾?X����z19_D�t(�@qk�H�k��tO�D��]Yz cP���\,��Jr��K�f�Zݵk׆�ܥK�-��EsGJr2�Ftt�\R��gϞ�ׯ�ģa��I�q��a+�� [��v����a����\�h(��̩��N���e˖͛7/�\��'O9b�̯�3v,	�HqyhJ111�W�~��F��rQ���;v�~���C<��o��߿��\�r���\(5gܳ�'��Y�~}�;�(�ʕ+	�ܿ�hѢʕ+�«�'�+�����#P�:u�Pns�υ����,�&�NװaCH8�����q=�W��cG۶�O�<^��ϡ1��ŋ7V���##��8�����;>>>᫯�8q��f�):���ed {���e��V#�]7n�M��(w$:d�3 ���8}�t�1�e\6�E�������G�;:�U���d�@���H
�teY0�Iv��Kw�sA_K�.�bD�T��W���#vv��<��4%� Y����(y_�禰NA	�b�fHH�P⠽jL-i�{�Er#�/�bg���,����Z`^;�\�ʢ�Bү����cǠ^h���|Zf� E�#�� -�$�@���]�j֬	��~�:�����9s�R�����^Q��b:�u��<=~������q�Wڕ�8�����Q�T��ڬM�ۂU&�m������YYz/���q7�' `��C�Ӧ����JՄ�ǎE׎���)�m�vS��&�XU6�ʻB�G�[e˖=�}&��r3�]�zz'�|�Y#��xV$�W��Q ��:��2�JPf�<��IP�B�s�K�Z�D��_������>�����j<|���#^}�7SyΨ���x���R��0,�5�4�!�[E%C�!�F�B�D���}�vf�϶x��+6,<�9EZ�}�E�Qf=�yد�;w.X�s���hk7�	����9g>x@������(,��СC������S��ј��)����ў~������.KQ;k��{���8p
�y�_сq��\�u�6J�Ү];������� ���U ����7`� ��{��ay��0�N��E�K0w��`(�;v˖-�/F�7n���������Dc���^��2�<}��k��A@�����t��S�N}7o��d�kX���3l}<(#�)�7���s炸���/�����Ve��_c��͝���ۅ����P�������tZ-�	ހ�`N�LV�h��: ������އ�-_�����T�Ũ͙3����=O����z�A'_�p��!���cLm����Ђ���k�{�̧0�4^���X���Y+�[x5�\AWa��`T�Xw�P�ֻ܋}E�/���[��N=�P�jc�jR�U71�OD��Y�J�+�;�N���5��=�)>�%����~�_)j��n�Թ��c�����Ϡ�`ކ�բ��/�L�0D�� :�gz &��J~�$44�
�VK��7o�H%hK�I(��@�b��< ���Pb ���"��6���l=���)�?v8^h��)� �II��w^�ּ��S ������Q�)_̻vj�l�xIPJ
fx�-��OS�J�P�TϠU��2&��w�*�zeWJDƜ!OL46+�<ɔ���UQ�;�'/O(=k2�@Z��E	K�VL�:������DO�G3��"k9���>:fߺu�Xi)�8Cb
�Z⌢��@�!�
�C:���C���S���QɁP����b,=�W�du�*�K����t+U��͈G����7h;�S�ॼ%�۔�'�RS�DAR��~ҝ��}Q\�|.�v�@�dV�E��>��R.8�б��;�+�%�G������T!l���oLV�c�� �ڷo�_x~7��,���G���^��R���T א)�
&�f�)kK�/۞gG[�oY�30�ȱG_������0eʕ/S��ٳK�.-�E|���	��.�$�|y��x4f�������wd H۶mkԨ�J�޽a��&�������G��ջs�.��ٳg6�Y���}	�ݺukZ�%B���nu�M��P4{ҤI0��%K�Pסߢ˕�?�/Y��"�_�`AJJ�� 
�?���jCS�+Ww�ںe��|R(oݺ��䂍^�Z5��Nb��q���݉F�"�q�8q�Ĺs��PP���)��ʕ+?���Ż#F��cǲeK@q��M�4���w��m���o����i�
,600̣G�֯_?{��:���HI��Z� N%T�\.w������=^��	�F��Ķ�K�W�V��+K3Љ�۸�fYBB�=�l�C'0j��V�Z�f�J�~��ШYt>N�[XN'�*Ϫ[yx���k׾��{$�W)������sOK��\m��� ��G3�R+V	�xa\bFk+DE�q����6?���'z����"Ur��U��+�5)�[��r�1æ����*����AmyffT��2�F���[o��,Y�aPjԭ��k�ܿ;��2Z���׫�c��5��E0h�:�IbcV��X��G����l۴�[.�M��?΃ƩP�B9�ۥ_~|lW|B!!A�4����4�6�!�
l*_��o�odkz��2�]��
��E?�h�ǩj%~>|�S?� ��h���)܋�9�Ρ\��p�7��*��1��6 m�5�r�����b��,�Y\�5�;��h���l{&p�sLBX*����KCu����Rb��GY M&����2�_!�'�R<�`C�ёi�G��� JKL��N��P8����!.K�֐i�_���Xe3��O�,W��F)��'��8Q��OtA|.�F:ae#Ξ� �L�aNR%^L���|�VȜ-��I�>}1%�j��q������b���r�Q(���x�T6)�����[�@�Ӊ��S�Ӻ3C4���/�D�sr�|���qq���d�\�04/��g��5Z�W1�ո�f��=�_���U�9A0`��j֩��o	U�
������O��٬�~aTyq�B��ۭ~~���u���)��ђ�e˂%ԭ[_�޽;��dCC����=`�;��L� �Ç����ڻw�?�h��+��R*U��`��?Ew�ԥJ��M�6���dɘ��zg�1ߨѩ3��9�ĉ���KE'I��n�fc��ͭ�d��m��ԩ���o��_�ӚK��5�����wG�߳w�M?�����s'������|�����U)?�:�ʥs_�5���o4lP?�Iϝ�"�Ռ��KB��W�q�<�(m��y}	�ި��YIxÌ+vHKiOd՛�ʟ\�D�'Č�8���ҽ]:v7a\�~�`��ICHBC��.��{��G���V�vm@>��/)�ѩ�'�l>0]贄�J��*N���<M�9*�K�eQ/�I�W�[����g����9ݛ�7���_`e	
��}��p�͛�����OmB�獤�) [k⏷�����zp��b�FVHM�������X��S �*ˀ�� ��Y�^�����@(w�t�U�Q#H%'4<B��C����\���$�}c!\�o�%�0��k]3�R��&�I�K\S�t�wOOK���E������V�	�쌗i��U�a�H������ŏ?�S��d�6�D��jK������3
�4S�	��䳄_���)i,�,K�S`�	(�ND�$##�. /?�R�H�:P*M����\�-��_1�q=ݐ�"�!��Z��m:x�v
��K*���z~��bU�T*�XC�
8��шJ',)����B��Gh��ܑ���s��x=�Z NDeh�O\�Q���Ii�pB~�;w��-%�'z,�:�*�3�~ݶXNn��%���6��ĉ4�U�V-����PH���w��J�@6 ���]Q���׫W�W_�Me	� X�[�nmب����.�]_��v�|�r���t�g�;w�}�����$��|󍇇{�v��l�taFGDD�[���0kL�j���}��߿��ɓ@���W�:���B�))_Zg�Eƫ݊�I��<��A�^��p�nb���w�ܺF�jkV��z���b;w��ʕ+���탇�{�֬�3�+ܥ�N�:����<O�0�vEcM��X�߃�,|Y�u���v�:1r��r����v�F�x�\�z�ڵkO�SZh;�\)�ý{�(c;JLqU��|�_�kx?�y��ڵkPJFc>&rI��b��+�/A��ȋB�?�
��Nzm������ K�7<�I��y{ɜ����y�]�x�
��9������lYU�g�as�w�1O[�7����sAA�'o
�C.�`��P�݁p9O��{��Ļ�n�������*�� �+ol�ȋ��1cnܸq���%ᨬ0	� �s-�-�p��(����?��R�C,%^Z�]Z���WM����E�@�8�����/KX���
"
����h�B"I�'r��f�e�,���H9�E�b��t����H9h��K����T��)`Y�2�V�V-2*�����b�7o�{zy{7m���_mݪ�b �*U��t���x��+���!dc�ԩU�V�����d�h�ziUu@��A�U*�С�~��-Z@���+�8.��D��F��0 ���˗)oOeM�G�jի^�
������;�Ao�Ix�5j���G����|X��>˖-�����xL[�Jm�Y��38˔�����"�݈j�����cv���))�˗g�Z��32&Z&4�M�6#F��ݻ��'����0L�����/))i�̙`],iߘ<�=O��$z��A��?u��g˟�i���Q��Y6��	{��A��"M������!����T I����4l������rԗ��Y xJ�U�Qcm�f�?�Cd����0�Ba9�g����V�O\-Fw��P��juxDf]x���g"�6Q�CC��=`�����?�y�2����)�%gP3�1���ͮ�T<G�ф��VIo�='NF���\o��<�3W�5 �rN?��m܋
���7ߔ�eP^��Dq�'�'�(^��#�8�_w�y�O��XW�B>��Z��6�V08��iz�9��ލ�+�
��YY�`D���;�װ����l�t���5����ʙ1����yb��%T�
\���7޽{��'�@Rׯ_I8�&T�͛7cbbϰ� @h���Ii ~�&_�˜�G�_��cǎǏ_�t)+^�U�a�({�=���$Z�i#��l��J��<x�S�vЕ+V����X�"{��������-�q����hH�O?�T����c���d�#�y��C�+U�����6h�`������"��s``5aU����d���������%��r�,߀�;P֬Y={����`�;����������aЃOpǣ�O�Ҁm�ϙ��&$B����y.-����U� ��]�reƌ>�^��Ų���c�x1$�mL�P��!e�	��l�&�mM\ �':t(���[7n��>~��70��ڌ�u��U|�B (���ݕ�$�����L|N5?YQ(�=��#44�H�����LI�>J�����)�G!�qz�_=�v�zA%e��>N[�>װV��l		���5^���q�6��ܙe�aq�V��@L�Xh%�-9��_��5'G�*I�l�W�`FI,�m���xfHY���3��5YH�U�>~�Bٲ2�Sc��UJ�"=�w�t�:w�|�)�qwZ���s��(,�]�vISŉ�����(���C�dh= �g1�SQ�b�k�Z��rq�@l���D=�?�?IOx���׬ٻw����y���]y�r5���~�՝�!�NzU���I�(i-`�,�w�d}������?�?%,
��K��s�l��Tq�G�$��E&{��	:�r�S�2�13>��PLcXٲb�8�+R�Zؤ���8�]��$E�0������g�ʆ�O��q�u�֓'O:t�7�⚝�t�ܹ3�����-��#� o@;��3Ǐ��wq�z�"B�կ\�"�J��Ӝ���-S�m`�,���"���O�ܺm�#G���9��^#)�4i�l�X4n<w����x���ի����==q�60z�����bרQ0F6������5"b�� Y���wB��m��@ES4]\��III}��E^�|H�N�|���ׯ���@n�����_�p!++��ܳ��o�����)))��D#���\�,yQl,��"'#���6^��Oq�b}H�&9˅E�++��,�`0<.�w�P��'����y`H$��l��pI�/�� `��� `�#LŮ���txrw�R��i]�.�9�W@ �-%���Ο&S�Ō��J��b\
�/���ԮA�����cn�B>P^�f͚�?p�B{��ȥ���Ǜ2�A)�N�si���ZU�*��:�ĥD�yo�|5��'�(��Ν������k׮��%ײe��>���U�Vdx�1?���'���v�����µBQ��z~��筃���Z�kw��#�����W^ ����Q,U�R����.���K�@8xB@�z�<���A� }�J;�χ@��8�tE��qOo�)�2ݍrxkX+��G���N���?P���=�1�=����'W3�V�����x:X���ć�LUzD�Sb�|7 00 ���*?�6_<�ծ��,�����������~�l�+��+��y8 L|B�7�|c��cx��{�XT�N���Or�3�d������;��~��irrr�T�v�;w�@�^��c�ʕ�5�jӦ�
*�^=<���_Ϟ� 1qӦM�:u:}�4��О��(�^��bŊ-Z�gd޻w��`cࡋ-3#gg<�����X�w*�ִiS�BQ�Ic�޽[�.�!)꓿3f�F�_�3NE�6���,��78�L�J^�\�}v���Ri1�ul����B(u����:���~� ��y0�����ޡ�
?�I�#�u2�xT�hi7K&�F�
����빑:�T���r!+`Æ����]�r�8-p8`^��~�����˗/�L=f���8�x��2e��l���e�h�"����P�"���dh޼��y����TT6Lz
3��a�[>-�Bo���6i�D�CB�V�\��o�Θ!PR�\:�V�v\k	P��IL�����.ߙRmY���4#ҥ��|)<���������_}</�;^�\׈����WМ9s7؝ ��g�������[Rw�@6����
ܲ��a,?z��},��]�~Qp奡rv�{�ޱc��b�!sp!�����}L���s��ip�V`2W�~.�P����Un�W|N��� �9S�|��k�J��v�k*n��_���VA+�m����@�B�86�#�TJ����U!�)��nh���t�JQ?;���r�^o�����Er�E��>.���;J����]�VY�l�֭�T�z��ao?_����͛��{��Z��|����wb��#G�ԩS�u뗞=˼y�vDD����i4�gd�<NIݱk���,�C�0[mF�EpEEFǖ�S�A���Ν?�q�=qℏ��wOLL��C�P��<�4~�~� � �+�S�565J�H���Uy�J��n���ye�>}�O�>��@�}~�(y����������HI� N$ӇT��˫xL�)߬Ֆb��A�>�3x\�y{yz�Y��Km�
|ؤ��5�"��Kl)�l�=�D��T+�\��p��?�
h͚5ǎ�V�^��C�u	�+W���x�lذa � �1Vkrrj�rQ?��S�Z� R}��ٵkW�ƍ��ƍ;z��`�oݺ�ڵ0�(
2,,���OL�6����_;v�E�	0d�1�� ZrÆ`<8'�ذaÝ��ԬY��4��>t+��;Q��̌�={��ujժ>N����OnݺzN�^�n�x��^_,t�����ٹ�s]�Čμ�] ~e�_!e�u��k/��d/Q�޽P��w贜�<�Ê��@ �!!!�}�9�8{��!�1�Cxx8:�Lh(���2�s]��Y���Z�j�xv����a�Z�C ʏ�Owo$�ȷ�����W4<UY��E$����p�v�O���A����G�C-�|n�1*ϙ-.3��^�[I2J�>���U^��Ee��8���
:�IV�H o7�����j��Z]�c>UZ-[��c��r�*۬�mp�C��?u_��Q�"BB���0` �4���ŋ��̓|�۷���0|���ƍ�+gϞ%�}饗 ����III��ၑ���r8(�K׮�"��cĈ�Fz��A�+�&=���0��R	�!f-v��#Hƈ|l1����Ŋ�/�yJ�4a�>>��G����r����d�Ւ�u��}j��2q
(��bӹ�%�f�J��@�����M$EE'�ͱ����;�Jn�Ye%K)�� d�{��5��|�G�c]c����ꫯnݶ͙~���ӦyށrB��VN�5`v�[��+�xu� �a��?�}���<#�UL`��*��������ھk�l�B� ��ݭww)^$�k���RJ)��N�@��{־g�����������䷹�{�ș�<g��9nnV�,׼��g̘�ײE�;w�ܼy6:y@�A��(�� ٨!^"r���|X0�.��v�Z����<`����H���!/\3�͒^��.]�<x� H@j��Jb.��%\�|1�re���/���P�Q�s�����P�S�LY�x)u��Gi[�l�ؘ��ݻ��T�9�gO�:��ɡ����aC��Y�VoЋ��}�����b\������ �s=#�"�h���p�G'�'ak2��쁾E�l�x�
p�o�-[��_����,[��E��y�)W�6w��CAW�Z$��3oiӦM*?W9|�p�F�{��۷��@��ܹ�y�,�?����\����0�0�fϙ3�|0�}���<qb̘1۷o�0a8%�h��ݧN�Z�l��Æ bbb�*��������>�6mFLt��i�V�X!�ԋ7�_�����_}4څ�4l�b���ŋ�~�iРA�rg�?w�*S�ti\�C�z2�/�x+PR��m�@��pC��i��f=>��߿��	`�E����bI7:�L�LNH���B��6�H��,<p�xLF�$	�WC$0�.\(7���M��&�]$�@����.�۫W/ ��*��رR�Ni��dڧ7��ߢ�d{+bb�^��-+T��cP�n݊��"* =�х����� �W&G��u���ꃜ�Y��D0 Pҙt@�:�< �w�>�'éS�h�|�v��?��R������={R�Ġd��M�ev��*b�8�j�ӧfлw�
,hm�@=Jq���?e�B!�+���c�x����65`��"""ʔ�����|��4`>V���Z�x��3::���畕B�K```��ͪT�|���"��!��A}î�߯ߏ6 �(Ǝ�������ŋ�i�A{��OOo��-� DYeZ���j9f惃�T!f/�y���(� D߅��8<��	� ӿj�j0�.Y]����}�A4(�-��9^����f�\�dI:���p�Q�k�λw@#8>�;�`�� ! G�ر#P���?�RQ�5���͛�;
-ߦuk���ɉ���_�&M0��L<��g�n Ǝ��.��
*�m�P�iӦ!!����Æ#�f��\��"��c��cӰaC��'��ƫs�N�W�Y�f;w� }�Iz:pt����ڵ�7o�G^A�v�ܹj�*��# ��� ����oÆx;�!�_�6(���}���+ �{����5a+EG`^L�4	�3f�\��ۛ�E�9u@�5<�z۶mA[��`rw�<�d�����"E��hB�{�˷�A��>�π��������ǆ?͛�� l����Q񖨨��-[�l�<99y��͛7����|�Q��/?��1(Q�ĉ'����5j�+�g���ؗ/_�,Y:~w��G�  1��z���x{�ߌ;v�1x����###��޿[�d�5�el,X�{�Fci	"ȏ�U@�%88x���h��{6?~�ݢE���8z�Hhh(T�H�P[Lp4��w�<�r��U�����!Օ߼~�A	�O��'F5��xfeZ�� `�;�B���2��AM�W�c��|�
RײU+�\�O�<�4%�̤Daޕ#��ׯ_w��O�+X�!D�At���(L|��2I��tfU���,Ǖ�t~�H$�իW0�M�Dj5�2���x`|�.�m��3e����7�E���G�y�U����b/�O!4���L��(� �e�2�6��s��W�>}0&����Mjj��haeM1��'����۳g,	R����4z�`��#c�R��CڗlL9�'��3�ֶ!�����mē'OB^��#9�� �ŋ��5ܿO�^����,�y������/`�O�8	x#�c��:�L����g�A߸A}�o��C��,S�B���'�N��Pܿs��	�寐��g����LM��V��P�s	�)�I֖K�,'>O�*���d�˔a��ǂ��I\�x1f >��i�Q��ց�������r,V��T�sX�!.\��e˖ѣG[iX��[�VM��9s�D���,�F��3��)�?�:k����g�<~���6n�(+[��ŋ%�'޸z���/����$WW|�⹳�N�5�U��Y�p��S'q�jw��y�v��?>&�� ��֬\ѩ}���w���Ջ�5+W�mۮr�*v�6;�n�����ѣ���q��dM�"u�0��+ ?�aK�Lޘ��!�B�.d��a. ����^�x�ǵk���ƍ۹u˷ݻ�U"�qd׮]QQ1�~�d�E��CyT��G�D s �P��<1��>;�ΗR��0��Ļ(��y��,0t����-�������s���N�aJ��؆9U��ͯ��>|�����**Z��C��Idm�U�@�ڵQ��7��ז�*| X0��@�����5��A`�<s��ojլ��ٳr��-^�x��aA�:�~��11Qj��ǵ�:t� h���)����h,.��P��`��u�-k׭C�Μ9�}ąKٕ0�0=Q��m�hT,�ް�#)P&_�f[����;����V.\x�����7JOI�7p��}?�΢��Ν{����=y�֥+�&�@�����={r���#G����/��ڵ�!3�_�^=�T}��Ƹ���cg͚YlX�ޛ7op?���m�2R�;�m��R�R$�m���<
�	�����[�n�hb�t�����ˀ7p�:���h,Ӓ��JE�4��|}0j���-`���6�ٻk'�C�vmw�#Bl ����V���@e:t��$6+7g�*	n�΄�C�B�@���d�\�lp���B��8^HP!��`L(�O/������d�R`��~^>��9��PPdvΐ���y���h�_���
�R�+1�������im��{ ��G�`�ݼ~�}�����L�B[�sp�N�����-�
֝F!<,�|������	4�2�=�V�����\�^=� [^��}�{��ϙ;��"�l�#�<��_<S���'MLc�b�J��?t�p�m��� �f>>�6�So����r��خ<���]+GG�۷nAK/^v�C�Z��cg�0
�{ya
���쀙�*���P�ջ�4��3�%l�3;t� ]`�LC��@�CO�?)<�O�*U�^��e�f�QAD\]�(�@zz	����[�,��8aT��8qȐ!���LNN%ȏ���V�nFBdrg�K���,���=̩I�&�,>�:D��+U���٘=�?�:7w�@(P 35)���4�BZr���,�5̣v܍t߾}+W���D����g�B:vl�o�/����"�k��o��1b�":鄱��@�Ё��	�mgo5
E	�v�e�beg��� x^|������/6nX�s�N-�H��--�������K��U�ޠ#G�,W�����s�F�Q�|��:���G��>>~���
�G�8�a)�9�!7~z/�4*o����hѴ)���ի�,-����%% N`��C�E|}QՖ-[��ؠ�$z�V�0Fϟ?$�ޣGxXXb"c �v�7�1dh#�Cd��瞧�b			A�0�##�߽{��?|�p��mڴ���������M[��Y	 N�� R�>{�(���w��0�PN��Z�nݶm�⍠Ԩ� @���Y�����bc1�N�9?i�8���M��U�7o�1�r��և�%�z�ʕ�̳g��*W�l�WY���H�`7���Q�n��ŋ������]�ft,XE�
�...����S�O��¯&�N
;u��CT��}�����r��$�:�u���Nf:����+��+�VZ�L
"����<P&y�Qhp�ܜ�D�-����#�<Ԓ�/��v�^Կr�
�����X�-�4$���
����a�V��H�F�<�iE����Ws�VKeDx$��;�ݺM��ʔ*������21	�9=?�͟@�����=��O�MFr��+��b�ٿq��W�^�������=ƕA�N�X�׏�7�SS�\r�3�4�Uy(�+|a?��&^�v�\\0UXԪ���ӦU�\yРAϟ���i$�}���"?��<�	���-[��42�Ew6!{� ��i�
]ଂV�<��&�h����C���[��FMM-W���c4G�Y�AR+Y���'K�=�33YY��P�:�W-�Ժ��FN��|�B�t�Ȣ�����,��l.���`�?� �ԥK�S�N	\���VMzJ
~�Z`ժ�Lqe|,F��{�^v�P�y����|���(��H=^�ݺ���vϗ���A>w"rq/0pz�i�<�J�@���7o��	�z���{�RT��0��ÿy���>�d.H�.���q5~�f}�re`�W`!�R�n��ÇM�0@��ր@�� |}����M�P��?�8Z�d�R���mH�P�L���B��y�^�z�T��ν{���p���Q+�u��y?�P��,�/��8FDRHcF�	)	��|�O�ޤy�x_]Fz ��'��$)!����-%)�Bc���-���..�8K�.E��nߡ�/���H�Q>bj[�;�V
Q4Rl8~&����j�>P�1�	��N������(Y�$
*1�T<l�_T�L����+����� ^[�`A�OΕ$*	�R�\�Z5k��d�ʟ_�T�'';9ضi�f}!�cRs3��twu�l΁F,�Lֽ{w4����[�nE����#N��)2"�XѢC��PJC߼�)X�d�qgη��\���޵kA��ܿ^�bŬ� Wg�ciJ��IJ�r�l-��dX�-������<�k	q���bY:`�q���m�e)F�+�G�����o��bZ�
�N����������1��S�^@�i��@���p�*���H939D���޽{�-^�~���!��޹�)�����*�	���hegGk-���/)Ϟ=�0�9 ��G�
t>PӠ+4dK��f笈�(2 ���A*�Zu��U/\�
��`�U%�`l4/�jc\^�#ȗ����-:�):�[�H�<���_/g��T��g�!,B�^Og���I��0:�Ű�6��-
原�z'G�Ǐ��Y�|9���l%@_�xTχ,A�@�Ox{B���5���T�������0��j�1-$ �W�Z5{{�*0��M�σ��Ȑ@��|�Pm+ѽ�`HHL!&�:��@"E8|�0̸�ްG�M>�y��z��X�+���d����ӧ-�pޮ}��ׯb*B�@��D�۵kנAT����`��$�˗/�����7@�p��ќ��تU�>�\��	�5Z�vUfݺU�X�@�Y�r%�,>.4�ߥ�:u�4kֈ�NAw�ih+�b
���ʘh���F����fժUm۵�U�֭[�v�ܩT��t�̙;��.CgB� W�6��`ܜ��@dd4l������'�R�B ���Λ7oҤIO7 a&˞)
K����0����Y�R%w�AA�'M
([��`�b0��G�Z��x�pU�!�Y��E3�����Ν;0�i�����̓���ș��CÆC���A�q���o|<[�#�w�"**�A.���3g�o����F��:��F#��B0�soY�Z��"Ņ{
(��@�i������4��$��PO6���	l*}i����"Nj��>��(���#r��ȃ_I1�����><��'���5�x�Y�|�	�(��#�B�I\�e씞������(�����Jܬm��V�T11��L���D@��/v���,�	j]�`H�K��M}L}���6�P댂6�ݛ]�vmް�ŋpg;�7K$%$��i������L��c�a9�^>�QCnŅs oke�c�3z�֣�AN@�e�R�Za�g��
�ש_�c���Ν�p`̠Q+M�=E0 ��T)W�̞={`y���@Aet��I�v1T��@�ðl��Q��<"����0[
�X�O�Q�DVAJ�N�|�P�GGH��C�3�OP@�Vj�Fͅ'�<}Z�X1tBRrl''�.' ��0|�l�r��]�-�+��Se���cKD��G`�'O��o�~5�AT`,z{{�����Vǎ-ZE��W�&a#�W1�/]�~��Ih.j��>�/�J�vA �㢣]\�Im�-)z?^�����]Ֆ�.]BA�����������9
�;�����'&$8p\ܖ7ovbhhMV/,P�����b���3��q�gϞ���aEceE�0�6jD�w!��� �RS�@1�(gR׮]AV0;������G��^�����:|X�����p�B:# DK=z�H9�	���4nx���{��_�>?)h ����p�)`����`�aPP��F?�Z�n�� �64n�X�ȧO��ׯ_��}?����S��+V���32�䰰���_��:t�w�ޓ'O�ի�L�u�D@z�\��`��o��ZP�B+�ё6X��c@llT�>���毿�j
�X:VN�a�RYn�(>�رc��"��c)՘態�O4�*T������M�*T���t��F�D<���3����a�k�n͚z��)�4�3�|���"L^(�@JcA)��_�C������ڂ��~�TnR&YJ:*�s��sPʗ!�p���Q��O><�QHN�����_2�����M�V�Ǉ����!rN��Z���/
�v���y��;�ׯ�����S�Nݽ{����B�A u�w`6}j*K�����RS���]J����R�'���!V ������J%>�vX�b6+�-[6x�`������,v��۷aF���D���3z��aòn�ή9����fϞS�*C��P��s�͍Ά}H�`�A��av����0ㄎs���>I�Y �Al�[��7�����}߾}��;��ƌ�w͘1w�-[���3�/��[�P�BP��._�8�~�@�x��b����AD��k���#ǌ�i�x�����j0����S��w���VA��؁�;��m�62�(�0U����L����Olw�`pqwG��4ή�u#Z����O��	 ��HMM����BY��"�8��x�XKq�h���PIP<1~�x�����G���X�4z>mM��ݘo��г�Ή��L�mtvq��ķؔ�K�^Z	 7u�3������j���������%���S�����99�<�`��۠��bG��(ڍb;��P't��M�?
�Š��]f�����1�s���U�j�y��+޹��Ճ!7��;u���/Ybx.Q��`*䞲x�b�]�v�R� � �|�
�֭[T�ɓ'�J x��ժ]�M�cF�d�iÜ�\==W�^M��^^^P)�d�L�~ԨQ��4ǭ̏Ȃ�8�d��P#իW��󵱁f`lC&�_�!@}����
.�`$�Y�R�A�A��K�23�S� � ����QQQYiV_�,��Q�9&O&�%�������|}�Q�NB9w��m��Y�	��z���2yE�&�A5tȨ���/������_��^�z��&�L���u2A�Yf-�s2S%�Y�)��zFZ�Ik:>+�;7���ѣ҅����%D�X���9�GF�EFE)�*�/8x�
��=��MLL���O��Xԧ��mC�7~d�)=#U����L�|8Dv���9���-��[����e*>x򜉔y�M|�{�1ag@��E2���i��+b� .]��d�r\i٢U���M��r�J�
��]��9�{�k�κu�zH2�h�l��"I��Ng��~�Ɏ�#�	T�2��88�4(.)�����_�ܚ��Ǐ���0bĈ�&�����S'z��������s�H^,P"'Μutu���OL7���n(T����[��5� V3f�]2���7�1���E����BŊ�x�gX��*T��4h����J�7��L��j��F���?C�ֆy�g�������ݼ}4>�y����#+V,kѢ�0����k�-��z��(]�����C�Ӓ8���@����ؘ��|��'&$�+,�ʴ�d��-����^0��MFp����|<��A�6S���)J��q&�3�:-��2Y�S�:��R����
%��K=@D(a���O#s�a��O�? f�j3@b)U`��Ɗ��Z�b�`!�,
P;

4���Uj���Q�t:���T��_4A>���R�0�����h����W\<��WkG��]����h�ZmiRbj'w���V��Yʃ��MN vNY<�K����'�$�i����?���b��e~ۓ�y�������+V��<2��6yд	�ܐɼ�˖�|�=�(ȏ�y�jx���8j�$�'�]��t�R���ջp�[��T�]ҷ}��ܫ�Ao�Y�?{��M��ITV?g�3�����t����/����T
��Y�L��*2�^����� �:�Q�$��&�1�J���Q9�Z`���`R��[�Ed��ɤӂ���֒��V�gB�|�t��v0E�^��F&�*�Y�Ef}�B�� �K��_�p$�2��ؾa�}�
�z��ٸqc����4�����$x6����#"z|�	��ƣɂ�&�}8X�"��v:~��D��90�������h&l)��gV=)f�9��'���t頥6t �J=�u?�N�e���g�~Ȭ�2|��	���ܳg�ŋa�رc�޽��v��9;;߻w�`�B��p;���J�N�"���]�hٲ%y�R2�A����y��n��
B���ag`�
��ʳm�K�.����9�X\]]a�㱰������c��c�7�2��ϟ�r�
;�٧�`>$���`i����B�K�5<<�Ν;>��	v��qt):�eȐ!1V��o���A� �dC�8q�����7S�r/�#�����ӧ��	&lܸ-�y��i�j֪e��k͚5+Vİ�=�t����~~�>�I�)8����6m�8��ff���� �c����\�:e�X�x&�}Ll�\ㆍ:t�اGO<y�ʕl	�l�:x�e�V�5)!aժUcǎ�HX����v���+W����a�G��CAP� TDRR��9X��{P�Y�=�:(۳�x|F#��P�t���2��#�V�SR�)�(�6 ��Uѯz�h:��!P:1���DE�!�Dn��W�7��̱�0�t�d���IN�JHZ�<�k+�����?�ia"vJ��#۱\?7އ�!IW�E)�����]�~�X�b�c��D}顅z�N7��{�.[�}���&XX�>��}Ȑ(�J����Qq�q٤E
��U��T���.\x��Yo/O�*���䤐�����F�ö�����a^�0�{{�����(��NnO��q���8R���TУr�o��������+<ܫc�6ӦM�ׯ���Ӷ��s���C����_��.]� ch�Bw@!�L�tZ�\�@����y'ђ ۸�Co�)�H��e�f=F^�b�H|͓>p�,!_0�ސ�`���y�+�}�ș����:�!�V�zu03�y���\�vm�R�
��?���`X�X��n�z�֭���G��n�g� ___vn�hD�ԬY��%�&W(�̞M9棣��xt�v�Z�)]�B�;vt@@��ի��%K)Z��*���w!Er(7<*���3-#:�����ѣa����q���T����ӧŋ��ڵ3(���E��ׯ_�D�?�������6l*��ݻ֭[3��׷i�� J��  w�pΰial=|� ��)[v��q�:,!�D�qW��3g޿<&,,�����L��IND���?�bٸFN�ȢP*�"��tbJ�Afб�)�8}�&*[S��/� z�7��s9eT�:O|�f��h

9�y2�Lω}�^!�.��C߆�Z[at�*��K�� ����++W7��ζZ�}�X��@3��ܔ�!�Ӹ7O3��r!�l"��}ȥ:G�����/��!x=�zY�H�FGb;w�<i�$���� ��OaȊfj�I~�E���a�⥯^�+R�o��	m۶�3��Mg�j���)����#5y��bR�q�M.�A��gu>T�p��M'�8�z����s��E���_;t� �8�[�aC#""�={F�lٲeɒ%P�...��]�T'Pt#����	����
��`v��'��yҋ����K���c�,�G����@��	�4ַ��]�����nkt��
�BxD�c�[ƔJ,R����G1!�ByF��p �_��~�-4Tݺu)b�ʕ�����Ա�g˖� W�]0��+W�x�ѪU���L�yH���۟<6�|n���ʿ~�zܸqM5Q�;w�_�	�b'N' ����q�:��͛��|G !�6�#������������K�L֭[�۷o?|��	I���/_�\�b�]�0��v�W�:���7o܀l_�zOF?�޼ys��%4�|Mr��D�� �@ڄ�a&�[Ze�jӵ�\��s���O�A������Dlll*O�da���])�&}+��'R��c�3u!g�|�^��i�\�2o��>��������c5(�������F�$��ݻ7<<T8-!������R�[k+K�'%9?[4m�k^�L��<s持�Fs���)xI�� �$�:�(�Ղ8�)S:s����T�m}�+$��~h"��czf�wĨ�C��	2�+kkg�#��)emF�������۶m�Hhzw7�^��������P��h)���f��I�T�X�"E�,\�0((��f�1��c�?�
�	Z��$��`�өzz	�\f��Z��E��P҉�仛��k�9BF��p\���{ѢE ����br^�~6����K��{��	WΜ=;{�쨘�bE���{K�/HΝ牯�5sS��ixدyD7�{���.YB$o��Xҕ$���:��Y˿?���d�0o^5�A����Kdҧ٘�����Vb{f�Q�6 :>x�} "�6,**j���ex�ٳ'������7::9�;{�����`dbb�)<��ַo_|��ٳ�׬�-�t�2\���P[�cbc B�<xpŀ�m@~fj�Jc���i�]�B�p`c׹sG|`n�����cǎ��lذa��M�k�޺u+��������wأQx,0�\�r����q4��G�}��904(_/�U(�7oΘ1�e˖�Ϝ��e\��Z>9|������QϘ+9NZ��0$�'����:u
4���h���}}}����nd��-,�*�%�	_���&�H!,������WH�S^��")�7'�
�/"d�P�"����ɲ����<��:`��������z%p�\I�L�HK�)^^\L�	�!5=�ҕ�<F�3��ٶ���uj��Q"���8\/���[� �)��N;�w/�P��U���\Ŗ*��٣���9���/�<M�E�)d��Ks���X��|�,H
�Y��T?}2s���V����fĂ'���<x��nЧ�޾���3{��-ZH�D�"��$/[�<Ϥ�::n̫ܞ�p7�CD��0�DL�_��u�3{�ܭc��1k�:u�ܺ��a�
4#���ƪIcSU�o��U�3��Lm��,���];�ׯ/�ʴ�%}��I�3�B)�b9E���s�4#����K{(u5�q��gϗ%��ɾ��\(~�(r��J��}G�L����3m��=�ww���޽{�7L
��/T�Ћ/������.0�S���@����w�؁�?t��#���ͅ����d�EЍ�}�]Dd$�gO����
<
��7��ًq��}��]�����b����3gNըQ���#}�ݰ{ϞĄ�5k�����fj1.6�ĉmڴK��v��hAMC}�������9s�8p�ʕ�%hᓝ��?1��A\�|��LKe9����ɩ��#G�8p $���yI�������YS�Q�)����>�,��F ��#
���h��GQ&vZmE	�зII)P;�Ν�����jժr��vv6d,��rs�q���p�+~���A��*~X�@Q4x���eEr<���۝��J�q7{
&��Ms;�:���ٱ#��
�1P�71ʙ�5�PG������A>Ǯ�w���]����ȈPu�_���Q�b��q��k�tI4�s�=$�����i�
����-�]���S�`s���I"""�ʣ�ddTJ�LIM��2�5��u�x59GQ�?���{�؄��x������x<|�������C�*5,,��2�U���nF� �Jb )��H{oܸqt�ļܝ�rv�����`18-T&�U�UÆ��j>��G�/��(�;7��R�0��|0s�(��-$F
�,3�§�˄|����D�r�J�>�	�"�1Y��좒C�h=C�{Z������z���ѣGa����wp(]��h������vl�Q�F��Mb�r*��wa�V�JNN�|L���X��<o�X�
�~��P�w��W�_N*R���g �6�6�����e�Ο9k��dom=eʔq�Oƈ�����ܩ��p��@�kצ�ʅ
3vl�,	?q�D����B[�JTM�e�/_>��իW�����b�crU�Zu�Νu��svr�[(U4�����]�@�b��W:`��/zt�'��:)1��?�ؾ};`��'T���h/Z�KH��/�ھeV�>}Uf4ʭ�>gwA�Q���-ڼy3�C��`G���+<��W����66v��N�<���k7Aڂ��aa--�9R=W&�
fof�'�0hu��܆��S�q		9�����II	x{RK���1���hI��e�,ռ��T�[a�i�?�����C�/�hq�Q�3!�B��]9�?�l~N����z�*Kocm-7��@�����_��䶶��$@�u�b�@�Qu74��Ǐ1�q�E�LֶlY���7G����&W�"�9�T(�-IBq��˸�9v4��]��܃(�W�FF^�.��ݺu��{���+88�����O��(������IZX��;[�;#�W<KV��Z���<':�%�~Q���۷�;Ń+�1]�q�DJ�ԩ�&40��i���t�L��e�>4��3��u�9�;@W���C�E���������A& �x�Μt�Ku#�V�+<��������"�{y��&�6m�
\=Al�N]�ؿn��E���k�N��d�_JJ�`ǻ���d|S��uȎi/�h��������/������QQQԜ�u�¾'�|08�3_>)�@W`;:::9;�'#���sǎ1q����!s�΅r��r�n���_�`��-@ �v����ʕ+V����L�(\�t���h���t}�i��z9�Z �޼u���yذa��0�U&4�i�7o�ܷoȟ�O1bĝ���M����ʂ~*�&�;M�={�̟?�H�"#X��W�Ƀ@3��F?3���������͛>|Р��+�6i^/�z��#1
����-Z4�r%hB@7�f�CQ�Yܡ�4����-Z����CLB2�w,��J��=����9.�]�>-�������⹋�'��O����޽3����h�������Y&��"7�N�<���c@�S+5��-[V�^rb�!~h��c�	��*#2,l��v6���A��,G�a�`=������D����C��:-�˼�(���ɓ'W�]ïϟ=۲eK�ڵ4d��af�@�q  F	%��J��G?�

_�dɷo߂�O�:jq�����%��>rF�/�����YiP�< ���=p�4��,��V\2������Ir����6��/�**s�O"�x��1(���3:
�
=���u������RSo߾��Hg���޹���t����:��\���*��BY��s\��"�+�
݁����Kwww�L�9�7;)*i��솒����r2��w���0_�q0o��q�ڒ�t�^�����<��)"�yA�`4�e��S����y{��(Dۊ��Y �F�6m�;v,������C��41�Cb����|�
A���T:8:�
�={6�b���"bQ�T)�����͏�P����G�Rr1Y��H=`�|4e��9�����5y�����;9:�i�
X^�tij��4�j��Xqƌim[5=�⾽{m��'O��B�MK�9�(=�31���X�1c�lݺ��6R4��6������h2T��JL��E�����y�^�ˮ]��ܜ0V��{�e*��=�,� ��`o�����Q90�M�6�,pdV;�@��h�VV��̛�����P1c���W7'{:f(�6�)�
zALHJ���z�#>P�h�����K���D��� �������E/����-�z,>�߸�fF���pPN�v����6j�Шc��>��.]dәC���S���6w�777Ph7L�	&̚5���ӧ�r�A�ӧO�mg�^T�0�0�`Ĭ[��X�b�:t����Q��3f��y�=z�(���~���D�u�&�600�]��t����,PnӦ��� �	'��-w�N�&%�Ճ�����Ա��}�L�r�E q������;���ݻ�� ~��Ӕ�Q�_T��ի�trr���=z�ŋ1F��0�0h^�~M�q��ҲU+�̙�������/��+V�"x	kae�fŊm۶�:u
��;p� *Og�Dy˱< �-���۷˔)�7�g�����,��5 �E�2�f'�~%H����)�B�V�SYp�<(&d���X
�M"]F�5-k�:��ʿ"�/�	���������`Íq׏
�Y�<���`+�
�?��?�1?�"[�.�Cj�N���6?Opy��'QE����.^G,3����]�����.^�8qb��E�/�d�o
Q+��m�H����y��ıc׭[c�`�B�������]�]Ws�1�9��?rX�T)#��HivvlO�E 8�ƻ��tA�V#?�Gq|�Pa�߱c�e��`��X��`
�<@cf
<Y��d���輸fIF�N�҃���s�]��W�ɰ9Y9;�����;��bd��o߸ioc��E�l�:��S�ؼV\=z���� �ONLkټ����)��Ѡ�ꘔg�90�C-EhZ =t���%K ��GL���-R1����m54����%u6ԯS�l����V����l�h��r��:u�̝;���!(h.��KO۽c��͛Ϟ:e��ķ�
y�V*vnۺq�:�����EJ����j��Q�0bٿ1����!&2�q���%{w�r�8
*�nݺr�ʍ9"�+�Ϙ:�ɓ'P
���;s�)�������O�b
��ПнC�ٱcǬ�7o܀�w�����;�^��T�㣣F�U�R�ԤD���7���===�3���yf��O�{����ǌ�:u*�!$$W�����������۷�߻׏�6���Ç`�^�|���?���+V��a&��?h���W������?m�������[[�eߕ+W ��|�i���V���箎�ڷ�Z�j�"E�u�� g��U�B��ׯ߻wo����ׯ��l���9�w�n�n࠾�Y'O� �nՊY�=���CU���u6�+7���DC��T>  P��E<u��TrquM�� `d�
��T��G,�wo�2����A�D?�t�rOg
�-J8�Ǌ��L��������Z�ל�����4
z ��M��VG�YG�cbc���q3 �SCZ:���T��~��9���SRS ����U����E��uxs����O�i�.�m
�����Z�>x(X��nkg�m��MO��{�(.�[����Q7oѢ/^^�v�~�Y�fai��\�N��	��c�p�½{�B�Vѓ>>>>dY����H��'_�������Wx#D($�$��������ȼ�/_�kgӦM..Yk' -��녤�d�\�J�����Ȑ"v���=��<t�c�a��p�h�����C����pd�>���}�6��I����߈�<8V�G5)��|�L�s1�߿O�pȧ�@� ��<n��%'�}�Q>G�>I�Al�6kG�rxK3�]ɾ�nEFFB�����-]��͛���e*lsc���@;L�J�*e������:u��tmذ�bŊe�֨q���ܹ3� �W��۷o�;4i��t��d���|^6nܸr��N]�6lúu �ٳg߽{��΄���Ν����9�;����� �p}Ĉ���0:���M)I���NnD�o��3��#�#޿���_�̙���c?��}�s��w����/_^�n]���I_]0��Lpp������/�566�*U��^�Zŝ}�lmgΜ	[#>l��@���pl7tK�~�ncA�޾����r�ӠA���ԑ#G�:G����Ǐ*TH�˰ ���{߾_��_�~]�`�Y�f6�	}��/Z��C�up�5��X�7�藐~��/?��s~�%]k�f�ҥK���Q�U�ƨI��N�N�)�cƌ�XH Y�i�C����GF���W�(��Oh�b�cƎ%�g`?:�����O?-[��֭[x5avbB¸q��� ��F�CQ�d^�L�ڴ	<s
b�iݺ��9P&��?aۭ��4V�i����ʹPYDDF`Vb"���guj�U��T@>>�y��2eʸ���<u�|���Y���B8�(\///���e�jլ�OHL �P�DI<��D���ĩ�o�>t�|�B��g��x-�.!p�)��`l�>#���1ׯߠ��=J�ltƁ�!*۷oG��H0�,y���LXt,;�;�3;��<���ٳ��_���澾�@}|@/b�N�<y�̩Ph�*�e����?R�,X1ڇ���C˟���ܜ���z������}z��]�o��a��(�XZZc�%�d���2�2���S����kFj���hԩӣ"�G�>y���<��S�ގE�MLI曀l��VN�FM$/�*�|C��n͍	����W@�񂿺���3������g�>�߿����T�*���j�V���Ԙ��Y�fО�<�(����\��3h�N��5|vBد���.�;7oޤ<�(�����v����{@��94;XN���W�Ykgvr<y�$��F'׫W��PVBi�L�����I[����( �E���))��� &&���z�oG}(��xl߾}��7jF���,���e*_��/K�Vm+V�r�ƻ����壼gЀ� �_��
��-Z��*��/�O�3��.����H׽A ���`?��&M�$%% -Г@T":p��iӦ4�2eʔB<�aDx$ �H���*�qb}�m��#F �'M���+�^�F�ڵk�8}
��|��|���ӧOcd�1 1�sԸ�I��7fК�k�ݽ�d�4y���,�`��<��a^�Jx)�k۶mu��5�U|���|L���v����8�l�q��M�6����E���q�^�cgܭ�B^>G�!�����A�Y�zkk\Ǔ1p !�4`�`4�:qr��u`*�yy��%�wque;/�]�jղ%K�?�?��B�
��*�W�`DX8*��@��߿ȇ
(�k�E�Ff2KK��];W�^���IO����I�5K������Z�8qo��y۷m�.ܾ}{��3�O��9^������
��ĉ�O�:O�A�@�������LK&����t~HmZ��	%K����͛�����/S�B�JI�Z98z(�o�^��3��*����Q)���+w93�e&�![m�b��2��-��-t����uX��l��(f����爅����!ƕ��#�������B�(��'��}]�,Ҍ%���V�^bMQH�3�*���d�����z5����A4w�s�"��dgd��0@�I5k�trrc��x��2���d����Q�,�ʹiВժU�E� )�Y��a&C��Z�k����	�υ�[�l,׽{�⽰{��((|}� �y���F�_,�G�mުUJb"z	�>�l ����'��u4����}� @DD��o�m��H	�`��k
F�_MA�F�i��e.���;�������ْ,p�K�.�yd5��˚5k�~-Z�gϞ�m�j���8�ǓH�9s��/^�X�zE���/]���}D?��6��1�ʓ#{yy�Q�Șؙ3gBZ Ɂ�+?��g*�ޭ���+�����֭0��5`� �3�,,&}���G�0_��G�V�ZU������=X{�T��ťQ�F66����N
�7WХ�� �:�7�<�RRSp����'VػQ����b%K#�sA��BW`A0X���&���J�9� ;v�h<�HZ�(��V�RibP[G'����j!0������իWc<<=�� e֬Y�{(Y��D(>!�����f�����l����^,i�p\�X1tT4/h,���H2��J�*����K��w�ލ���E�+\�0j��^�p��ӑ��gFǓ&�x����˗=��1d�W�B̔��/����ɩM�6Ѝ�I���U�.X�d鲕�"�f@Ŋz����4q�D�'�Nn�P��=�Q�Z�c̛J0
��eұ� �exK�������	�	���u��:�6�N���r�*�+C��C��G�ꥡS��@�K_��s�勎�_��µ��2D���E}�%a�d����e���w�t���ևA�Z]��7J���Ս�nXPG{��2S��4F�^g4�1�!SN$��v���Sf��@ �(�VRa0 ���>\��>���#yM�������G�R-Y�|�0� �Pm��3��k���+�9'�d7l��"E�@�A+�8��C۶P��g/�H�b����"S*��t�}�����bA �z���s�Ώ?�����w�&  �'�P��
*����
޾}�=��&�H� �U�V7o݂� �r��LKN+�V���+��:t��[�����/Y���],pP�s�o� �a��+�w����<9:jw��}J1 ӴEjP��ںjժ���T�ڭ�<y�[��������r*��e��ф��M�0v�����
I�u*oy̓�@��R�- �XB?�'a�ƍ��ԩ+�s�h4�#ն]K�ia��������.@�a��?~�����m����ޠ^B��عs���z��ŗ^��0��
�2�5 $�Ή5�R�S�(Qs�s�.�b��AT)�;��6Y�7 ���߼y3ĉe�5����S=D,�����ΞEͧN�
ȧT��O�J��,=v��?�(�0����&B_�H�0v�I0������#y���p?f"��N�V�Z�/��ѣGhFѵkW�o��APP�p�B �B5֮]kŭ�/3�ԇ���gϝ��@(
�!;cm�W�!��/�wv:l����[�h�]ϞӧO��!O��~��#/��ߊ+�W���:�eFvv��`�3�֐ζ�[!��z��\ik������K�e��=�֭ݱ�w��+�Uuz�1=#i��Y[�nub�)ٶ)��Se,�y^���~��*�O����A!����s�����]|�8k��BV�g�#�;Q�4�2Rx8�Q��8�_Q�X"�tn��kL��X�h��:���:��l�W��QгI�E�x��Ҭ��?`��ΐ�;#)9�+~��'�G���Q�����G�޴�?f�8�W1�ws�t؋0��o��n��5k,��5آ�U'W�%K� �Ю�m;�D2������@���g 7����S����f̘ulmgeܠA�����۷����Ρ��� �a��x�p`^A���||`�Yi4 
�.^�gfB�9r���P( �"�6�N��x),����C���˿��0a����|ۭǩ��qqȐ!��{�ݳ�� �a�@�`�.]�\�S�I�&�f͚E`�̠��0��4��V\�:t�������Z�xFsi�Cq�&&�N;�{<�f#�Cɒ%QVL�Ԙ���
�����@�Ǝ�ރYY�t�իVB�W
�������˗+���B���ۃ���V�]1h� �\�A�
��h��NƝ��]@�/d�u�֓�L�Q>x�`ӝ;w���o_�E��ރ�E��A_ �}�����̝�B�i�cy^>�t׮]���֭��Ƹ�:�{���
��СC]:w.�������i�aZ��|!�-:�����Q��N�u�����A�v���>��A��;w�vU�X MCI�|��&映�lܸ1���*�.oNNNqqa^��Aak===����6l� �{����E�.^"1.���łg��b��	e���1c�T�NQG�yK�i��>���R)d
[k[Z�O�H�r� ��x��bk/��C?Й4���C�aÆ9vH��P(�������a��"��I��Z<��j@Ǣ��'�$�����?��4�]f��O�ZY�W9�E��I�q���_�d_�e�=S2]b?�M`*=�uFRX�;�j�3B�a��u�~�O��J����`�A��=8�Nk0ge�9�ع#K-��oo�V-�+�i&>���	�+p���3�F�ھk7�5b�y��L1���vT{R�Rl&���,�������9(L�Q�-�m2��Q�6ӽ@��k��/�Q���L����*J��(Wd�^m���x@��s�9BtQ,[��{8�P3��6+�}��I�m|ݒQ(�E�o�"�C`��������dـw���:�����@j�6��Sv6�3�K�|���G" W[V�?�T�ۨ1�Uf�>y��ׯ�'??fm�\��@DS�fF��CQ�r�)>p���8��+��x�ر�u�i��-�srZ�k�o���æ-�
�A6��ɑ�qvN��! 
ģ��!�^��U-Z4;}������W�U;:> ��yxx�%����N�0���At�կ/��y(0R�/��z�K��AqJLJ,\����7d�U떏�<��8u���!%5�����ϳ���/���&͚�9.`a��5��i߹�ݳO����?~�^�z$�~>W�\�*U�\bJj���¸�N����~�d09s'�H��y�-�h��a�$5j�)qvr.\���y�N�N�޾>U�WKNM�4�{������=_��gΞ/G�<|�d��ΡZ���j�u���֪5RN��ɳ���� ����{~s��u��ʕE |��ǣ{� "���;�v鞐�;f̸�ׯò�ُ��=�Y�zjj"`�jkg���٢E�Voo�!>.n�޽��0���E�H����>Q����1qjK�����E���p�+Ø�ȵ
�޽?o۶�ڵ��v�N���0��&b�V�N���ٴq㕫Wy�����nt:~��(l޴%9.�Nc�g	d�x�r܄�M�`=3���#��r���w�޳�,eƺA��}纋/�9y�\�
� ��F0j����`��蓼_��ؿx��t�����߫ϳg�T�))��<.�Z�t
�^i�+�T�Q��00a�J��#��k��
f��"uKKb����huF�A���VjK�Dod�Q�� G��g�yez؊��&�|s�Ba���PZi�:���{4*��W>sTLt��y='[�!`%�$���H�֙ 1��"gr2�l��l��i;ҳF��<~��9�KEȵ���Wo+U�D���R҉�j4�����X��0[[ۏ�j���v����))l��Ғ|���]=<|B+���m�)�>D�j�2 @t�@<m"��!�.��B��f�P�H�|(��Ϥʩ�D�J@��@!�M�ts��v	��¦33�S,[t#l/<֑q#-��o�@��N�D�P�_rcD+�.i���[�"��8Ѱ:�R,q���D��
z;_�|��%:!S7��O)��=JD}r�m<�_�x1�i��s������'1��3�i�AAA�-f�;y{Vi:_����V���jw����>-��Yɸ�8GG�NK��_Qᄔ�g�t�*�V�bŊ�g���K~y {W����e��dk��B!��!�&M�
��3�G�a�|��a1�fWp���[g
�&0�5��"��H�w�%�n�*p�o�g�,]�4�Eh�ߖ�ީS'�o�:u��SV����ۓ���M�M�6�)h��|�O�;w.f=��j�DfGul���~��g0ȩS'�%Pm��0R==�ủN�*S�<�I7oN�>j��ׯ[��hȶ�KK<� m������֏��A} �P/�i���R���{��D�A�j�\�W+V�����fEw6��3��L���>zv!�mh�%@Umy�)��p�ԙ5��ʢID.&	��Ȏ]�Q[7W�z��	�����I�&)�5x�������b���T��a�����ݖ-[��aim����]�Q�����ω��t����q��$�@��z�y�/5��ߒ���"""�
��3���/�R��R�#Ƞ�1߬��[j
s]������r'ed�ӑP=�`����E������i��� �~'��A�g5s��i�/˸�;[Eh���$��8�,&��=�hj��ȧ[���L��g�	h)�r�f))���;gY��D�J�Bi��Bo�P�s�\ ��(g;����A��։N�b
�K/��~��U�6m�V��|��'Ov��&�#��ꄇGFFB����[�zy=y����?�o%y�G
��S�k
0���=��?���
���D��<19%MY�'�%=��1�DW^
I&��ѣD`��,�^e����X�L�b�޽{���64�7��vv��jժ��vrv�b�H�|���W��bce͒J�4|������Vq�,��!��{�|� �F�����d٨�J��N��"��E٩����ye�Uda�x(�����-��I�����'�LZ�����b����ku��(��G5�|�8��.T�C�]V��0�+@,��*S�S�=l\�D�W���\�gᰴ���L�8Q�G�6�=z􌋋�a1 ء���
�J�IIN�0QƯR�K�_�[�xr<�'�'�����=0�_�|	��_+V��'����T�P��			������PMC�� Aa��9R�~NLHNH����f
#�����E��YZ�EF�3�~��L�r��yAA/�@M��,r���K�z����7,��?~���̬�A������~���jϞ={��ձ}�-۷����ݻ��][�
n�[�qg^9y�Ӳ ���gȏ��dll����f�k�h{,!����ٟ/�B@��/��տ���[�� ��m?�Ė+���9��)��Q�3d�x��/_V[0�_�h�/^<�s�TٲRU.v�W�*y"Nf�&%�;��ӟ>{��טDPn"",��`h�p����#g��}��}�������� �j+��U�6�h�Z����Ry�1>	]H�KM
j�t@�N�=-���Ќ��B|8���FL:'H,	�C=7L�Fl�C�0tb����N�q���˖-��=~��̙s�֭ƍ��{(�b>�
BP��5k�@��]�v�%,j��/'H���c�ò�m����R4���hF\�+���DV>9���,J����w�rN�N!<׭[��B���-[�D?x��!t 0�.��=z@����788:jy�1���#�h�m:v���3����S�L��ƕ.]���B�!6�'O�ؑ98���_~�944�z���˗���Te�3�,5%e�̙Çg�r$	�(�@Bl������[aXR(�O�բ�k�"���3-����r7�����bc�y:"0s5Vv��a�����]�[�yC�u�p��4d7p8cy��Bh �R�-(4Y��Z�z��u�S��& @T5�XbBH�og�5Yg<f�@��O��ں��6j؈F�������;�BBBF��wvw߽};8e����7jĂ������>z��x�|�1U�w@�-��+j�ƨ<v�ص�w��jTB[b޾�leÔ�UO`�Y�V-��,!������+w���� �S��ȇ%V�fM��ϟ6o�r�'Sd1�"~摺�\�u�`�e�eEm6i�ޫ��2���`e(|v�xST s}(�Sttt�Ĥy�ŵG)��/d9��%���:00�P!?#�� 7[�n]�t)?ti�ja!Wf���Z����;����Ea�R+��V�Q/S�Y+M�ȼf�My�����O� S���N�
��׹s���_����?��>��k�n�f���z� H�^�WA� �G����(�R�&�ҥ���H'�I���~��ٝ�l
	��;�wo�;s��9%$|G�Jم�Scy%)L;�\HĘ����MZ��Z7�m�5�|��ԁW���Y1���/�.%���jJ�pvUi��]�(�)k
n�����!r
��ܹ}[��B�k��ɒ%K�M���v��?����U*�������(	��5�e�#�l;#�ҚӤRn�iF��ٗ�e-:�8+�S:��4u"Z��2�Q3/��h�bg߯\��_�;7k=b�Z��#&�j�j���ȏ7n޼y+V���lyy�`̜�:9߾ywϮ�?�`�JR�>qr����n�9x�Z�n}��U+��׿Vݺ������~��}�?x�8��٧N�

z~7����q��d����ڵk�J��;������ |+�;�:�yz2_���X�d��%�"���3� ��K
�Α	$K�Œƛҙ���S\Ll??OH���s�ӌ㦎�;w��~m"�U,j��ͯ���qwc�<������^�ٖ�X���@;������P�--fs̘�Z��wO� L�����py�ҥP��:�'O�L�y��[�An�~ժV>v��޽���o���ʫ�e+'"""v��u��A�쁼���_~�ӯ/����lM�(��M�S�%��9ʖ!��0�i,kБ��ُ�U�L�h ����#������*r���z��\���:`��f�n݊�f޷ ��,�/�pdh)>>��]�=�drn#w�wwc>[X�.^X�*%3�3D£��o?�Q�s�ʵ�N6Sa��}����۷1�EB��J�{ː�f�˗vqH�I�`j�>W�V���%�Rؼy3�� F���IԢ`��ϻ�[�B��%K`�M��\��&��.X�f�&��hV�o2a�:�˖-[ܜ]j׮ݥK�뤇��4*�	���~hٲ���{�R�̪W._�6|��I\�;s�L��d�4��̙3x�:qO�@���)�۝;wBCC���Ѐ�@�}���X�v-����yŊ�-
���5h��*U�R�/]���/�6g=rĚ�G�b
XuN�\�stL���|���P��<BZ�q�F*�ҿ舛6m*R����R������Z��,��D"����)]��o0E���۱�]�I|��HRe�8i�UF�tˍ����0���X��׌.�VEV��e��|�4nf�믿R�G�d%w�^��A�6���y���@������&�y�eQ���n·K�g~^�W��pw�n�S{��mӮݱc�|}��R�ѬY�Ԥ$�;�ܲu�n�;c��Z�
R�Of�!�`H�s5�1; z�'�����2}�t@�=z�ٟ�I�9CX�^=J����S�؇~���	�cԨQ,���);�n-S�LѢEcbb�V�o�W���bժUK�)CܷpѢ7x{��3ZΔs�Հd��Ϟ={�ԩ8��nѲ%͵8Ӝ��c��HV՟�(�O�FI�V��q����"*<<|ǎlҤ	tn�,$&؈I}nsRk�m�w��p���=|��K�5l� �w`%��v	�!�!J�H�G?|�x�b��Y�d��&?FQ7��
� (R�������n\����ۛY�e
�tp�lZ8e�f�+n������H�ڵ�룷8���܏�P������?w�\RRO��v�Ǝ��!s>u�;��;&fR�(W:Aة���k��eF@�(#��B�������ra�!����ȟ�8s#8�E�p��!ǃ�8,	,`���'�:x��r���k�%rA�7J�/i�R%K�-�g��4��0�>���7`+*G�`���Z��>Y'�,.Q���{�E���17]P3@kJ��s�=e9(0���=�*U�f��y����������� F,Z����{���ŋ6lZ�h�u͖�K��oHp�ÿܷoxGؽp�B�4��+T�>7u����ZMJ�}Ē�$nܤɃ�|2mƌժUQq5eÆu�f��߿�cGڴy��ʸlpw�(�D�b?��S��P�	�_��L����!q�X&{��~�oݦ����?��ʕ+�Ѓo[���"�	��xqdT^����AÆx�2e
$�-�7������٭@��"#��@�l���`E�U�Xj�9M��(� @�&.��_�0#6qC�����j[X�*�|���d�6�"�$�M��i�A�+���}��ݷn�&�,�I���..AF=|X�D��ǏC��;b���"9�ɓk���g��9��Ʈ_�nŊ:^�N��洴������nҔ)��NuPiDm_���
F�ּy�b	 L`N��A Zv��AD�N�ЧO��G��T�p:v�x�ȑ�6n��M7�q�b�~� f�<\�b��۷׬Ys�Ν�K�bɂ||�����A�6����ڶ�4iR(�<�b�lx�*���;j+�
H=  �ҥ+�7��F<y�hc4���0P��zT�P9�`������ӷl�� ���0�
V���{�����/U�t��:|��EcJ�����:�Z�Z�a��޴qs���aw/K�{h�햚*��.�R4@x;w�t��h۶����pb�$���*�N����&1��.���,�
gY�x�?P��y7���!�xM��)0��T���C�=)��>4V>��4�9ھm����=��7n|��~L�єγt�
��!��t#�)LG���Z�1�mߌ1����2���V�۵k���QL��<Y����7˜ �\@�XҲ��9�A�����x�� q��4O�7����iͰQ ��l%�^�f7p$<\=<0�[�n�� BBB���}���v���3�V Kau��>�[3)�P*�j0�䧢X��i�>3�T��&��Nʧ����oР�Q�P��
����{ �Њ�5�����ϛ�`ݺuk֭�ծ�g����PSD��C+�R���T���D>��<���W^
Z�~=�J\L��0��/�Lrqy��V�F��JjşW���V�6m�?����&��:��T|3�p�N�����.|��'�T,o�|�.@��7,�����ׯc`K�.���)#;�P��ݻwy2r��͛�.����I�8Yt�y0n6 \�5lX�`Æx
%�g��\�͙3��ի�xAB�e�Y :�&6��kO�����:}�4(
#C��� ُ?�x��%���c�QJas�'a/0�F��	��� m�@���U�)ҒxMR:���ٳ}�ιx�qH�� \�|²k׮_/���ܹ�{�^ ��A�T�I"����k��	=I�׃��A����=���*�g�uX1L�4�K>\@	��b4�&C件��Ӹ808��@�5j��߿�[�Z�ݳg�С���
`���p`�f͚Vm�b�0ݸ��͛�d'N�h�/\�s�v,o�p��T���?񚸪b�P�6��1cƄ/nJK�c8PV�%�2T�-^L�<���{{oݲ�}���F� �m�e4��l��g0 l����ի%�{�	��
���*{�w�o�	R��ɓ8X�A�U�������6ܲe���1�x"Պ%�����D&ۤpt<��/cǎ�nӦ��u�̌���,�7�V�$>`�q*�������/��_�5�T:<T���7MLHe��ܺ�ҡ���&��;PN��p��1�Y��͛�1zx����.����/.�yc�M����Q�i1%�
UD���.���M�"����=�%����o��4C$*u6�|�*���� 2H׷��CO sY=��c�g�FF� d�!G��N˷d
[����ԴEs�ٮ]�� ��}PPA0(u�ճ�l�VF���c$��Tr�Z�n�n]/_�s��  C
s����w࠷��%�Z�B���$k7�9M�x�t��&N�*?w�����N��u�-Z�\O��@$�)��Jd��������O�f�l`��Ç!u���TD1�P'g� �u�᯻�Wj2�0�n�]��Z��H�`�*��)[�{��۷o�h��Hi�C�a�Ǥ�D05O`U˖-���3�����^a�3�)[�U�֐[-Z���oٲp�% �f��ŋϞ=;!!b��͛��z��S��](�a�FfI@,*H|�S0S�1��ܹ��v�ֻw�m۶6�*�?~��_�Y�����j:(�,���P�$BZX�`X�F����o`�*9�yzY�'<ckϞ=����k�?A6����n0�/����� �,Vn.A�__͞]�N��u�H\i��g,���q���D�ƍ����6�~�Ν7n���Y/B��F����w0;@�b���f�Хf}9�h6�>������g7y�����h��[��`�H%_�J^�!�H������9e!���5<6���'�=�fΜ	�I~�6���I$�ƺ���¬A��]����	0�'`)5i�%2��;^¦Th�_=vԨ�{����J!f
h)�dI�Mnݺ�n�U>�$�	$i��M���f��^<>�rذ���[���N�6M��>f�+�Qh8���yܸ	k���/�����6o~�];���E�x{y�8;?������2�K7j�0�� �-J�N���vc5	�w�?���9mZ4k��ƍ�쳙�h@U�\ Q�-��}�m�}�f �G11��4c��`���<R|/��Å��nG��Z����O��E1n�D���e˂9����9O�0�g��Z>Ƞ@=t���#���.�N��+���#&�#/B4��6}�T�_	��+�& �.ݺ��޻�شiK�#f�ר(�;�Yf,�I�
��0��$��Iщl��'����$��D���F��({F��pr�I���BA4�I���[(�����"#}�\��10*>�i����? ୷����� ��$��h���=x�T��F�U�<�'�l���upr��t��q����n����M��}�9H5�8��^S���2�r0)�e0ЦT\l���N8t(�Yw1�<�$=|/,��<A&�v��	0kb�"�,�x��mHY�
�X��d�|JDϨS�I�y�������kh�����͛X��j���I�E��.�5�G�Z=ˀm�I<�$��i�f�8��i�®nn�˗�p�t<�K7		�Tv�e���3Fܿr/�E7�7(d6l�ѣ��y�|[��L��U���V�Z� ���?xz�S�h�j�
(�5�Γ��1��D&MtРA����;��pcf���=���ӧ��3gJ�Ғ
2�����ᇨ��Ŋ���V888�����K������իeʄ�h�����<N�4i������#�BU�|�Νۡ�����%`��˗Ԯ][�ֵk�XxUj*�eNr|<�B39�
���(A**�`�ԩ�>���P/Y�dʔ)@�п!S!��(��T�� �����T]�t�ۯ>�:u
X�\�����2:}�t '�4,�ݲe�@�� M����+W�?�������dHr�ѻ�޸z,~������ဉ2g	���yON0�����y�����`Q��dg��s�^�x�믿.�+�@G�� ���J%D>���D~��E
T�R��}�lL�8�τ�Y�bňѣ�J%��իW��`dM�D�s%.��[�6�ntX� �hG�bccAB�-�F���dY� ��{���e��ݺva����[!�-`B�@G�#@f�R���,#���s]���ع�%Ā;굘\�5� �p	26�l7=��	��Gr�	���̢(�M���8�x`(5�ĳ�3ĲVs0�X�L)�g]i�*o�����w��Ù���x��ϝ�	��9��M�"W� 3�%�� ���W0��\����������8�۵k-��T� �?�����KӧLV+$�P=+x�[ˡH"�̢�Mϛ͚^�r�ڜ9 5�f+)�R�
\�:�9s4n��f� �����j�\������<�8;��LOr�:���A)�I�K��5pK�MKI�rw�Ҹ����OMNMIL0��*�1�bL�\��4^�s(\���j�ݬuһ��Z�T^$���9_-]���_�0n���1Q$%%;:B(&��dZ���M�T�j���b�hV��qϐ!C"#"��������j
��#Iz��;�䞢8���� �@�a��׮��PAC}z�j��m-w�^�be�Fo8s�I,ܤe��͚7�x��R��O�p��eOrvNMd�*K7T���QQ���D��k�0�~����iD�M58��qG����KZ�l6z���M��غe�ȑP2(�O�ܱ�GjV�\�s�hӒ�W��Z�h�����$n����C[���T�`�d�0�$��a��R�[�DF{
E�5�\@�V�V�HѢd".��7�y��Q��t[7/��K�T�Tu�����gHK�i4Q���P�~D��-�5J.I��c.<d���	'���.�b-_p$<<D�R�$'���_kڼ���ۡ�c� �FDx��]Oυ�mٺ��8���߼e���C?AAATM�~��;�k�j1�`18��K�&L?b�p����Ө?�,�����s ��~�N�EK7�R-F�}HR(�K��|�E=|���R+C��J�v�p���2ޅ2�`��>}�����*U�ի�p*�_�֭E�r�F�e�Gl;hJOO�#��7o�cذK�.�P�AA��
���/�?�T<]�����sԨQ�)o7İ�{_�H��&�����p���zu�׬QB���`6�ճgϦo5�+�$ֱ�l��N���$4���71!��`r��3��K쫅�`"##��c�C�����#CJ�Q�T��]�2y!)y�xG�2Y���}Z�e\ ϼ|���v�T�X��3�=�B^5'R�l�f���t5_!�=m,�4k��3�����ϩ��c^�z����t�,J�^�|Y0��ܷ@:�2�����Ǖ2�*U�_����~��y�rC�A' C49r�G����U�#��Yٯ�Δ�$G'g0tH�ӧO7x�������@F������v��1bsFnU��Ⱥ�MI�˖//v�U�V@k�"A� ^���G��.�Lp(D~g�c)T�P�Νj������!^ėe�2@(�+�:�z�S��n���y�sT7	ு����yv
�*��$�t��D�C zy��l&�2�Pa�O?�

����q�u�	J�V��{�6x�ɓ'�qW�t^E7��t��H�c�&[�v�uJ�f1�`
G�<��9$Ͼ�\��~<{���Ǿ�8~:�t�7ި[��Ν;��D��V���X:���?�5�Y���31я�<=�DG<b�=W�O?��~�l&y�����aÆ�<�LRbb����Ƣo=��a�G�nݺ���E�����쌟�ת�w�^�2^���ǡ*<�}Y���O|�4(8��~�l:�=��o�>z(�Ɉ�����Ry�:f�x�R���/��-��"OMJ�[��W���d�Rx��[7��ҫ,���7�d�s���K�1j�=�w�-[��p�WL^���:�G�dS3TCn�ݲiӪU�ʗ/7`����ﮟ�:��nu�޽��?:t�Zu1���mGیYȌO?=��/X����|����:y� �������ϟ�REG �/_�1���Р��Z�^�|y۶m!¹�/�����J��"��+�2J�u�֮]}��%�NRrJ"ŸC�!6c٧a7n)d9plM���S�f�N���q��N�;U�\���0���`i�~��|�P�"e�pyܖ
�Y󑸺b�+xNC� ^�r� {Zj
�aҝ|����A�Lk�ʓ�mL�GXd�V���<쒓�}e�s��k�d#�EZ<{��׵<��� ����)���`��8�Զ����ԇz�0k�,�����/U*$�I�kPP���!�W�\�g�nHk �F��H�2`[ooe��#��\�C,S����W/@�� `Uy�.Ŋ��>mƯ�� �ءs!��X��/m@��=T�\_Ǎ.��JUG�I�}ة<��È,u`����ׯ��_�aB����t��Jʴj�
�X�b�!�8׭��C���`�hN�OJ���q��G�RS<����'�{�n�N���f0�k}��?��"\���ͻ�v�,��R��4p���?�@�� A.⯲n��Zgxw��	}�LZ{�@{ �D󳿜5f��ŋE�7U�^}����}`�x�W>7l� �(�~2ע�Æ����ٳ`�	��c�v�rݺubG�}*T�бc'ɖ��I�g��e֕i�\�/�l>|k3��Z@�lڴ��[�!!i<u����A�b+�ʤ�]�6�` ���P���h����<2BTsfR_&�+A{�B�(��{RN�V��S�Q��Dstqf�j-w�2�k%UBr�O�?���^�nI���S�i�
�`p�oA�C��Rq�T�hѧqq�+XD�Htp �� ,jr�q�`��Y������+Yֺv���9B���2��&�V:�I�f�hD�y����f͚����u����Y��W/_�Թ���s�r� �1�͛7?v���e� ͪ5j������n��A�9��?E�7e5����ӪuK��qOc��\\��;���1K�,Q�-uk�U��9sJ�۹m��Ag��jV��k�.��{�A999&������"������^�L:~]�h��)S�׳R�d�����ʊ�1ԋ�M�<�S�P���
aH�t���U�\�@�5l�Ϙg+,&�&ml[x�!�ZÌ꒵v�Һ׽ӭkH�,�C�������d3myPH���@�|*��Y�C/V�p-�D���<�:ܓ)'iiŝ��țdCo,�����Z��܄��¢c���&1t���a;<,㧔����b�W,��������/�i4�̞�$��N��9�]�$�)r�B��kR���e�,\�p��q�&}_@]�%�1�`͚5�'��X;�f�{�:$4��!WǨL^�\C�Q���E����x�r�Ԡ� Ly�ł����K�,Y�^=0qP~���%��H��R�W��reCA,E��,�8gg`�,�.��cQ͞=ۓ{c�N�:i�$��C��y�:;=zj=`�ҥKѥ/����p
���6��1c�@t��;v�(^��f�+��������-��e˖��d�oWם;v�Y�CTйw�Ֆ@����&��ˑÇ!\����Ёб:�%a V1S�n�t�����V�v��(�b�� �YNC��������f{x���;u��Ø�oS�4<M!�~J0'�ԡ�dှ���z�������y&���R�R��L�s���S�YM[��x�5�/э�����{�r�ܹ��@���̌��%�bbb��A�u���%a��7!1���GG{��8;��SP� a�\!)�J�!5��(K�c��f��d1�x�B2�;f���z@0�;�s��������Ǥ�����PP�H�����g�7B�(�Q�ug7.���2]
�Rv3&[E>��!,oܸ��,�'��h��Y��b ]]��*U�rrڷoTv���]��lɁ3�  ��IDAT�|X)#F��p�ԩ+����	���>���nq��Y���P�����A���>>M�6�4y*N�Gg�����ٳ[7nl۵+� qt,_�<~Ţ��/T�дi�<<=�R�HS�2:�O���r)����F�d�G�dG�&Y����B�)��)��|��7w��л�6�WC=l����8�'���ۓ�L;k�t<>>^�)�B���0�XP������w����C��c�Q�1b�ifI�s7dVP�5+γ3%�����|T%���Ud��[lI�����aG�y&V|�
�x��˳�-Z�*
E�d�k��v�����U�R�믿�\ܲyG���0���xeV������-���اX��g�9��l�F�6mnt�V�����,�5����<�R�h�����ͧ�7__��TH� 0��0C�3�{����Uھ};ȕdC*�<o�@����\���+�ʰrjc��J�ɓ'�-[I����~���:''��M�5۰aF�%�I���g �����A^o���i��%��$��O&NY�;�;�4���K�Tw���Uŋ�a�6�?��c�ĉ�Gݽ{7���	<�ȑ#�J��s<؞�s�ع�O>�����m�vŊ��L�eYΜ9������?.��ǎ+Nk����c��QD ��>q����|���$����ǂ�<<HV�H��O!��2�l-G�g.0w�-�f�b��@fL�����9�J8p� ���6o��Tj`����w���E��w:��cj*�U�פA�@Kf�L������cp��}ʄ�nUV��`���q�L���^�x�"�k�bō&��۷�T��jU��������y ���::�c�<Wś�o��9IA$�=�sws���)�zG�è�~�~�RA�l�4�Zʳ�b������K6mI|���A~X�z^�v�<�4� �ǯ��\���fP����`������'PxJ�UʆV�lI���~��[��ӧ=�yB4�֯_?h�!���k)�ڸ1c�:������_.\�z�N�z.V�7�xl�c�ƩT*g5[\�� ,=�.lƅ�˕e<����r���B`���v�h��Hvi�~�/�?,(0
f����q(X�ɖ�U�!���,ց�D���ķ��x:�P`y\<۲�XD%0�~��b�r�"j��G׮�����g�n��yn�����.Nճ�>Er�]���խ�jI�l�8Pf
1�@��`�F�t2�nt��4<$���3d������.���t�)K�&��$�ȃ$�R�O�Y����J������r��3�xF215��J�����96��o@f�.J�-;�|7��۷A��FGGn�Q�@��L�a�r�f[�>f�2�sc�T�R%�H�];w�nP�0+D@@���1��0�I��@�6����!ff͚�p�"�4nт�Q�_~���s�n�p@���dK9�
�,|?�-��
���ۯy�X� }ɒܸiS�c!��`rx��o���\�Ȯ��d��k��P�m� ��%KB�x������.���E� �)%8��1�*� ]h���Ç/_���̅��i_}��²�K�^�J=�\�����B����9BUO��b�1c�Y�
+F�R�
�@��`��|Hk�;&K"�I:�i��jd��r��[�ך5??!�P!��ٳgCX�:u
G>��C��	0_Q��G�n��o��w�aD���y,���z�`kX�q}�&M�:Hz��BE�t���2d���+����L"y��7Y�/��3WF�"$|��́�&L�0m�4��U���C~p�}�!� �s�N��J+��<=<C��@!�	={��"��?r��#�L�ʕ+>|�Io���رc˖-�W�F��~��g�9�gĈ5k�0p ���K�in(�W�^�+��ݻw���;�,�gΜ�B��Ç�gNc��ԩ�'B޳�%K��d�R�q��u��k��M�����VG9@!`�Пw�{�I���\���ۛ��6nRw��©O��d��i'�]֮]ֽ���ӧC��k��Xy<�ٖ�j��rj��˗/?��ը�t�>����i]�`1yڋ�(S��k׮	�
� {��� �'O�"������]۴6�d]0?�lMs))RRYJG�Z�'g�_� ��R�"���_"I�K��r2�/;�{�Fu0��(0��r�A���7 ��Iej�N׬ES0��#��}A!����$
�rg5ϘK?�3�L} ���@ ��m9+�Lf,ԅ"�p�0���/Rf��dS�F��'8���죫�����Y��t�T�I�k��C|���Ð>/R�������-n��Ӳ���g>��~A��/k�cǢE���0�Xx<�� Cɣ;��μ�sb���?Q��H�T+�jV[p�ҟ~�E�5@vN��xP�9=͘��XM��(�f����U�U�89��%�Xu;��h������9]�vZ�a��j=]<�!BJ�D=���)��:t8�w�+�.5;ꘘw�;X�$^/���T(3���2m�<
񋛻��%�����L�J���f�'�89[�/,�b�K�����]���L��qO�Φt�[��@����=s�Y�fl3L���[��`֎9>`���t�q��N�;��3���j(���{Æ��7zS��7P�g.H��ޅ���jU&���E����Y��g6%.d~�ܛGaQ*?���0��ئfҴ�!%K��V�Y�%IT����h�o����Y@�`�=�a��������Gz����&���b�C�	�.�d��t���C=��O���ީ[W�Ң%�C�����ȑ#Y�F+�D�	��c@��<���֍?M�2M��n۴9�iB��>c=����M���}�v�.V��͝[�~�i}���?�nZ0 p�)XJ)Ii��ߥ}7p4[�J3(������칺:_����qIbb��3�
�9P�y��È�Zժ�l>=
"��/�ED�8�fL���	�S��N?��G�����#�׮Y���v'�2e
d��J���ڶe+`���K>}�Q�@��Z_��JbB���P����(/�E����2��y떟�|0����=��]�0�X����'N�={����'}���_����ߴ~=�{�n}##bƎ�q�L��� ޶n���o�+�i��~[vn��i�}$��ϻ�2ސ�N޸�!.L7�׭_߹sg�ϸq�@cƎݽgORr2����'v4]�paϞ=���C��:~��o�NC�6i�,)>����ǎkи���S�BBB|
0_����C��ʀ�I2Q� ʧ��-���p����*%�������D�u���� �|||��v���Yf'T�[���Ժv�˿��+�%��Q�z�����	N�q�V�b��X�Bp�kw� �'�#zp*�R�蜞������dC2t����TI�J�Ots�Hg--ijV��%�d������uT��qk����3;�����E�n�vi������s�_�l�!1�Q���#��	OY�Ti��E����ѻ���0G&`�Ⱦ���5�$Y1!)3�nѺu��ա�B]�zle��P�B
�e ��%�i�(����;����7o��	�2�V蓴�4��(YzZ//%�Y�ǆ7Ʋ�[�p7��G}�y���K �	�=t�
�[&sX9���*c�F>��R^v�&чLZ����Mz���׺uk�cG��l��`gP���1}���P�s�Nɒ%��Ю�����W҄�Y�_zxxP%h���y����i��\���୷m�FN<w��J/[�lTT�y��KA�s�ν}�����? �DОG�x�������A#��aÆ5lذI�&�5J�j��r����>�4�7�t�f	�jw �����v�M&�Nh�x�vw������t�)�.P`�����"���v@\]���b��k`�
����Q����SX� ����I��;f�,"��k7o6�_�����6��~��Z8�g��5(�e~��0�P%A��[Ъ(C΄ȿu��2���+&Q0���gͣ�,X(ʇB�7n߾��	w,��P'G�ݵk��͛C����CjFGE�Y�׶n�?mڴ	��uѰQ#��S88���/ٓ���6Z�dq��$6=/Y��|ud�~�6%H�r��7oޤ��������#�Ps@�+.\ط{7B����e�Yo����C�~ޱky������C��7d��e�T�N�L������1|�p�<����@�k׮�jK�C�B:���Ҧf��߿Cǎd�I�f|��l�%�\�㘘�K�մiS77��@���&=�N�i ���w��l�ʗ���X. __t�˖�+�Ҡ��o�^�F��nJ�|�fݤQYEr�n�@��ؠZ�Ѭ��>'Q�W^��9�
E:�vSj�e+T([�|�k׾��`i'$����홁:A� 7�Zْ�U���'G�	��?�z�m:�L#�U�V�ʕ�js�����d;P��R�PK���Nx��]ҨQ��Ǐ�*U
�:+t�V�JU2��uB�D��-U���%��1��ν�x�ͫ�][���-j��E"���S<1bI�(Ķr�J���x
�e���;@f�Laaa�Ν�ׯ_�.]ڷo������I�&}������n`�-��o���X�n-��S�N�`���q	�
�&��s��:��CH3�[�Xjll<�70�m�R?��##AQ�\8h� R� ��T�Ɯ������+.<��oŋGg�.#��O���`}|��w#�>T�VԵo�>T�z#��~~>������j��Y5g� 	</����*�@��qO��� W��y�eoo���Fi޼y�E8  � ��aL�f�k�fE>@&r������a��A-Z� �����i>���c���	<��K������D�<��ԈK�G�j��H�Ӻn�:`t�7��@P��Z�:���_QA�6�gΜ9�믣ǌJ���߿��K)���G��"P��Rx�'����!)1�z� ��!0{����L{R�		{���b�g@!��Ƥ�WW�	j�S�>U��D
��i��&���Oh��_fEB��3y#�ݼK^JVA��H*׈�.P����Y$,C�Ӈ�·�nLɇ3++�lJ8٘�$�X��N�����n�f���@̙�Y>��4�
��f�����ъ�*�͂�����W�^��C�<�Y����f�(��v����@��С&\	Vx�(��t��;e!2�M�6��LK����!e�Dk׮�^�������3H��+Voߺł���䳱ԗ�����z��Ja�@ ��q[�-��2���
�7W�[	�_p:h��B�X������&�|�|�G�ѷo_-�w�blJa����r:��!`���|�����C��� WJN~�nBb
�%��Y2����3�R��<��_���l���U�_�P!`\�6�ҽ�s?a-�'W�\�h� k�Pd���3Yp�&<}j�Y�0qO˔)��s ��h|�ؚL�5j@��A(�����IO�:��A�A�bEϚ5/\t��S�o|�:u�ѣǇ:~�S*s����ѣn�ו+�ʖ�T:t("�b+��y�ܹs�v��U��=f����ׯ��O�
���_l��~���1�`,�k׆��T�R�:uN�8��9r���@?�q�/6l �� Q�gP����S�dڧ��߳B������ŋ���@j@(�9�v@߾��ţAl@-֌r\I���qӦM���ĉ��l+[�,h�F�4i<��(KC��<���i�^Xt��K�zy�=z��c|�]*V*߿z"(?C�+ؒ��X�M�./�Q���Z�9���5�jN���ʟ�u�����!��Rz�Y�))GN�� 2�c�jV��!�3O��7�XB��uƔ���u�$Y�L!ŋ�(QT���=x��k��YJ�F��A����� ��֭>2"�4'�|�Gh���\�{+Y�V�CB�$/ab;W�`_R��+�h�>��*�*�$�W副^�8�ɋ8�,.Y��4:v�)��A�y���{�c"�JB��O�|
����3��[LL++����L$�!'|}}!3 &�C:i�~6j�����\���ˏ���Z�J�aެ`�8��g�M�8\[�sx��R��O�~��^}z��b�Ě���*�wsu+T�p��yY�y����c�F�!���+V��6�� xt^����矵��%����o�H�����t�V�����6��;3�/]�� �0*j�M��L
��h�wo݊x�h��������s��
QE�!�,,�D��+�ϟ_�N-*e��up�Q�6�'��?����ɓq�il���gO�<z���ě:���6w���}2�V}C�F �@
z��H�V�l�nݺA6ԫW�cǎjE��b��]6o�N����J�"���%K��}���l���U̦M�� �!�+W����ԪU+ಮݻ�V�۽�nf��:ud�}�G�&��c�F^����kܸQ�^=x�@���'
x���bL�6mҾ}��f|���dފ�ɰf�X���{J�8�wﮧ�;����g�=\A�AA��i<�ޑ�
����*B}�]�4���O��Q�2c����m�+쥧�g/XI�R)o��Sʧ�T
�p���z���N�'�JP	�6�C;����i8<U�\�ļ�T�!R��� r���]C���6Ke��Dw)Q⣏>Rٽ�3�/F��%��왹��v��G�j9!k�S�)2�P�L�9=Z��D�$7�5���r��$���'>��7�&n��^?o޼���՞I�Y�(�����B��^�>}Z�!C��᫼dΧ(>�Y�Vu�	Y���� �O�:��A������{���[��M�4���M�>�"Y�2$%�nv���X�;����_�<��4C�͜9�+dO�*���B,]�v���5kF�m2�Y	�T�& ��[��add$1_�K�fPp0��i�f���Rxd#��Ŋ��ׯW�V�����L~�4� ��}/�ǧ�~Z�x�'��z-5�%��֭[���֭u�u�ָ"��ӧ���a^�<�(6&���x�ر9s�@r1�V*l�ܹ�C�jԬ	s��Թs�5j�ݳo�����(dt�ر͚5xZ�h�f�mw����In�'��>�.�(��o@@:�c.X����?� ��H�i��k,�����.@���,2P��C||��5kBCC1\��ɫ�>0k˖-A!4�kB���a��v�����?c�@�E��}(�JE�0�~����1��`��z����u�� �Q�&-wǗl!Kr�E�v�6�Ks���+�������<y���v:�R�#��/���|�U1��w�޾};&G@1�w��hgT��Ji-�N�I�!���S)���
�����㒔E��2�qt� @܄�Ia2p�D��J��d�`�M&�
[Q��M�Y5�u�,9���X}�Ԛ�4c6u�_�B�K��2mJ2�.��%�V�4q�\ϐ���[(��J)JH��U�����D�XK�/���ŘO|n�/�9�;w���qS�JZ�5o��mۖ,a�T֯__�P!:H�#e'��<�A���1ƤPΘ����"mپ�<�8ɚJ�s�������`�,-D�&իWwqf��B˖��񔈈�B��lxhxd2�EQ�5oo�1�X�ݻ�T(����:���/$'�jXz>�����֣���-���\�d��n�K=)��HѢXb1qO˖��r���D<��	N�n~����G+V�޽o?��L�ݸ9��o��ha�%�*W����22&/B�Rg��߻w�.m�SbZ���E���=��	&����E�:o���˖��Vkp+�
�����F�\۲e���7$��0�X1L��A�H���������Hi֜e��v�<J���w�1���PBK�,=bGI}�s�6.� �	�Dˉ��r��<�nn�I�Tb�ڍ�����n��/�pg�x2�=@���~��z�ҥ�߿O�.K�+�/]�4I���r�E{a����8c.�z��ܢǍ׭[7�Α�t�B�b�Xd9�i�k0Xi��F�	����#�,I���V���N������Ȓ*F����E���*��w�^ÆI�A���@��c�IV�3&rՁ�'l���� �{�9��:QM���u!�!i�Ur����L^�
LB��(�J1�q��+qX<�l�@�TX�Tk�[V
���7�B:�<b
��#������d%q�"�����ϔX�=G�-54���#�Eˇ��~�l��m)l!�r�o���#�FJ��I[V�GR܄T|Z�v;�49��l�ܘ/@���?���ޅ�<��/�C���ةq�իWc��<y�"U$+W�����q��]��\�R�R�e˖�s��!�)��'�6d��:���x�	��M�J��Su��Փx����*���wޱ+m�8#gy����ҨQ#��II4�˖/Ӥ�`͔_��3ƏO1�8���]�xQ��DA3f�x���=��q��i��������@ܞ8qr?�]��j�j����C�������K� }p!��m^�P %9��8�x)p�j�i��ݷo�ٯ_���.RJ����Ϥ�J���*���&n�[]U*gp��7oR�y(�i<Y=�#p�jժ)Y�#����	�#� ��H�ױ��a�Bj&�F�w�={�{�7p���˗����"E������.]
���~/7���ڶ��c�K�H��&rb�|�� ��̙���9�s�e��\i]�9�qER�H	�i^^�W�^�k~��'���T���e�5��D�ZC�����Z���'+�D,�ۧO_�bIr��s�7��Z@G�	����r8�k��P�Wb\HJ=_8п���-'�s#��Mib"�_4� B��Ot\� �PAg$� ,"��L9��$�ƫ��%�TTd����Y�zm�re1Vtgab�uK'�h��2�=��Be3lܠ"�t�߄���T&R��x!��
!*�WC�<8��� -h��k�S�uH���dw�G�j�8Nϥ���H`,�9��#8��Rb'��W�t9O��ݓ��9�j�/�!�7o�	f
�x�ڵ��H�4hW@��!<���ޗ���趨IY�$[ɖ䇾�
�'|,�9Y%Y��$���<�el�v!�Sy�+|P�*(F�/��8I<���~�
	�x�v������gv�7¯���D���R�KSR9(���`������8>�+;	�>}��%JI<M� ��k�2�Ν;׶m[9w�j%x:ϓxo۶�K�>�;�Z��+�+V�:t�uѢE�����=�`�^�T�dI(��5`@3�/ݸq������}#O���TI0���B�
�4@N��=z� ��ѽ;d�m� S,��)�D�/ W���l�e"-�f�#ց�M�8�T�R�|�����Xiӄ��B���bm������r2=v�����ݻ7�Q�ց��{<ȝ�J�%��63iue˖�s'lʔ�ܖ��tt����ӓR2$&�~��2��V�=��t�`h2�Gh��-@�O��}�)�����\�x���}��V/j7�y�qH��ٳV�`4���������1虥�k�*s�T�~��}ҤIo4n��)y5�ӫ���������P�l˘ �8N&�I@"9Z�C!�Yt�P혐�����f9���t���'����ْ,xF�tʭ8b1K���l�G�q{ۉ����.�VX��bp�υ,�7�W�{�j'�C�L.���5�N��ANP�22��Q�P��N�_�`A��|�����uG�Z~; �O��W���x��$��>=[�e�"I�_~?�R ��={9rDi����W��*��Q���BZ@Y��s�k�����W�reI��l� ,��+�ӑ����'n5`��������ۀ���"|{
�@@˖-���*��Y�f�u�ҥF�P�\�����9s��wߝ;w.�|���Ο]�dɄ	yyzQr�Tc�h�EK RǋT�Xh��fU
�
���ʛ�|H�Ga��[�p!�:�h��-�$%0`2Zk�[x�D,X�X��Q��D�%Lw��Q�J.�Ր&Ѳe�0�B�
~��׬+7����bk|�Y�A�-����G�����%51C�y�חK}���N�Ov�x��;]��&h�������Q�>�RN�.�=�������ל������/��S,X�@�F?�	S�:��g�y�B��w��V,��qq��j��Iƛy5 �%C�گ�������Mtn�������d�s�ߜ�>�1#QD8�b�Q�7����3k�s�⹄B �v6:�匒ޑwOMV���q7^�G-k�|��#�?�y�H��U�,E����ۤH@`�����_�'�Y5]A��ZD�E �����%�H�\;b�h�իW�����W�N�!C�4i��uO����˖-�̾v�F�p�-_��m׮]�A]�MqêU����>���a4�h�,`�<>!�RPЌ��x�w��kT�R����+W�ܽ{���d��o5�F�Ŗ������S��yV�B�7�|���eg���H�7�R��&'��\_g�;�Kł~-z���G$'��lZ��8�G_@a�̏7e�&
E�I��,�������h�$�uj����UT��ORf�#���_k��g��/�M��������O!VV�S����r��v��Ќ_�)%��Ȝ@>�F��}E�p�ː���n5j4lذ�;f���摶rِ����h_�~�^��]�x��Na+��l:I5�|r�;S����cݍ�����(����(���˃Qܣ$�p�����ٮD7ww;�2��M�>�
C'���ih�ȗ�U��e(��TQ�~�y_�,t;���R*!�EZ=Q�B�i#�ןը�stlѢ�=y%1�<�>��s������>�<*T�Dɒ5k�)`W�0o��|T�W0` Y���{zz�
$^"�^V� �ᠵ�,�d�fP^�!��a )^�y��7n�X0�ۈ�|���!mX`H � �jժU�vm��rr'|yc�̜(�FC͚5�ǤR�$3!�C*�Fh0���!�05����;����F��a��\b�[�2f,ﲓӥ�,%I� �/��5j t;�_�|��Ȑ�Bޙ���,,�_�k�!��Ҽzi'zD�Sِ��"|!-����p�b�����~Ra��Xf�C�cG�u�,�Ś��b�nP�_�\��pg�.�"�{�#v���m``�P�8A�i��fq<� 1t�_%C����Ϛ5c8a��ɤq�
��ܟ��ځ�'oݺ%�4E�#*���p�I���yr6ۼ�!h�)�W���R�{It�Ty);��B_	4��lG̉7�Y�z�*�H��W�\�jKޯ111����\����"E�0@��]�QH2/I� p"$ �Z�F�qz�3Y�i���/ �BBB��`����:9yz������ǂ�|��
x��:�9i�`pqq�Hs�'�(Q��s%�'������g��U+��YhUaVkU��^իw����+����y>nH'��*�*���//Ve �i��;�-�W�x��0�.z@�!%2���ꫯR��j��t�M�=�t�9[�%�۠����p�t�a@�%o�`��F���\Zޥ�����sQ�����ײ)$�&R�(�Y�;.��.�-�[���d���M`$,�B����-��2�?~��?f����׮��xw��R�%VN�.@��R�X������ �?��� ����H��b�O�>=z�h ��'���޿��Ƀ��޽�K���cy�02zS~#Oll�(HR�.�7.p$�m&-��$`��y��)���\���\��,g���{��1�`���HL���N������,ւ�V!�	I(��aΘ�;��ŅP�޻t+�)�&-v�$��7��v�U����ˋeF� ��+��#?������� ������ݘ�b2gl���Q�NS�థ�v�R�(QTa*����*̼(<K� c#�sj���"(c�KX���t˷n����O5EXeP����M��/=։�-"m�Yqv��BV��ܢ�;w�@�yt)�I�m1ϼ���`��Tv��m�%�]�_m��JE>mc��$� �*���e�7�|��I�6�)�m�J�+J\6T�T)o�ɯ��|y�@��X��r�P�x��w���E�l�*4y��@�t[|�B�0�]!��hY�ݔ��h���b�� �8��R4Э�&�3��fL�a��j5�HDyV��(C��6��e�qvv��xxxA���,��<=�g�R�ƶW�.��ٙ�C����E˳;p?|�
T�1�~`Sr�e�z���TY˅����듌��.9�'D(��ެ��R�.�_���"er��x��_��&[Ͷ��3� &�9����R�M^o���[��"y���o�V��1cF�z����K�\�8�Zr��k�H�P�m���J�����:+�`SH�Ņ�%Ĭ���LM/��;��IY1��:v[Tr���#����"K��9K��-ᶖ��_�;������h���s�Z�	,��lf���$�L\�+1�z�S�-��9陗����Ȃ�,
fq㥢S��R�yf@�;�q\KSh�F��
b�'�Z��YV8���KX�xq�m#���c����;w�(x���,�+�l��������'/�k���N�M�ij��D�J!����11n^O���|��_�
�����I:�T�GD���:Zi]�p��\���$����?n2�=9��Zr�Wf^V@��e|�"7���9o¢rvu��(��V��]�m�`���k�:�o���K�K�F����)����Y�s���SU�Qc�`��_Z�g6��e��6%���&�|����#t&�JiH�w��>�g��t����A�L�5�ݲ�͵��>*2�A� �Kj����?�O%^:!?XK&�ڬ�i)��<���RR�{0㊃�F��Z�/]i�H�.�ց��f �q/..�����F	�LeN3e��Ls��#�_�M��4��-�Y:�!��9�k׮m۶��d�����X=�L&�>22���Ònv���Vg�6�_��M)���(�w4�"�j��&��+}0�(�����5�"����J��?�+���L�&t�v�I/��Ǣ�(��3O#HE�u.�\B�٢
��#�+���P�����<CקT���^j�#�G��ٳ�V�R��o巽��9k��6�ѣ��Ǉ��U�\���e+�cI��A�3.\X�tPj�f�Z�$/��Y?%�������h2Y����5��l�C���+��"�E��x�/�] �ټ˫r5�ecD�Ѩi�_P��I���T�s!��y�msb��G�\x>��!�ͫo��Q���ȫ7%⹇T�oF�s������@ze�R%��F$�"RD�q�N��s����7��,[�\��&��ʕ+k׮M��D-�_��茝�˫l�#NNv�324`k�/kc���"	���^R8T���f��꠳Wd�'S{�~$�<�nyMԍ̱�������nY^�f�4{�XZz>E_4K���r�WA?�P��5B'�Ck����x������*�)�������F̈�qZ1>��&����Km�˃*�����n۶�C�N�7&ĭ��]�x�;n����J�KHH0�,}�SO��4V8�͂��6���X�u�e�[����={���<����B��ڿo����1��;w���6�<kܧ�E����jE�=�tЪ�3�'�Ŕ����{����[��y�@<��]�v��})c]Jr�a��}�݊+>��B��`��h�14��F�yZ�3�Ɍ�P�4QJ��Ϛ�_��\B���skFM�HyeR_4�Ó�C��G�Ϛ5�Q�F����MÂ��uԞ���f T�O4�*��,j�,�In���}ٺ��V鄾B�HLL�?��o�5j4z�� �	�{�����_�U�F�&M�xaO��b{E�Z�G[xx��˗1顡��^^r���k���Kf�T�xq�0�������9 �҄	�w�N��ɓ?��Ӏ^8��w=I@��.f��4(�w)�`����P�$e-����J=��eQf��ӌ�J�R[]�m>կ�YlU�_���#.�~IL���-R8�P�BG�]�p�СC��1)���y	�������a5R*V���ח�����1-�b�I>�/t�7����S ��O����j�
		�y��Ν;!����M�Ο� �W ��%JH9�U��]z��l�.]�ݻ7�~���#F��ˬ��A���� Bjڢ����?��G/9��H.[��Ν;%J��׭[���*���,6A-TΎj7���"�_`��l����VT�Ai�z�)lE��o_�e4�N�J��W [�b�Fv����3gv�҅I}�[���9*�f[�\����+��We��K�p�=w��߱ce�.�,e������U�jUQ��6����|�E�_��(���5m���M&�1��&qO�8;;���ӧ�BB����S�����d��?�GI�iݺu}||nܸ����bH}a�O3>�jH�R�J�z��5��o���fއ4{��R�v���`f�V��v6o�<~�x��ׯ�2e
�9�����gΜٷoߕ+W([���,W��Jշ�����F�4^b���c��Չ~fcR���<P���y�qA����o'&b��%�E��`-��2Wx5+���,��+4wxKNI.]��+�tl�o��I�&�_�@�%(�Oc�<a�
����"m5�^����f�\���￧��+��l����k�n~�����+*h0�^\���vo���9��G@���ڵ[0~DDıc�4h��6�9?��#~/[�,%(��/t����?_-�<6��\�I�z���նm�Y�f�Z�j�ȑ�U��O�:u��e������|������%b�W`���<�Fp\`G�"���޻w��'O�f��ޫW��k׎�0��T�6m�\�Gy��Žq��`��LL�ԩS!�����P���/��3&,,lȐ!'N��^0�$J)��HY�_َ ��*>�W@I��&�0%SV?I�����#3���'�K.lw_a3��M/����*!ig����.]ڶm�u��5���SSS�ח��2�ڄ6Om�ʕT?��`q�,)�����Q(�l�Z�̡�%��@�Wn���'Z��N%w�א��� ����Fo�A�㏋O�<	�NU�p�9��l�l�/����U򺨂�۹�w��a��٠�'Nt��I�j��Eb���y=+�n�[�WV�f��r�O9�o��:�2>44+����d4�l�r�ܹ���v��Y�n�g�V��3��̙3,X�u�V��4���-&&
��c�M�,��{�3�s�[suUW��t7͠J�Q�8�S�y������8�SC$����ט�D"N
��@�"4�� M�s���=��ڿsv���F�y���r��s����k���k �>��S˖-�������aT���Z,@WQ�H4cƌ�����@��׈Tt6��^r�4� ���V�4B�>��hb���1;��j����_�\s͏�����m؄�f�Y*�xL5m�f
ϳ�l\��.�h��X�x�Z��_�d�}gzLk��)�D��PQs�b%���烫�z����~�6�W����Y���fͼ��&�~�zv,��ˬ�d�/RRF$�XL��}ʪ��̇�x�ݿx��J�*~�������sϝI��[4[��{h�~ަ���U�N��h_�v���������W��7��q�g�\��3��̣�>�7�7���C��_����������}��_��?�S�n����Q���IђT ���k��Q�i��G7�㉆�j���7��cX�`�2����0��2�S�\]
%�,q�u���}��'�X�s�NC�1I���gUU��t�Y�E>F
E��Ϸ�,�71���6Rڔ�?:�-�����
��R��������k�>{td���E:�X�r���ǌ�im��҆��
��@P
���������T�Q"A3�d&�y����O<�D)���c�yf��]�v��׿����ͼR�U;/�����+����7��x��u˖�N;"��+�`Y�?���s��:������G�c��+�͛���}�}�{�����3�<J�iÆ��v�qDM��}�~<Ǚ亮�:ԏ��*�J}�*��B71"E��?Z���1�S��(�lVI�nE��g��R_�y�]S�:p��~�����7gϞ��؈�O랙�Ƚ��b(��/h�e=�*v][�&Z�Οe���ox�.��\�ijcuӕʦ�n4�H��o���lc��^�z5��9眙3; ��nH���~��T*_&^��;��6����p�nĚ7�B�,�Z*Ł\#f����
RϞ=O>��Y�q�;�(W�V�X�n���/}���Ȇy=Լ9s������s�r�nY^xa6�~�;�����_a�%���'����mZ�G�ڴ=�������w]t�����hn�@F���L߄I���B�H��PR�����mV�����C�ï��n����
��/G�UZ��۷����fv����N`ǖ�R�u��Dxztd��j'^��~j�b��k���~�}�v �M[�Lk�0��zn�Çoܸ�G�x�5�	��TR���;���r��\p�1m��V�kX���D��h��S@���G-Z�!ϙ;���}�m�� �>~�u�V��t:���6=ld�D ˷�T��Qbee�����i�A��]�v钅�m�x��gc������Λ�B6:x�d�J��GR)�=��$zR����L)3g���w���-����W���عs'��j�s�>�LV*_��W���7���8�3h��E܏t�����3��|���/�y�6���XM��I�O@&�?��ոJ��
2����w����uuJ����y����K�~���r'󣶗�\�Pij�z�)���=���g>�3�K��J���Gۼy���/��Mozv&U�j%Oo�����7�NSs�x�Ϲ��[dL����r�\0�������n��ttz/��H}0�;�3p^��+��xu�c��t��===@�---�=��޽{��>x��/_����N(�0'���w�u��>�1hc[�lɤ�]v����YS��J?�Ղ*p/SF�� F�\^*��P'bW]}5��7;6-���+��rpp0��8d�jR�φ0��]w���o���?��T���ۿ��>��)Ot�Fv� a~!�=Hu�EH}}��G�?�M�d���J�X�����}n��x2U(�\[r$�j.���?�a�-2)�ejۉ�v��>�Ԝnl|�[����Ȳ��4'�B�imPs���h�|����-�S]�奏�V}�A�]����/}����,�u����wպu�:;g:t�ӟ���={
�ҵ�^Ka_-��)���"xx���}�O�SlO60���>84��������]t������mۆ}N?�����_�܆��%|���*B4?6F�����?ml���ѽ"��ޏ|�#��ຌ�?��;���1�xGG�3<g�C����������{����#��_�҃�imm=|���_S�іńD4�a�R$F	ݬ�*�z�aV/�_��3���ŕ"��ze��'��!�
-�����w��P�3�O29e�8'-��C�2�G/r�e|����3eP��{��Pr�=��Ys>r�G�F��a�̺e����=ys�X
�娧O_Oo{k��o5=W(��ؙ���li�ρ��g�}��tr�����z�ܐ�O�g�����I:����ɋ;PpbPLA/vt��x�'_7���b��3�x�O����}+�Z[k۫�<��J$ғWaJ�mh`PLG�k�n}!������!u�~��� ���<��nh�N�n�N6��k'�z�ŋ���rյ�q���?}G<���zu䮜�[�T+�X�>��O^�ҙE��\��\����ۭ��B����rćz�44dU!��O(������o�t�M�l�^�&��A}���/���?�0��'?���&�s�.Z���V+Ɇ�1�}���-�J�?4LK���:l���Iʑ��KA�D���B1�FT��Q����j��*m���㪌�[���c\�����~��w�Ws�ҥP�8pꩧ��Ŕ؃�p�ڵ�jӦMر��Q3����qW�>'ҎF��o}��o���` �b2��������8w޼���Q�pO�$`�/�����<��_�mllR���<.x���_��v����7��T]*��~��pe�VM8	�����:��n�o��S����cS͎��������W�Zu�ik���a455����ݻ�p��"R�44~�fl(��a����fE\�߿?׉%��?s�-�d�`_lnn�_��ls\ �9�ëU�	"��/�/:
�x��Y~����Q�珙X��c{)M�������K\�̚O�7�i���G��Y�`�?��?�}FONG�N�7yG�X�C�F�!���H9o�:t����'
� �K:|(�JCaJ��?�G���	�g��/}	�	#��]�b���|��e�/��[n�"
T�p��5k�Ny�^�'�T�,������;::x�h?��?��?����������T*	9�ɼ��K<UY�79|�����~�|�\���O|�˗/Q�����I�����Ѧ������=��G]�d	�.6;�
�m@��^��o����C�(�&0�YX�C�87Bs�>����haO�s�������~c�^K��&��|������?�>)���ӑ#��E~�PHg�" �'ӱp'�`����5k����ba�炆��KO9����/S[�x�u�]w�w�^��=w��1��;QB�j��g>�E�M�K���k^������l*}�&�0�)l�\/l�8L �'�>4�m۶�衳�p�嶶����'g�y&��|��w�}��e�U��@�̙3�V'�Yռ�����Gg���S�{�_��?4�\��#"l߾�3�������C�wwwg[�x1�ҧP�הm��u�i�7ot������?�:<_����Ej�Hz|)�4Lۂ�w=Aa��cŞo1�(z4�"�T�5ۉy�oM�8�m�������*�u��v����Vs��	�Ŗ��W���G��5��ɣ�J�
�^�^j ��:i_�����g�C{kik�ʙ?�� �=9\��|5d��O0�E�A���I����m��6�#*d������K��Ȥ+���0�ʿҥ>����7n���w��?�������_���^�l9�ӂ���o.^���|�_VBCR�A�����v4�hǩG9�����<��3g��_�����g?�v�Z���3�O�k:��>�e}�7�?�	���9����tO������6
E���e�eu����dUGM�r��;2c�T���w<�1h��ei,��f����3��7f{{����%�v��.����Ə��@���7_�����I��)_�)��+9��X,A���r���'W�\y�G>������fAQƇа�T^,��:��^��W�q�7�tS�����9�xC��N���qNё������O����5���A���t���ɳ�s ����iY��S�����x�{A�����	(&�?���l�w:ɠ�I�m��<�M��bg��o�vݑ#:r�졹�&�<a���i/o@g���Y�sJ�t�(AJ�=Cy�c��֤S3�n����x���R1�Nm�^ќB������;wn[[�駟����wuvͩW��C=c#��XqƌF,�U�+��ڵc���0İ��R��R)��OR�ٴ�0b�?zOh29
8�c��~F��"5H�5���ށ�ƖV1䨯e�|O�����sxhh˖-)��q�l
��0F�̑�_s��s ��v��0)����	�&e;��»�t�xNq<�#'�:�aB�R{~�ݴ6Mc�1M�?s��\㭖��LZ��j�?Zj�Z��N��7^���Yڹs�M�֬Y��l۶m�b���ի�MM�� H��ފ�y�0�֎��*\���쎎ۑ�N���N�14-�=/\�} ��&���׿��h�)�|F8�W �1p�(���ݻ0�����fGbO�yL+��R)|N�b #&�0�4�\c���!J˄�,G��G��и]�1�
�qD)eݘՀ��P(�PXI�Dl(:����O��� �)hb�w�f` ���B&r7��Fd�k�fh!z�U�{�Zgg��_|���g�zڧJ�Ǵ@����(+u$�?ӧ���2�S�ab� ��=%^y<枯���|69�2���;�`-t�)y���(�y���Y�O��n��r`PW_}5�5w~��}�n�W{��mlnjhj�4>���;w��曋��E��\��~�+,����!�q��1<�u{�9�T�N_�{��_�ҩ�����-��-G�M�L쥯r�3��\�����c�
����[ч���x�����-$�4�b#��^11�/��P(�y%�ѕ�Y�D�^C����ʣ3���^���*�o�?�����G2x�hH�G�F��H�A�o���O��~TxtB�!щVm� 'XcHf_Q�G�>����3��K �*)2���������ãw��1c��t>f�'�"Js�&D����ږ�N�?:œ��+\8���d������JS�q���,�:?�q4���������0��+���9֦���C�����통Ϋxc�k+�`{~�6�j�<dr��WBۼy�����O|�7�p������������?�A��?p��_��E]��O����ݼy����7�s9H�|������<���x�v�{5a�L��$�1/K��jPMg(���0�O�@������B����eɠy>>k(�����aɑ�x���o]�2zϣ�c1��D�v?
H3�~5��~����!��@߲�F(�)�Hv�2|��%"�����rQ�h�-QK}�T#��R@r]�6�?R>�q"s�b��A3�Ư�r����輱�J4"_�DS�^�����F<:���#FFF�.�F �
�3´����mUކ��Ohv�����`nq���o��8��O|��[�!sZq�찱o�-	�˪Ͽ����Q�o�^m���o5�qfH��h�=t�e���Τ"�?����W�����X;��j��pbD�s�����Ȕ�����,^���0�>�u�z���馭[zz�W�|�ʓV�����n������ןw뭷��Η��A��V�(�JW]u�>����r'z�}�;��\�1ş�
�G6��'�P˴���d޲������jy����g`L�hL�MC�ܧ���k�kD�U�Za})4}$/�۸������Jv6�M�K:���D{|h�;<���@��TC�q�>�2ì�'x��D��z	�P�]�6*3�'��4�XD�O��>�""�}0¤~x�!%(�#jf<2U��6�Y����:w�����/3"{/��k�=��.���V� >�"9��'�!Y�T�1cƒ%K�x�	G��.�J����^��p�ŵ6z�j/�>�؍6��=������=�9��2���q�č��W�߸W\O#���'r���r�g�[���On�����I����E��!�J� ����>r�j�8i5:��lMSh��W�\	:7NT��"	�H�dȘsP;���˩��n�u�{����IK,ρ���~�����o�u�xG]ѡ.���ׇ�N?�h�7nW:�s &Yw���R���v�{�DŢ)@�����?�C��<x�� ��ɾ���L7�<g�W�ՙ3gJ�Q��F�r�@� ��Z��ɺf%�*;lDt ���q�h�Ä��2�Ro�4T�@ʤRR���
W*��ټ��`�|j��i6��-?�<rƣj��H��a�~`�'��񙃁��n=��R_��X�XTW�d�Ԝd᧴�
	݈E�:(?Lg3պL�!��-��{��xv���u��i����&�D�FIj�J�r)j��x��%l:��3��i/����?*����[g��Cӈ����M��IF�Vɍ"�ڥ��>�$R�Xb9>�C?q� ]A]n�����ҞZ�[4j��q[N��N���GQNT��%A�"�xR���ǜ����'�VM�i���u���7��p&��J�M�=-B	���T�ڎ@#)fd$S ��۷c��p��븾[��2A����ޒ��4��56�A�)��~$o�Ck���#Z�섦Zȸ�5�
s�K�7,��ݣ�
c���	|�;��w���_ܯR�L*��CS
Ͽ�݌|�74�1��!+��q�kC �LŒ�v����P�%}�ߦJO�
r����&����=�x���J�Y�L��0�6���`���;u0:o�B��z����u$>p=�R)3���5ͦ��"�*����|>?�7o���:��7�10쁴��B�?<<l(� ��q�aK@����JO�9FF Bήe<�f��I6�[�Ta����~,9�|SS�Yg��b�
tUpM&��[UP�V��'o���Fz��S�=P�F�!�ܨN��jУO��ځ�m�f�QL�D�Gi��y64r��z�Sm�ࠢ��"S)H>�K$>�kV�V�
�����V�QhD6���IS�����5|��Sۢ�'V�bcb���F�����v���E��E�v ��D;�&�@���F�����e~�Dȟ+[���Ħ��^/��=�n�����s\�OUQ&���)��h��R)�t�g,l�� ��A:���$낞m�
��X�ctt���Q;�[ks�n���4��U5s�ҳ������G-[�O��I���L[��h��T��=e0�{oo�ҥK��ك��A�����|b �uq�R=�̧oe�S�W���|��`2����e�T�t��{`�ZUm� �
ìK�?жʣ"z�D9Ƅ��*g#+�jRv5?@���u���CCC���U.�����[έ���r��������a*~�7�&K
����1�~}"%�h��Hm�e=M�C'3Z��	�yCC:�9�8�02�)7�ogg'v�����I44*r�<�N�FU��������NN(-��ĆO�GF���C/9�nܸ����{�l͜9s�ܹ|���d��fx���}д6�U�I���"�CZt�[�ʄ���訯G�=Y(��5 2�c#���T@���S-c0?�s}/4������L��[۩��=�Dk�P,�����$Bs�v��'*�zPF��"�H�<=��5d1�Ch?4���0F�+�D�y�7�a�]k�-���N8�(�r����*���l�JU��TsIޓd��@9��>گ�`E,d�8�PÏ����Za�Ht*�l�wӸ��n��)�$fǽ�#M`,Y�O�-e���q����5�i��f��ǁGG���,��1�� ��]5Ms�F�7��G܃�&'��m��
۳�ZC.ǧS��[|H/WZD�s��G�%C����1fx��b+yJe�WI'b;x����5�(@$Z�ީx:8�EW\V�?R�ת�C�64�ǲ�>�@��Ҵ`��ٳg��]1H8��(P�X�� �{KE���I}Ck�iD�Q��#_�}�4�y���V�i�U�Y�w"uL�6��J �b��J�h��k��]3��c�xU�l^ı�S�D��H�I�f���7̘�V(Wd����{�ʍ/^�(ƊR��E�[� ��dt��y�V����PS#L�jC4��r�]v�I'���l\p�b߾}�{/4-���D�"Y��QR�ǜfXsIo	
Z�R�VA�//�L���4#�M/���m�O֣7��՛�o������0.��hM9�}����	�2q��|�ZC�O�&��3B!*��HjK���1|[�Vh��q�(ʘIHB^� `�a�8�RGx�����0%�~,4�7쪯���!�9c��4�2���yx��N
t&/7�4U5U/<U�x�:.��� ږe0�0BN�5�&-M$d�Z���D�a�D"	���C�D�"�Ո@��R�>:F���^��4�k�N종\t�`����"{-�u���O-�I*~h\�D5�\�=kA
�/��Z��ڒās��+:oj��	@�'M��Ԯ-$l�#Ѥ���R�~��X�K��)W:ؾ�1 |�1����r�i��J�(;�"_��
u}���k>�X��RA���>��
�h�eD����D�Bm U?*�� �aCH�z}5�d�1yQ��@C�n1FX��y�0K�򻣣��g�`P��9�>M���b���7<�'|ŝp��`r�����9�d��=���E��N����5o��&S6i�k�^�f]|���A�g̘�#|�����<��78�T�a�h��|�Ȧ��$h��d�p�ڄtB���Gj�O��?X(�.�𢮮.�xss�s�=G���ܶA7��Qkd�TQ:��m�T��Ǚ^�W�T�~tlP�T�2�L���(�P.56I@#htѢE�
mA��7�4�r�Z�v��=V�T(OZ�_���@��[+�56�,���@���-���J����pǃ |L�1����bl(�R
�&'��>�pcC�{K�(ϬU�o�aO��x�=f:q�^
 ٴ��z5�U(��n�4tY��:�㘎�1Tݒ�
�[��U1/����W�e.�X�q���`�p�|~�����KX��a�w�L�`HA+�y}�q;`�U�\� �^`T.	� �+����g�Z�niǮ�ʶ/�B�Z�rR�\C�"bˉ����=����0�)���ۡZ+�#f�:mL̐c[������~),�D�����Q��n�?�W + ^n6�V��{��L�`@�.V�Yn�({P�Q�)@+�ah#��3�uaw����plύ'�����w�mZq����Z�)n@�o�n�jۖ �����/�f�ؚ�&P��M$�3:�p�LR%�	�B�@d?��<�M��Mr�Ki�����o� ��n=�ĺ:;�,�$�k����tCF�:��%��N�G�m\PQ��즸/�TĜ�X�t:��:��
�S��D���%./e�n�b��l"�����`�#CC�}�3gv�/C����X2�)�FG����R/ȶ-�;��A�,>W�e�3c�oE
�k�6�D��ox0Ր/�f�X%+pP1-�����u׬֤Z����L��x�-�i"����3j�j��.V7�����ޞHg��Zf*+���C�f��x��4SdP#Aʩ�ft�~���(p�J��)��d�����s���X�ּ�l�:��%��|	2�qñ�RSc[ss3g�R�k�\If��tww�+\@�)�z���,��Ρ�!��d�� ��B�UA9�2xO�C*�AWk��]�Jq:�I$����*uO�:�J�0�C��ϔ]\��Wh�*��lh��A��ض�{���`���])�&�m�GOO��O���Z����(�xt��q��Mb��M̑ƹl��}@i6-om:�O�~#<3��(��1� ��Z�qO���,˫��u�!��JJ}�:[����a׉XR=���w�v=��x.Hr�i�������-B�;��SI1��UJ)�yǎ���t������C��Qg��菪�@���E��,)`\LU��f���,��^���DqR��B�M�ik��L�*�����0M���5\�E=�á���bW�BgpL`c������i�vW2Yl?�Rp��"�;�WG��x��#&5���-����L$�^ZG�h+��
����4�������1���;ZڨV�����g���ǨE1J��F$��5��ۜ	�0BrTM�)˄:!	�M͊G�D�ŊR���P&�U���k�V-���vP\���`^J�X�R��Y��@���*y����.G[�Z3����D�ݪ�0
ƈ�~yz��8�0� [���]��YǊ���*�U&Gy6@8�<�2�k}e���[?��'.��6��|e��:=�]|���U�Q:#�����I���3#[���̕M���CZepm�����B�� ƕ��x���>AX�G����X-�M�tw�'�� d�Vz�,n��0s�5[�w�2��A�+��<��8n�,����)�@T�;p|��}�L0���Y��D�~\5�Hd����Ib|���d/��\�Zu�j�KA�[�����㚡��(s5ɓ�Τ�D���9^Ѭ<�_ϗ}�*9�r츚F	�on��㗿���MO�󧭖ھv2������X��?#o��T�ǱzF�����z�cI�cI�c}�G�&]��觀?�Ν��Q��Oh��t[�/�S��˗��j�*�L�[����/������v�{(O
������[7���`�=�S��DR)Uc�u�S�B����:$
McN��1Se*�q���V���\=�xHj�6�>A�|k<�K����y�/��]���X����z	�̠Q}f�"Q���M1G��V�T��e����Z��Ҧ,��CK1?�E�~^AW@-�:�ŝ�C�7�w�&T�e�$���2�4iD�m�f�eU�LdԊ�G��6��y�GMV�Z �N�Ov8�D�����4㶀ojo�|���j�h6ti���k�����u�"_շ���f�~�� �:�&gZ���CZ��$���E�损�!�(U8��Sf�>WJ6�1Oa9���o����RnE�����=7Ȝ��%8z��*�@�n�xz��J�q��!B�|���+��}�}ʣ��7�`�I�"����Z)	���x�e�mx1q�c���sL ��Ƞm�ô�c��SxUh�)������Z�5e{Ckjh��Wd,"*�c�T2�z�ݗ�����p��A�t�9�����z�k�6���L���A�Փ`J�/p�b�FV��ztڕ;���f���wD���s����X�� ���S�I�F/�q��O�XZ{IzK����1'I.Z��KeG=7[S�cd�>�^���@�K��<�"a%���Gyà'&�¬�_Ǐ�0骐VP��bI�R�1/��З3
�)4�)	��Mcc3�}�lrF��d2��T�N�i�H3�d�;P�������I^s<�,���c�cf��&�\��E�ȋ����v����w,�կ~�ܮ���޲�Oe�y�<��{��>w8�Eѽ7a>o�����y]�9֡�q��=!aiBZ��l���z�g�v�*GԞ�e����oݿ����.������3gΜJ�|��fNz��q``��uƺu�N>yuk+�Q�B�
)����۾c'TI�x�6)����r18��MGz��b6�h�((�jJ~lP�Iu�k��
 G|�}�E��e�vb.�5Kb/�`�zH�ܹ|���]�c�s�?B�G굶��'K�,A�<�Ndi�ß�����Q݈�xX���ƚJ��b�si�ey���f]s�����R
�W�0	 ����^�~��L�`o� 5��TN��+5F���iE���g�\:�Ϟ�P1�?����ƴ1#1n(���=���G4#48c5���nh>.R_?�1��B�N_�r���QMuLa����T9?�2����+Ϗ��J�4u�-Z*�	�ɵ�I��0���X�$�>i�OB9�����ɔ����-j�ji�H�����|u[AO�8���j9̫��a���9���>�hN�
w+W+Z����c^lmQ.OH���(EB��P�}���e%2|P����BG��*�T�fU�si�����#�6�t��Ko��Dm��hU��/�;��H�y^�f��oR�&j4���P�:;���t�.~��B.A���wB4�J�2�N�0,����Chn�p�L68� t �iii��6�/�q�
���h!SH+�H4����F���EZ-�I`M�$KO�����#e�@��-_���1�����������g�s-3�)u�y���կS�\�8����J�imZ�'�8j{)���,��[&��[�=���X��)%'�֊+����z��o��;::zz��Z��%��w����.�H�|6��B������o�}�3�%� ?v���d29R*h�U�9Չ�_�l�C=t����3gBd2^yt�W��ߝXJ�]B�>��ͱ�:q<i��~R�>��,�?��矯�,XΎ�ժ����� ����������1��R�����M&�#�rˌ�o Yc�Ѩ���υΘ�Y�>|x���L,��2�kaI�l��:��+�kQ��dO:Ѭ�T����5ˉ�(<q��9|Pv~LS���=��31��
��r���#Ε�I.רUs�I'���G��6:��GB�(ڥ��)G#��`����ʵ��^��!��[��!�*���;�U8n�S���j��W:���e�uW�q��7�(��%ӫ�r���M�2f�2>z<-�[�G�|��6��q\ ���+0�R����������
[�L����X�b��C�՚W�Ts��eE⍣bO���yY5��Ols< ��ᡇb���lnN������I|��Pb�p�T�l�!q��5�v�����b�r��Z�1���Uԫ&�T�8��B�1�am �,��1�Zg%��:AѨ��D�x���2E�b:���/�-L���Z���J�mT�-e4�--�K�x��x��č��b)��@������j��_�@5 Q����|	l��؁���j^:D`�K)�k�
�r��K_W'�Ȥ�dB��X�II'���u�Ig,5<,��g����F

�Iy��SVCT� �c���5H��m�4{gv�A���V����͝�M���.���T~��
/灝q��I�I��� ��N����w���L����$�vt����O_p��W���w�͵������k�/�t�,ׯZ���-��L\�*��~׭��������A�����>��.ӧ��R�W��o�B�X �̝�k�����g��:�>-��#Z�?��	�����ͧ>�)LŤ>C��@�h����ַ�u�]wa~�;��뮻�Rv��o<���d*�h�\&�*��t#\VfP'�noo�������S�А޳g����|��ݻw��dY��T7caF��kȵ��Q㬇�xj���U�|��3 V����"�?���߿?�L:th�Mb�M$�����Z��;���W3������I;���h W4�RZf`�� ��DUXv�n�i��mFtnJ}P��	��,��_�͠aF?�/KLTC��E��y�ҘE"�d��J��Q�+O�qgðI�E���	6�ƪ ���'Iwm���!�?4���A�F������mߊ$�r�I}g^�z���h�Xb`��)���m��T7�F�����hw���H-/L6���D���L]��{����dJ��L(�����E'�3vpW)�� 8����PuV-�x^��̳���l*J�� c*"?��\�&�j��c^4K����l�X=K�{#L��M����)
<���_�B4k7/�9.���1C�Rߥ)Q���.����դ3��}���s^6�r�О1z����	wq�֡������m�B����������<�W�N�����;o��bH��4�����Jf�Y�L��`��Ym��I��̞n�}�-r*�N��L%3�ʈ�Zu9�4�lٺv���N;Ӛ�f��Z�:�Q�n�$_ B1��*fWY�����G�}�����W���֭�\���ƹ�VF�^2I�@�f4���X���������p�X�5k&� �Ic.��;(�|L��a��s��Ԇ%^g21��Q� 	���k�a|ǤV.W˥���z�'?��}�=��O~��+�<��5jj����JE|���t�;2�%��\��-����O�X���+.Ûݻ�b�474W��(��zN����V,�<O��%5T�9���d��!�X:��d�c�w��Ȯ8{/^<��U+N[��J����~h��%K�`�?��g�m�V>OUX� #�1#��T��σ�sPT�������������[�xl!hO��TF?�6��QV��W�����j�@���'�֭���q�;v���-|'���6hn�S �v��9�?�0�2)$3��v���-Rib�錒�ͤ3�7�ZPy�[r�[pb�L3֯��V_���r措Bf��E����e�:���`��VD�%�<X(%)*���¦уiTZ�&���q����p)P�W�b��)�!幭�9�$���7t�U�f�'�a�}fQO	�2Ƥ�Ĉ:�H҈�P $�Wxf�X�%XxW��1Bd�0��v]Ѳ!�͖RM�1��O P��%�?f�d�,��ЉLFP�PJq�1(<���4l!B�j��ezj��c��t�5ʌ!\Jp�J+NSq����T#0�Ǥ��d�d��VJF-����z)��rG`�R	z�ԁp�6��ܭɅ��)��g��p60!�"~��<���2����l��}�7n����Q�N�N�Bmj�$̰Ø�Ba]Z�f���Izܣ86�ٿ����Zx�g�{���dG{�34�^5ex��$?���D�}v��{��{ｻv킴�(��3<*Á.��K��&3b	��iկ~��~�Gv����I��@�� ��ad���EuAm%f=i+L�_�=���g��fC�[�.^���m� %[�\��0W����Md=l��yhM�K�
Rv����Ѭ5@B�p��}��jlH�k_y���팧F6.��"<��#��O�F9~Xމ�΀)�������7n���}�\�̝;o���@�$��0>�X@z�ݵO67��*桫�˧���۴����E;\}�՟�ԧ�s��\q����~��K.��X�pO������	UϓO>Y[Gٴ��u�$-�'�"zާH+�gq���TY�Q�++��ӟ�Q��Y&I_���I� ��ݘ�'x���|��x��v�Ŋ��׿ݾ}���������w�y�0�@�X��{D�Z�)�*H��좋/8묳�<���O>�f]��� x'8\P�RE"x��H���gA��{'̊�'b�*�"uD�`6+�o���Z[[��2M)��M����qE#n��&�R��G�F��W�+4����S�v�hc�Rщ㎶ 5�4ˇ�@4��7Ub�d�QgX"�Ao�M�����Kp@BM��sbSk�J&٬��!5��Q�hc2.��)v��p�oAY�r��{`�w��OB��hZ�t���f� ��I9Y��m9|m��0���L��"^X+K�KbrYLS:�{a��i~����'�D/Q�u�����*p��i&n
N1ԞUY����&
S�JnE/��|;�0=��\�jZ��ۚ��T+WtЙ1ф��eHf`��Ԁ���|�I���6�] ���8������k=��Q�M0��|ܦ��T*Q,����R��>����F��|2Z�-r<6V+auvv�h��߼y�����MO?�5k�����^kIK�	�Pث`[�  ��=!�(#!!�a���4_ӫnÆL�
!�}�=����ܥ�\�`���>�}��͛gu�3R�rM��c�W��H��'�7bb8�����׽x�Y(��ri�w�w�#�-Mo��M׿�w��3��k��|C)K/ٱb�Oۛ.{�����ɠ�k��@�U�\��ͥE���o`�@�d���� 憛[�m#��V��hw뭷^��L]bD�l�ʩ��<88T���Q��LO�A������굪��< ��ܾ�\lnڴidx���9_.oٲ�5|)/0X,k���Б���7��]������Ո�"�7�ʙdr��%�磣c�}��L7��ȤsL/����t�5�0n�,�p �m[�Y�pQSsÞ={��Z�馔T��OZ��𽍏?�.�ʗ_z�'7���&�����[6mƳfϦOF����q1G���r��@!�W�s�>���o^�h�����,�?�/r *�����Q��|�b��(vĂ�nu�)yw�(f�L:�^�+�š������N��
���v�٠�o~�x��?���w�y�Y����Uq��`���q�Q���s������z��U�	��ş� _��ˊ]����OBi�`&��U����H8`u����U�(��)����l����p��aM��̛�9�|ۧIy�����XB	?9ӭU�l�R�)���g�`eINg"����f�4��#i���hFέDp�֤�[���^�ʥ�J|Rw�v\ٮU���Ng�J���QIvm�ш:h��T���@䆉yN9���Ch�5�7��<=:��	���<	̥m�1ҩX*�2�4�H�!�QhόY�w)
OM<
!�U�,)��3u��mʥ��7b�u۰��"ͽc���zA�2pN�2�A9H�V*�g�w�Q�u_�}�V�z���1�W�\1�k׮�ႥpF�R�����/ɫ�\F�l�#��(��f��Y	�������T�`p<�*Kl��ڞ}�ٯ~����j��>����_7BM�R�� b��eOV�R��^r�&�0,*�`���e�x�(���]>�9�h���y�Ν@ 
ʨ+�tH8@'+����kn��[F�d��<�#p�
w��dD�c~��/x=S@���>=�SV��ap�76'��t�(ǌT|�#���)�AGzh۳:%3���/�%G����q[�j��R1\(�3��r
x��ŋ���-�Hk/L�}��H�*ۥ)l��H���];v�y�����U�Vu͜}���1"@���Q��P���V�)&id����{U�ꆇ╪�Y鎁`��͛�	n��]�vU� ��a��?V�@ce���0 ��uwz������q��զ�V B�:H ��ojjP��@�*����y���F� y�-�)?2�_=��#�>�(���7ߌ��=�P�?��nP��ЀMq���>mѶͼ���M'�`S-�9`��Y�TYz��$����Y�?�Ќ�מ�>�p�̙m�p���3gt���V��[�ba�}��TX��C{{�����b��a]J&�Y�K����K�� �*zBN�}/8^�����qb}�Z
i*�3C�eÐ�]���0��?��8L�$gwC/pn��9����9H����M%jV�Ĭ��Ϊ����i�����U��K7�S�
b��'�U�2p�ɑl�Ɯ���".K���!���S�)�Y�cv$�A��Q�b��tu��d����H�$,�N�$T�)f[mnn��*�D���_�2NxL2��Z~͖�U���19��'���0}�-r��y�r^O5�e�`��d0�M`���*�Z1m3R�y���]����ԏ:�M(�K�P��x��"�FG���Աk�sdc��ck=�ؓ��G�ͣ�:%U	8�nnF���$�t�"Z�@`����%��\sͶm����k(��,Yr��am@6B+�f3���{ч
}@���P��A�Ӥ��JE�cK�R_�a�g\�QO��hQ�²~���>���k߼��WG���'�����}򓟔���\S����-[�t��}������&�8�b��(��0M�?a�'��8d+i$)�b����]�w\}��d���7(ևG���g��=��Y���ޒ��s=��^ãc���I$O��L"���%��s+NG��-��B._�
�ݸi��g����:T�u��q�d��d�T[Mx=, �mo�U���jB�c�+�`������m�N;�S��Z��C݇�{�pg�rR��9T��J�:X2$�eٯ�M/�s�N	w[�p����;;���_�|類�}{���"0�*&"�^~llT�2gA/�/�rp�t"�6���k���+?��Zgv	 U6��1ɴ�ַ_�Q
H,��3ׂ��\r+EP�E�Z�i;!�,��v%�#�x�ƌ &A��8�� !�N<����̤
F�UJ�t*w�N�X�~�_���2F��݋>܍�x��^�y�T���y�ɫ�֭[w�]w�̘-��ܛ`���<mn���&Yr"�I%��� ��a)l��`�ee4�b�mhh�Uf��V�k He�0�:l���s'n{*2-��ǹV2� !K�@��Cz��c�����AZ�0W� �F�Xk�%�[%��\3%$��G3��H׀ͅ�/�+$��%�����s
"��K)}U������0V�.꾲$���66*Gf�[��@� ��J���؀ynomy���m-�=��B=*��02vR���P��8766����@��z1O1�k�!�̶z�k*�ѓ�ԍ�M��&M�*N��ͦ�5�XRYS�44J����P$R���(�ԖT���P<��E��"p��g����=�����u�|CE��@'���6:�O������5�©�ҿE)���Ctɜ�<+�����^'f3}^OOߧ>��G�LV49����d-�C޿�ugCŶ�F�cǎݻw�����@g�y�$�]c#���)F͘�n�|R�~Ų��O([;�S/��U ��H���xF@���z�'$���g�E�A%2��=3&A�z�����$��;��7�i�ҥP)�G�M')i��mc����?[m�"q^�A���
�?1��8$�$/r�*.����Ӣ����[�l��9G�CC�F��0:��i���ca�>B=������B<��W^y%8�ƍ1�;���?�y�Z�%D�`��=4�Є���t{�zUgsrUeC��*!(%G^��4ܔ�ϝ�0�O�ǔ���-��>=}�0ù�����\fhj"��E{zrh<��l{�Ǟxz3�\(J$7����'��.,QX�H�ҙ�J���cZ�\p��v'��`��S�k����?����z+@��D���y�a05\��X�\ww�0ā�3&���#�tjo�y�UV��]��Y�Td2Ky�Ve�l�.۰a�X�2�g�y�X*�~�?���g?���}�c�m؀��@×^v�Z}TIό�m
Be!���\Ď�F)iA�`�MKR���fl�x� kY��>i���nXgRYb��*�h�;�"9����4�jˊh��FG���-R�ɵz�so�s�.vŌ���黠�XK͸c�4*f� /JY�&����?Q���VA�V�U��
������n�f%é�K$��D�,�c�B� �p2��~��V���9��С>�6�9�>��s��- �H$P#�W�5y6��#*����B�8�Sw�@�]x��@���O�3j*�È/Z���Ԍ�q�m?��m��L2�]A��F�{,�$_�|I9���Ay흼|nnS)�ٖݨ��t��l�R_�)�ּ6���Z��D{2�F`��V�|�P�b9���5S'&��t�|�p�gnܸ����<��ؘS�ϰx*VMDŊ+p��sA=�^��d��ٳf�y�g�}6�x6��?y������o�S���'��5������&o�G�x�E������pl
�L�nl%9J�,�.e��LA�4��Mn0�J +����6>�!���R1L]<�z����￿���>r���p��\qU����yVg����߄�.����J��p����sP�x�(���H!�=��Ҕ�W)˹r�4gv�q���������e�әm۞�@J�c�Y�6��s,}r,ױ<(�`1��U+�����{�/.��M��'�~�{�~[ͳ��w��!'o��=��텕�Ռ�P5�*�u�T��-����~w�=� z�f@��C�jyVg��zu�T+h[��	h�AT=����e�<����T��AU���c���{��߿g����>�<�����b��H�عt��,X}�/�
��#+�-w,����軱��b�qι��o�zρý�-3z{{��t__?o�"��2*��C�[�/\��L�$���ի�Bx�T"e�1U�FR12��2,���(��s%��;֯nV@���}��ކ	ms׾���R�:�� D�sL����������m��qPK<���{��0h�j�L����v:����+U)��� C�Z�R,��	���9�0�>F�Nɪ�kR�S��r��l���բ�"�%ݒ+�r)�|3E�4�\OR�EBN�}ݩ����lWB�W��V抓������J�*���8�הTS�"̗0���ݨ�7t�H:a�uC*
Ip�<Db񕷦o�C3��%�<�̫�X��RŞ�*�P�Y��55A��m�Sr=%{ˏ�u�R�8Rqɹ�t}?�
�j**F1fb�mK�1t��d��քP-�Ri�b��$}쵶�L�l��h���<�S��C9�rp+��$�d䔣z�q���G�4vG��	��щ�@���b���'~��2y*��T���WU�D[[�K����ke	�I$���w�6�a��Ib��PE")qѝ�f)�X$勾'	�E���@������A�Ш�0wM��
��~I��6���>j��M"ɳV�\�y�����x �a]q[+,��[A�5��c�PBI���N>�d:�Y�٫�B�����C���)ij@���JZ�]�xa`�+��7�d)a�*�Ԟ����{qųL���<$־KvX���F�̙3i��[����r���5�Re���׼�5��wߣ�>z�R��Jg�ao�X��Aeg�>{n��pUs?L�������� ��I���s��k�����[|������F��.���!cW����x�b,�� (>��+gz�~dt��S"bh,'���),�u�C_E���XB��=��4z+;��� � �7a{{;�36����(��yS|�Yy��H|����Jt#��u�9����oy�[0Q˖-���?��'��x���Z��*�����XQF�/�p�j�V�1���v���k˕2�=Z`,��mT�k᱑([n��X�\�d�N;�c\���#��F�U�
����U�3]�aθr��Þ��S[��}��U1��������5{��9x��#�<�.`b1��u�7���Xˊ�4P����Tr��V����q$�r���P����ʌUMA��R����)���м���!�8YK,?�%*�8�a�B��9%������5$HR-R<AK�&g��:�Qu}:5�1��w�b��)���H�\��ԗ�96.���KV�1�X��-ST�֖&q��\*S���ʜl<j
Ҝ��|R3�쓬ؤSz�<}<e]DO�`'�����!�Zߪ�����	Ta�ę:�gK���>m6�Q���c��)�s��\rP�̶��c٪�X��װ�Б��.��P�����<�j���4nPu����c�M��� �>�{?|���L��n0���c/��_�0rp,�޽e��_3#m��R}�_����
r��=�|āoA�K�.=���W�^��u��WH߿��{!������}��������ϙ3�����ͱԕ�����P<+L�Ƀ|�ؔkhWA��W*��*Gh
�8�$�=$�x�n�IB�d���T�G��I���Wt�P�O�����{���n���N;c��׿r�%� ���߶^��W����O>�$�+'��ll?�~3�.��S�J�ul?;�La����P�î�\��z�3��
�Ǘ ���Dʃ�pǒ���Py���E���x�RʥD��$����+1����|��~LpFGǜ75
~��_n�&+��3���́���@Z+�c1���b�L��\���P����k%` )�dY����=�3g�s�����\&c�j�	u���r��+U�X*�s�'�k�t��.O/����G~}���i�� ��cP��G�@!�\�d��]�醌:�OA��HlK1��-_�����S���G���U�U����}�׾�5��Ɠݽ��M9�T���t
304�;���7��S:w��������̊G*4��k,.��
����/�̏����w���Ξ�%'t� 1ctt���k��������N��/��[rM��{�����iaǉk��a\$�XXR��dW���q7���ml΃�A���٠��B�.8��F���%߭��g`�ㅃ�Z�G>���ǬV���Ǿ0$���Р�
yг�쑦D��$VWȠ���埢�`�	�B��dm�q�%y�IVU-JY�s��ub�/�����o҃�WոDt}��~��@�6m��@�/�%0�Iġ��c)"�3���X�mK~����~����jHf?vUL�m���W����Uvhõ�g���1_��
^m������)��^�D��[5���,���H�0�ޜK'̢Y���U���<6��C�:$%!�dattd�w���֝��P�Ý�V6Љ�\)�ڮ|�X��4��x{,@��<�|G������M>���A�'f�a�l�e�dm�M�*�����󇇇�(��X�~
��鏎��O�3�R
��K/����/�3gv������ݻ~��}����A�cr�;v|�;�y�_�-��<�����؅+���2̔T�	��0������X ����ɲ���ik?U���*�rp8
��7�>�,x��]�����ぱ�x�ϚՂ>��sЖ z7m���}�����:�\�������;��r��.�����ͰXu�� ������ѷ]�m�e�	~�I���������yެ�s������~;H�(�bE��x�������*�kw�`wSSs]�nPu��!���0<���#�]�z5�ゅ�3��g�\3��:����dL5�ʑS�U�Cp���
�y�>J��a�К*U��J��@�,s��/|b���C'4�� �s�wKK� 'Z���v�V�úH@��tM]]w���?<� �����&}�U�ЍTZ܎�ؤ��I�Q�c�LF�Dr u=?Qlm�i��P�έ\SWY�TcQ���\KkK+�^m%\&�e˖\Fr>��Ҋ+�[l��͛7_y啄���J��xh�AW���z� E�H�W�G�LqSM��y�(KI�]T����8ɺ����T�&���<>|��C]_��Pnܺ������A=IQLk\q�"�B~��%wT�oEu~NSA,L�M2�@2'֛��d�#6U,���7��
T[�������ۓWM"e�mOR�@��ҠC!{����z�x���V��Ol��X�)f7^c�G#0MZ����Ya�`Ó7�H�+�R�~<�"-N�2:VF���h<�oĮQ�D0��m۶e�����DC���w ]uw⍕õ��N:1m�$�Ed4�/p�w���
k��0�z�k-̀l�#j���<��C�m�*�IR��'��Q�ǆ�:U������9�\Y��!Cyc�ԁ��X�Z�[f̉�,3��/�Xؽ�J1����ӕ�ЮW����y����R��ٲT.9v|�}�sX�w��m�4?������I*椹wǳ��-q;Kf���c��3ۛ�,X�u˳�|&�����B�1�|���Z���|ٴ�iӮU�@�����n����h�0m'!*r�<��&@��Z�W�=A�1;	��pUȰ*�F�mmm������:d!����ع��Sj	6�v�E��m�ܶ9���:8���f'����}j㖦���P_6#��8t���^8��{�9t������zT:t�Ю�{ G�}n����R�����P�b~�c�=��ņF;ښ�ڦ??<6kFs̯:���<(��,0�B:�"��R,��x�' ��˙�[Z�xv�vG��;c5w���K6m�����H���6�X,K�t.cI�~1��(W���}���p"��A2�c��vP�_�������ypR��rY���&���'-�����6�cPv�l�x�.&�X"��ܾ}�����̬����gS����:�s6�	p���X�!W7�$D}ܩ�C����
�N��d|�x��� #nX;����/?r����߽���}�p�P�V2�MY�0��%+V<����'����sa8�Nmۺ��K�����};�;��S[�3�=�4`Ļ��^�����G?�ы�p�Z.�<K� $߉�7f\3f�F[�cl,�xB\DOC&Ƣ����V�i�Jl_��l�j_7v��Y�Ճ�w���k*���dY���⩆�{z�L{=�ㄆk��DL���8����R����'��ٻ}���#�mM�矄�4�A�K�c�_vɏ��R�����5�`hHj�;1�挸a�����p�U0n�!��T̬��[-�_2VM4'�%gt�M�ܸ]ojj@��نb3+�F*�u=AE�WB'�*�pl���Ew�U��`XNQ���'r<B�W܉��f�f��t�]ժ�kõ����5�`���'���P�3���'ih�iq�%��� �b�T]��5����yN_�5�3��RC��礒�p�E�5$W�W�ͭ��j���^�nL�eSmC�%�b���tے�'��y��|��E��2�����3m�5e���������� �$�BL�y����Rn�UuG-��񹖃.��ң����w�\u�?~��wv����l�w� ����4�>QD��<*�#V�X0�A���@�릷�n���fvz�s��}>g��$��|����}嵙���r�y��>���R�*NN��ƌd��k�fՌE��:�D�[���p<eu{}��l^��2�lV���pE���2���,9K��u�4/:g�ţ�'��c��B�}e���E��Q�����M�4y��q�G�U�W	�ETyHN�'�*�'��d�h�S�Nk=|�~S��|����������ʗ��A
�wwI������r�Ν�7�#��klә�uq����n���?�������~��S�w�1{����__�� ��=���ĭ.��­[������馛`-���SEPz��������4X���20��ǜb6�p2%K�Qc�Bl<|>�n3$�U��g4�	���0�0�;c�+Vlذ�Cx0�kj*c��=��
�+��b�ҥ���/������ۖ-[6cƌ���7T����Q2�0�a��ф�}ԛ��AN�0�"��, <�D")l�BS>&$0�XS<9D�%�f�.)C
3i&N�/�R7/"�����]w�x�OsXڬ�w{=�K���͛7f�ȧM4����-�Cu��<�y�f�Pf���������tuuq���X�J� E��f����(� �I�B�2~X3�F�����ݢ�2���)R3'�1>�}�nݺ7uv�8E�.E ��H@��s7�E��G ��Fc/}���`��晪�PCC>�����<{[�a�ݻ��,Gt��&P�^����q�y�,��V��x��Y�����L��ܪ�C�f)
�G)i��s��xD���P�B�2��q,��Y���X_��g�}�ԩSxO}�h���0���M����`�Pܝ�d�$*Q�^sD�c����f;'p�Up�2�'�d�E�n�p�l�Oh��=���|^N���t&azM�/"�]f�bYW�c0��t~'o��� _8�dm�-E�%�������B���r�t����Y��9�Ns���.������Lb��Dg&�����f��3 �P_��Q������E�.o~�4d��Q�'Deed �?3>�I9��Ñ9x�Մ��Co/%�hF}�6���$� �xWSUԙ�	'���,��������]jsy��g֯_��G�+b��+-	RI�\V�M���M?3�$Š�erG��g� �O3�K��O}�Fj")�n�������?y��5k���cƌIC�f3�M���qc>���@e��i��lkODcs�/\�`��]-��>7i>��"ԩD�*3$I��./)Z�f�ȭLߡm�,��Ow�4Y*�؁WV�^ǹT��)Li&�n+��/�����;I�߷x��ѣ��w_82T[_/�9ܫ$ܹm�O<��u������сY�Q��
��xJ�СC�[8Ӏ�U�jƬ\��6��$��y���d&j.o0(�ĊU�Yu�9�ˎ�-iլO�:89�����/�~�wh��H�9�Dt:�@�_t�E_��W'65d��D��|�ı��Jo=���?}�[����?��ߗ��G����i=zw�8q���ɜJ��gsX�X�Я���lM-<08RL�ĀQ��&g3��/�rN����`i�n|��ǉ$X%�L�FO@.��s���^�{��b�Ă1����rSg^��%�JRVhҀ�<���)uS&�����_��ן~�),�S��żw�ͺg��`i��5o�Hu����l��{�)�l�X�0�[2�5Y�X�+E�(���Pȡ�T<l"����b�bp$г+�P
;�u�j�U��DTf"Ռ��2��x@A�	Ő:�J��{ө�Ǐ�vX0��L��#��=��$H؅���ik�����e�p�A1K*O��u�/4�j���J3S��R,?r6G�Ѽ�n\ȟ7��i�����:���	`�e��7n���|�>��CMt ��2��E�E3E%ߟ���	��5fW�E�*O͐�Ğ'c_'өH�2�<^�B.|���'SX7mZ�B@_���c&����$�a�dՈs<%��l"@�R~�,��}6cj�sG1����"j+����BT� �\'��U�m��tҠ�e+1+N2S�ј��n�:}����Z���d��������4�С#>Q���9�����T�/H#�"��s�HH-��'�
	}��DS&�a�"��uZ���D䞸�J�dK���G	d�FΑ��T��ț��,#�2�i��z3�JV,V��R����	����$^���Q�@������ �������Ë**�L�R�wvv2��Ν;�ʈ
�r�&��e^�^�hs{ �9���s9�dqP"��m�d�7R��@�* LȞ=���`0`��>HO���K/���˽/[�ꡟ�{�?��S?��O�;�K�p��+y뭷`�~������O�\�2@�	�w��u�v zSa�=}��H((�Ri���xL�s-/a�@��ق�L�fx��)y��<�Q�xyU5� dJ���������ŧxYas�f��}}�߼�_��(���]�x�]��F'Z�b��Rf�G>v3`b(X����׮]���W������� �w��uU��(�[M�Y��H�X���|���I�j���O��p� �
����!Q�����.L1�b	�aQ,��Fa���Ʉ`�r766��$u�%�O��lM��������O�8�9'Z򼆃Scw�����.\�j�Bʸ[�>�D+O�L7� �9��J���FƜE9C듷@��GZ�B! �PxE@��RӁB7#j��2�ϑ���ꅖ�8>ӛ'a��~���W��g���ԩS1���8�[$�;ٕM�c�Yd3�ω`V�dN�K�Fe
�lkjF5c43T�7������`o��l�%�Vh:�;@�@�S�C(&*�!�YpZ\�06C�?�b}C֝֎|�L}iޓ_0u�dd��i)E�F]x�ʹy1:�)d�kC�5	�X7�Y���<q{f��k��H�;"����Q�c+<vJ���L]:�A����'U�^�F�)K~�BjJD�'-M�`/Q�!�`�� ğ5k�~��&�
�I��_R�n�U�i��N����}����'6o��<i"?��O\��Z�ؽ/���TTT�(;7F� %ۓ��b8HEֆ�!κ��C��!Z����S����rɺ���S_[3{�M�6As�-`��a��rC�˯�䓟������ٳ�����;e���O�z����u��-�('N�äu{\B�X�fDUyE__.�L$R^����̤��FutƆ���Uu�x*<m�E��[-F���Z�i�*�s����%�>�/�m�񩒠_�
�ݦ_����n������������7��߷S`�L�c��~z�����c�~������͞3s��/6Mh<|� f&�f�;����%�q����:�>�eL�:�2��р�9zt����r:/�q�����v���1����,9�m۶s��5k�P)�Uq���������G������ݛn��i+l�p$��W��k׮��@��㋦5����S�^~�����r%U�&�h$<�__]����l��ys�P���]]]�d"C#�6��x�N���&c��S���'s��`�q�g�Q'-�|fŢH��iI�Dc�C�Zs���x�l&�y}A��H,���	5mڴٳg�w�y�&6���y�X*V�����x}}-�dֺ��`-�Py�3k�L|aKK���m����, �6;5��˸��g`i�	5+�6���?��F�A�zV��̘Rҋm֝9��ޔw�.���g7v,����>d�
�vӧO��_v�%�����r�<^�=bɦSe��,��5W?���6�%��ϥ�Y!�m� cM\
�dџɸ� ���F��"�SS52�p�T����I 7�*��fu8�9��;]9�ٲQU7~t
���;dE�M��8�lN3
��El]DQ�k.�a��L6g�d�g�2�P@O�VD��׍�u,������U�?M�, �y��0�������t+pyN�6�;���%�;��M$3j^V�.�#���q2M��@��B��'�BEƱ���W���ģ�X�B�ElxM"���+t��z\�����A�DC�ۄ|+�l67�y�L�Ͽ�M&����b�	CV4���DҐȦ��U�X��j�Y�Rɬ�⬫SUU����82�����2�|��d$u�<\Xk:�8˒9ˉ3MW��+� ��o�<yr�Oe��$=߿���^.g�5G��,�F3�m�|ˈ6�Ef�Y�f[��*qr����4�P}`�;��)�;���qf��a�={���>1����{���⋿{��_xᅙ��]qŇ���!ұ0W�>;/d�ӕ�v�֧���r��PiH�T�)���U��]eD�iEp����n��1Y7jdE)���A�Ñx�(�)/�rq��!����\�ׯ�����7|�÷�v[6o�����w_~���p����;���
<��o;,��_��pQ}x(&L&������c+����L�$����k�e��(}�6���0���^k[-���|���#�׮��/~��%��;$ڶl���[o�Μ��o�nL�� ��c�ؓ˗�Mg����\�`4�YY�b&'L�����AaK�;���E��>�����Be�j��0{�t�v����zT�^ٴ�0�W�p� �N`�������|��W_v�eӚ'IB�������띝��F�b<C��Ԭ����_�V0�� ����3f��81<0 �{��:)cig
�Z"�^1*� 1s\z���N�ш�L����7Z���`�)�4x�66�h2��PيC}`++�����\qU�jkkΝ�'��/衇p$O�:���8s_�	�8e��G����������'3�J��Q6�nrK�֋�
,���3���"+[6X"���@�4:<C� f����H���3�[��r���R��w�²��K��>��� 6������&���N������D�zZĭD����tX���2�q��ȹ��u"T鐈q΄.(�E�r���ʈ��*ٌ�?��,��&����.��l��^ÙdX���/���}��� 4�0R<J�_6+��R+lV7�����v�yD
6*0={�D��E�������3y�2T5k�
x]�\p���{�������/l�Bݶ���:���-��a�\nxx�#�'���K2d�\l�a��/v�d7�]�t¢.]�TU���/�p���.ǎ��o|��[o���F`K�R	���x�g̘���~�ҋ/�:5�������E'�b��Zxp(TR�Ñ�h"Y]Q��/}	[��Kd��w�.U{I*іN��1xo�A���q�0ՋP��c9�Y�"�Mbg gQḆ�OΜ5��s�q9�n�r]�ӹp��7�y�ml�L*���qRC_WWy�X�t<v�W�<����e�B�@ScD-�����ȑ#��_��2g�����ģѺ���x�&bfNG*���c �<4�?80�Py!L&�.�Av��{F����CH*���O��a=ɸp����-\p�_t�-�z�[K�]zQt�{Ŋ�+���UW�30�Nf~��G���|�[��w�]��S�SN�kۀ�8zkQYQ[��>)�Σ��%ı��DK����2XHG���G"#1��lV�n4��q]�x��QZ����*���Sݪ$_Q%�ӥ[�p��8q"l��o�Њ���o���6
i��]�mmm���M�ݶ}�ĉM�����M�E'�5��0~������wڭ��D�L&���r$R���0I&d�=�y����d�6�,�z�y�n�M�In�_��Bmoo��Z
U[� �'�o�,����3aI_qɅu��;O�3gN]}�Ɏ��VU�{��oϫ���'N��N�vm�\UY����ؓ�!�Ê����z�5�X'�6eP�*�_Fw�Rٜ�S�LNG5�1�y��1�KZ
��`0�2�,����>+KS�.kJD��� �'>O��@��H:�f��e4b��*���YJ8��^>)3""�u�.I�S֝Ȍ �N�_��ů0):ⳅ�C�7XMd�������`�⽊;�t�j�����$Z�Y�MB0�A��J�4�j6'�#	�S�Z�����Pʺ��%L�%���D��h��Q�j٩kO./�֠�A`}3�_��?�ɠQ��_�5䕨o��p{BeAnO�1CTB���Q]KA�TWvw&�浄�鱉6��Ñ����-t[��l�ɦ2YlX�.���%�Ҽ^��I-s)�i�$��N7:2�hBJS�����o����d��B��9�#u8��=�����1L�b�o� ����I:�H��u�jcS��Xp,Ɏ;Ȍi��O��x 2������G��52�I�?��O�ˌ3<� ��A%��?ؾ}��~��	&A��ݻ#=z4D������/��5k�3�<s�=_ްq�����zz�XVR����1KIC�JDy��'#��`=���ب7Fy9ce]0�JdP�mUm���������k�}���ԖC�'Sʂ��w�W~�k_���~O����曇�)�;V8p`��ӦM[���S�frp���2��1@�|6���a�q�l��s��V�c)b�*T<�`	58���k�����K�^3�̲��'%Fc�&ҟf,��m֋.��w��j]�������M���{﷠J��ԧ`{u����9�6�t�-^a�%������ܘϞ~��7n�k����i�'�,~4e,�Q���P226�Bk�B3���(���"�SY^#���/Q,�rڪ�+�?����|���uvv��x�����ڎ�������zw=�@�D*���'��ݚ5kF��`հd�~��2� ͼ(�g詈���.%3w�����n�B�)�(�B$X)"�������3Y,�E�Ƶ;MǅŅ�}�-�͟?��.�͔)S�Ιz��Q��E����o�s&[y��-[ �s�N��ȱ�������ٰ(]}�|V�O �$�pބ�Q�3�]q�>/U�zy~���P�@/c�ٙ�߅���%�DM��D$��B�[Q{I��`�Ta?(���Y5Q~1�Dn�^(�e�#�b%��:���0���P_l�'�&��͉ؕL�<̭W�Je2	΅��
Z;)�_H�����&a�E��"tE�M�ByNNW�@���颃3�N7����o�I�/��h>)bRRR��3!a��r�N@@&cy��
�;��d@HUU~���<]�+uA�+%:�X�)+���p�(Y��:��r���i��yŢ�L [� ����v.o�z}>A�K¤��2|��� m=�=X�	&�{�|�y�v�+�6s�@�r��={��C���,��ߢ��>|�UQ�v�5�b�/��2�G��g������y! �Ϟ��@���G?��`Q|po����;k/��S���74�e�J�)ESwoߺd�@�)�H�ڬ��Ñ�KR��� �J�XK����N5b�2�#�#s��d�:mP�Mco���;w���<>(\W P*�x\��1��>�4a�Ha��0��?�mۖn��W����o��M�b}�.\x�e���V��q��Wv��A��K'�յ�8n�t�9��a������]�I$��{�8��؈���G�=����g-K
,P$<��2�9��|"N����|� �q���.���$�*�&9��
0����D����f�����H�X���}�W]��G�	�w�z�^H'p�mu�u�K����{x���э����>�ʞ����[o�n��[o[��q�����]���
8)�H8-���,�|Q?��h4n���{�ÃCU5�
��w8�V�] AJ�f�y��s���Md��W�- ~�ڱ%���x�%͛=���r������ݚʤGU���W�$�}�����~L}˾�R�o�����㨩���PQذe��a�Ĉ�����ܩ�����X:guS6��4\ߤΙ|���U��al���T�0S��� f _��{�>���{Z���CfD4N��^���r; �`������]��*�A����+���5��,^1�u��������믿������c�[����>��O�N����!���~�ر�ƴ�������r� FbQ��莖=�ʪ�Z�l����u�hh�I�Xt�d�/��<�����ѣ�������e�}=7�2����f(�)�ۉ +/�9`�Ќ�V31B6��㓝��<�66J�I�.	�G@�tꭲ Ʀ_fUEl]P�X
��9E��﷊j��H\$2{FD�Ѿ����j��5kS&M�%e(���d*':R�m:K�/�(%�n�F�.�fRDRQ+l-���ɚ�ثN�%P�To�EDe��S���kY�j[[pԼy���mt���w8������p>�L�-��S�����<-�ڸ:3�浜�`Qܢᅇ��X*Ɇ�Q�,�;k��Nu��nmfK�d =2s�O�A����RMϛ$��B!n�G��10�n���R��Ʋ�����N"��ά.'s�\��������7�>��x���b������|�~/���?�Mu,*�(�R��Kn��G�_F
5OL�:u
��аm۶u��AЯ]��СC���S������ϥ�V���fΜ	�4��/|��{a(��@|8������x�K��&E��e�G���X}f���{_�U	Ͽ�������qi�3w�f�kJ�@�e�g�^q�� OY���������d��58h��kj5�k�.<��W������?�q�]wY��;w����饗z|^<~tx���[ny衇�#�3�/FB�q�٠��M��x@3�w��N�jFg�"��)�z<X٦,�ڬx�!�]��a�V�$��/�2�saB`Z�w�y���X__w?�o{{;��o\v�]���-[(d`����1���/$m�R�!���.���+��.Ћ���5��<�(�����/S���9�^v�	`Y���8͍"6��?�i+�J�8s[���k���g?�7_s�57n�_��_1��S�Pa��U��ʕ�=�����s�����⪫���w�ich��m�ox�kE�$�2��>�LoBR�]��b"3nF����bt�1T�ݰ1f͚��g�|�4��Iex#��ٳf���-Z�����c�555ao�S##0�_}�u�����e�ՙ��l޼��l2+j,"8�v�QHau	b��3� ��<����Lz�<G����㉰�0pC�Mg�)l�P�B�����X��t�VS��I��?.�Hr7�l���SK2�&>f�>��o�;!��I`>��r@�X6Uw��5��v�Ώ�
�E��:�s�=�x��d2�5�k
-�c�ϥ���al`�513��l4���V3�렑�GhA,ִi�v�܎;�|�Z�4y�٢��~S2Y!���%�Y�QH�����aD�8��3��ġ8��y�����IWL�J���
eo5�5L<BI!E�!]a�c�=����׿�������B�K%�s\J(9�@s}�m�(��ע�|�2��WK��˖-[�`�$�������ڰ�͓�7�7������ys�J|@�W�Z�v�|��W^y�s@�c�u�W~���F"#==��w�L�8B�a�oݼ��p;�
�rۍ���ˡK�̙�z�j�;��h������_y��y���P�����vY.�Hy���<�U���`��\D`g�J;�!�:�O��a<���&i��� b^uy���lܹc�I�`��}][7o�8iz�ёH��VE�'O��p�|�f(	 ���;����:l����q��Ӛ�9�^ZZҲ��"ʾ�\��A/eT)�W����txd$-b-�����	�Y��7r�N�S)��q	7@FU%��@/CB�4*X�I�&���&�5��I��{JK��jO�� ?���Nn=�]*����P�n��^{�q�y^����#N�cJ�����D*=.���|:ݎL.=͡�7o�6w�1��[��jc�l!��l�|0�9)�M���QP	!�/��u�Ω��x=��෬��Jv����!>ג�����D�b�����HMհ;����Z�%��ߐ��_w�SO=��]�CK�eؔ��������Ο���7�n����%���ኒ`UiI��nu;��T9�lU�����ֶ��
�>2g7s�pH^1�1��23<G4��[:���f�IT�@U�>���%v)��.�h��g
	H��,T���r�W�y����eee���zoϩT2��]�v�e�^�c�6	T.����yuh �d�[�	�O��CH�bw��>q���������X�"���"#������d������l���:&�x���4T��������!v�~������W���\}@/�^��6����S�"?�8��i���8B�"1<M��|=�j
�ɚJ~Z�+/+T�.Yu�>�abe�:���|��\w-���[�aN�h+��B��!�p����MX-�3�5��tXD�I�6Ra��I�6ҥ��Y�ʲ�\�����j�����uw�]��n�65̀�!�YCbxu-.�Y�'�I	��Zq*��eи�Y�dX�!,c�X�7:���5�ۈP���r����N�5�]Ib�-�Ã��L��+#��8�3�ͱ	�@����q:�/.L�#�f���������F뛗~f
��ŕ7�g��С�܊�����ۊi��k��YdF*�b���|�.7C�M�6�;v���%
�f���G'����;�=c�D��	�' =�p���_�K�:*Um:�d�r�9���|�3Ɍ3�i�9Y�~=0
D!�+>ԅ��Y����#��{�	��-ľ"H�9��;�5릊O_��4�fT��͘1c�;�������ʭ�~�x��/��+���ȑ#��Y�xqS�xL��Y�q�z��+W�ty=555�fL�|{�4���9眎�^n&��K�Z�*.��q?{���N_��N�#�ccf�9b��#�ɔ�@��Bn"^���j�r),Li���Ȋ`�{��䊶Änk*0�.qU�j�Ǐ������}/1�`����p����ϣ�w��7��bN��AjD���q+�|�����u���-��ĶL����L&+Q!������O∸©�^C�M�2�N�+1��������?������-���/�ُC��"�&��-s�Vv׮]�7QPNe&'N�p��ƍ�$�TM����vv����E�E�[9;�b��=���s	�8�:{��rI���)d�7PS[�ϟ�d$SZ���` 	�M'K�z�� 	��ﾋ�O�~�����__�t������T^V��܇�y�_���O�9i�p>�#.��tD�/�{�S��F�3O�e��[9V�v�c}b��.��v;�vN��+\�X�-���{���(I�V/pyOo�� ,��c�)�\$�˖3�-�h���8k�l��adDt(P�TL��>|��gB��o$?�D�Ў��N�}UM&��/a�(fi��q�`�g�ڷo����t��N��J��u����0B�cJC�$F:{�	�T<2{�t`����?m�,�%%h���B��+��D�śߐ�)M��b�����0�,6Q�`ޭ@�'4:�;�|%���t �����4��J�@"��H����}s�v��ux�>ܤ�,T��K������ӕ?���'G�~a3����k�c_���H�,�t8�D��uݞqeRih�\&;�?0�~TMu��'؈�j�Ӂ}��]8��O�49�L���۫^��s�=es�8�d(�֣ǰ�q��H��q���ȣǎ"��*���`�.ǿ�_Y���q^}͕/�~�"��p���Sz�U��f2�����{�a�	:���U�dX���d�T�
�A����f�ϝ9O��|:�v:h6m^��}�g?y��ޛ4�����g�����5oM�0�s�펚ѣ�����ؚJ'Ǐ;�o��w�~kM4h$:r�W|�+�B%?�ۧҙN;oz�%T)��1��pd�j
춑xlL�h�hDd�X�!��y�e�Z�&���c�Ƥ�d'0dSa�[VHg�����v�ȡ��K>odx�����p,�wwK��N�g��%�7O�T��w� �O��$���ں6���9k��������Z7f<$xמ��O�./[�T�X<���N���[��߅!�A�"T&�P����Ɋ7SO=��
�55[Q[�E!寸�J���O���}e5���%�ϛ7��TǱc�.�`��7��կܙ�|��y�7��'�^�(�Pl9�L[�N���}�d r�/}��./��(F��W�S�3%�����P�{�qWh6�R�,'��/s���1�$�*��0������y����+y�X嫙<'��V{� �f�ݲ���jj4�����a�������];n��Ƶk�nۺ��*^�#�%p�y�,�w���ժ�s�T�f�9�.ԵX"100T][<�Ɓ�H�c؜�o�(�6#OI�4��B��eJ`q�juC2%�E��ޒ�J�;0<�#z�VQ��p�{L�D���y9O�H�(̊7H�O��aax��Ot�%��h��a�z�R��'&���ڿ�o):��u���;�ރG�>��I'�Ν]Zjm=���X�&H*�Ε�*0�d"�z���������
U�7lڼgOK0�UVՕ�����_}>Oݨ��������e�_��N;�m���clNG�����	ѥ�:�N��%�.g�ՌW��W_6僩`t;/x8�"
8PJ�X��A� E�Cn�a��UvLJ�x��Om^@K`�[E���Y=	�VN��%�w�u��c�`�ٔ�,%��,���h�����1_)/��7����2�^|P�"���ō�3�����f�s�Tokkks���/�%L���75Ţу ��yU�m�ª:u�6`�p�Ho7 �o_������O?M�rT����Ҳ������B�\]�ns��9y�$�����7n�x��:g�ZE����U0���Č���"�v��ǆ!]E9�S�h,�?�z�M7Q��tf��ys�,���w���.�p)��__{�����?;GU9�
���|��1��	M�G��K6m����u��c]Z�M�'�O, $�Mr�a�&7��Kg&$�E
�� ��"�Ib!�Y��K�(��E3�T2�Ux�Ͻ���~��@��}�@SSӛo��$qzs�@*P{94����ݻ r�������Q
��VH��~��O~��nj��koL���De��rQ��PT�8���Q|�,��n�RF��&�q
c�.��B|������K/�̯Z��{��^<��[��j��n����/��
N�0�l;�4��U@����u5u���GR̬�	�i�� U�\��T���Z�u�kq�������9�L5X�9+bp��`�w~X�>�={63�ol�*�?�e�]T�����ٳ ���=g͚���8���箿�z<��B�<L4�/�u׉'�����v8JM#���ʜ`�T8o��LIfj^D��q�mN�7�t��ɦ�I�'
���UU7k&��)�.:.((��P�<�\N��2�烬s�!DF���*Ř1ucGU�oƦ�G^7��iw1��O��p*Yy��kU �	j�m�Pͺ87
o���f��sI�b0fbCΝ;���y�����lll�H��$�N�/��ʀI�q�&N�vt�~�z���q�V��é�S"���Hp�vG�0�Gg4�H������Ҍ=s&֗����E�uax�Z!	��B>�uh���/��Mj6ƿ��23�����b��Y�
\88�I^韸�m��\���3.2�����Y��}�κ��k�09����nTH�!$,�Ͱ]|����,Fp�#��^��J��P����n�<e�$<�X$�J�3g�ٶ�q������d:�?��ݾ}���|��@y���--	�����\�ay��#�}���S�Y~�	�&�����ή?�� Bw���w�y���������ݻ�Ν������'������3)��������L&	@�֎~��DS&Oq9�}ߺuoCJΛ5�y�Q����k�p8̓'Omٵ�a��~�%@XKK˘Q��j�����ϯ\��l;&ᖏ�X"rsShB�d�"�Bq�RF�h�T�<'��y��.��*MA#r�g�2a�;���#_�����f�*���M���O<1�����η;��d�������.�g��%3�.��Y�m����������r��S�ݣ��C�������J+�|���z�����n>�zxƌ���g�Q6n�����b�#`��{��H�dԌI���[���hzᤘ$�< x���paaCL�:�a�P��Q��jk6�����血�#W_�<e�H*�bŊ��mث�����YR1�y�fl03vlE�h��W���[o���@��B$�29Pu4� �;�6 tQ�G=����
���YU�@��N�'̋�1��l�(��2�j��vC�k!�d1za@��qꉖ�^p������ö�Ї�b��Z��mi7�4ܴa=�;��%��˫_����:�k��VO���Y�xqEu�d��t����W��6��n͢� r�dV�R�±�4��Mo�D�HȤ:|� 
�ى�.�fJJ�c��px����3��j^�YƏd#q�t7)5-���Z_6�q8,`�B�h��Ɋ��a��s����Ԕ�Y��
��dj}�c�$
mc���6��iR#F2y��r����lAE?�?�ؔycu�y�_�V��z2��3{>��RYY�{����AF%��I���x��X2:N��K.X���j�Ν�t�t�3��P �;k�8��2\p4Cww�)��&�a] ��G��z�Ƈ��@�DHsB��N)M8��h�f�LL�L�#	dAI6T=a��}�=ĽC�C��+���"-'*��lx	d��2X��N��Y�ђ	�U�5�,����o����&�t�|ZN���n�b;�x�L�B�.z����ş2鿑F����,mV/f�
�r"�ʾ�^(�{����� ���PT�M��WO��;C����Ż�����4�M��b~ҤI_��5��5k�瞓;>��#�w�q���9����^5j	����ft'6�D
�`h�\+��a�"����ӡ�Q�3L�mP� �l��z��G������K?�d	p�Hx��_t;=��~;N&��߿���;��އ��
ӂ����{����eɒ%˟|k�r�+�G�->g!��,
d;����-�煐8�"�)F��\X�f�B��z�%��J��@���sG7&g(�W��V��+V��7��E�X�MƩ{���HŊ�������k�mٺ��/�L=	�+��rA��d K�קN�
�o��V��|���4�=�{(��:db��b	��Z������l�H�M�kJQn
'���Wb$�P�uL��b@����駟>p��	z�Z`���M���ZXd�dm�� �`�aY��ڰo/�袭[���U�r2v>%U�sr�ь�An������_=z�����#��b�4q��.�zE܄4�؛�f�.�;S0��^�'��I�����𙌈��d�m9�y�H0�؊�>��e�^��/|���V����.,PŨQ4��8���F gߡVJ@>�fv9�Kt�y��^*�$����2g���R��������p��gU�fL�(+1�>5'�e�YUЋ� �D�*���`�K�;���G*��^�
��X���M$�fq��%�^r�ϛ7v3F	M����4��S�9��@	^�D�����Ź ����� ��E�4�pv�"v�܎ŝ=��*'5�� ��0axh ���sa�����a�`�/��� /4׎3���R���q����b���P�4-��Fax�N%�fS��
�$�mMvEM�b}DT%��JiP1�z���/��5
u�9j�I�d6�Ym$��*�Ã��^�(˪hg��,�7-<��� ��fuʲ�vY���������@ �O��~�#0_:MJ�4 �G+�tٽ>7��g�2%G�j�����G6^*��zI �|*��;"�6�g�8��]�7C@ �.:gAO_/�P�����K�i�͓>|Ӎ�DbÆ�v�����k�-N+�qEe��e{�g?��in�>q�ľ�~`��-��]�V%Bp��Hg���rΒ���S�z�:�]�d���aS%��,NF^p�Q��Q	�Y�Wl� }L���->����~8�(�d���� ��~L͵�^e!��ܷ���yӚǕǅ��ǎ�Y��M���`�=��]�,���,�vvzB�=�-���G����3�����ۨ��ؑ�}��{���֖�SN�̾�4�z�s�K|e.���ҡ@�'��K}>�k���X�{��</&ۇ;	�<��E�A)�p������8�6��[��"�>8~���`��w~�K$-#~I����/���uZ�«.�mi�˨Q����h��?^m	8��]�7�ڴ��7�=�"�6�J�w�+���T$�U��#�=�sw��Oh��4��l}1M��?�s�cB�9J�AM�bY&Njؾ}{�`?��ꤌ��P)	t*<������!E(a*@�C%K�U�ūg�ل�4�'J*�+r9}ǎ�@yiY͜�;w��'G56yC��_x��2�Hve�j�?��~�`�f�Ɏ֌�U5��D��[�-O��1�f�9c^�������d�Db��#�W�^o�˸ Tԅ/���h�[V76�u?�a�e�{Oesi�"�2j6�K����%�g���I�ŖH���򔋮e�67+T���9��_2�0�A��#٤]d2��"'=�~�G�[[���]c������ջv�쪫gΜ��ǳR$�{�w�ͯ���;�F�^���O���q��'I�
"�u�ͳfXd˽_��%����"�Yo� fL�Q�U&	�l��R�=��쮨I�L?�5e��횚�(��ld����a�}}*E��q4=O�@)����"�1OÑt"�;��5���n���݀� ԄƢZ%)��QF�D�2�+Oj95��gs���ϋ�A���F^-�]���G2��f�$��b��F ٬�T!�]�4������=vlC�h��R�=�PG������h���{8"rq�|���A��iLաC����K.��dt9p,�K.�����|~��#{}�X,��ק˩K��Ѱ�_���J'�<��"'+F�aT��9�[;��A|x�iu�s8+D?�7I�lIL�U�]V;Y<�{��;ɪъ(r�A�h�&aQ�@��'�cV�J��)e'1��0"��©�$�%��|��q�R:�(���-�;v��&X^Q�M%�{IM����Ag��o�=���-a���qK��["+�D�,֊�ꫮ�𛯽��h�TN�-��7Ϳ��?��#+u�[����<��|���/����p+fL�p����P�8��m:Y4�f7��?�o���Տ�;;��/�g`�����H�zp` m�����'`��O�6m���([���/\�b����믿��DY-���F��2rj�л�:&ߑ�ZS�@���ǡ᠖�Cx}�޽C��qIl5�"Փ�-�D�[^V�_��7`~8"
� �8����"ǭ���J��=���V��5kִ�Ʒ�zk��uW_}um��v�i�^ٷ��ӟ���0/�1x�]n}��O�{��#�`&NK8FW�3/5_�@��DRC$Qb0�<�H��T1}t��ҒT��ƎI�!�HF��@�s��C%~'jT]��`9D�����{챬J��[o�j`����B::NTTT �c��'N<��c�ԢE����� ���qqmٌ��|��o���/��y�-_�������d5���Q��lvї�K)*X=嘾>��>�'Ҏ��ڙ\ϕ?F����T�Ib�8S���nU^Q&8����͛�\Ē�ihX�z��o��9?̟?ߦ��{�=KF���������o,zZ���t�r:QG���("���8T,.|�f6�d\镜�)r\��RMS��=�H����t���Z�|,۵i{KK���۟}v���]6nܸm۷?�䓽�ð���/ ��^}Vm�s�FP?X�}{[ y��Xe�2,QL�!|)������`K�D'N �j$����B�8�6��/e�E�G탄&�����#�3���T��O���t���~P��ܪ���s-�ʦ]󑼛��:݉V���bh*m,�DF�`Y���'ʘE��"�~.�@��blV�Z�����o�R����	�3luؙ�k�H�Q���f�
�ה)� ��/;� ٨�#wR�o�c��2r����V`�sD�Ӌ��L�9��3R��BE��H"��%�UT�7<���E����)9�j�mr�4��,*�)x�H������.����q����	IV,E�_���O\�rZ�/^�TVQ/�%��))W��X̪��� �y��GFF؅�Z�=�ز�!(��eE��̮�l|�j7�����r�\��()M��X0���;r{� |���@[���]|���M$7l�G���{��@�P��I�c5��O����b����/�{���Ϟ5��˯||�S��l��<�whS4�B�:���D��p�V<��;Zx���ə���B�'|����;�˩�X��s�-C�4�i��h�T�ｻV$~mUmI���~Tݸɾ~xpp���]���i5ucG��7g��--�R%� d��͛�+k �Z��y|�C�־{��_��<��(��\���S��E�NQ)����=t��ap(�<m���oP�%6#���"	EB�5~/�uummm.������뮅4������-[ƍ}�h�-\v�ek֬ʇ��)�8��`J&�ӛ�L��+J�r�������khjصkwWw︆��{��gnב�(f8�N���L����'��G���f���9��|(&x��d��S_��zaڨk�L	\�k�^�&`� ��0v��ٲk���=x�ȵ�Hxdx۶m�L�K��Y0Yּ��M����o���N�:��{��e��cƜ<|��Tǁ]{`�^u͕�ӧ���Mr(	��9���)Fe�	����	����6�����;��~��1�/jق� 쒣*��K�{��EW$X� ΰe�h�~�zDEUQVn�����{�y���S��2}ƄCG��w��%␰.���s����X����`���={N]Uņ��LYi(Y8�pxd��}#CéX��0S(X��ՙLe>E9����x��~ʪ�6��.�N�N���~�R�H��s�_�{d�2:�����1C��q7����\�֗N��)y�c,t��: ����Y6�y,������Zd�3���b�$}�q�r%Q���"ky���B�%49N5i��
�Ce��%� �=f�H���/:�3�唍�ˠ�eI�g�.{�������0�Jf�I�;y�D']���0DM}}}ee9�pxh$)a�b[�t�����V�N*ju)NQCHi�z�й��u�"Ӽf�� Ǟ��4ѿ���Df�E�Pb
��R܂�@�g%�8���� ��r_(T�+ >(<�*�'!F�^��Q�U�dH�&�	J�Q$�>+>�P�����L*�:K�D�;i�{k}ft糠j���B��DKf��]�O�|ڋ ��pA3z.q0�&�?+ l�|�	�!���6)[�X��˗C�_��8Hǎú-\��L�:��SS�N�����xz��G�#����m˗?	�x�u9����j~��Ǐk ���kl"��W��ճ+��S�g&�E��X'!�uss0B���r�9-��J9pX&:�A�
ǉ�b�ԩS��5I�96ń�050�ptDd��쉦R����㕊� �BSSSkk+W<x��޽s'�<�B|#�ݼ��q����㋢�̑���,��n����z0���N/�H�DhS3��h�l��R�?������K��
R�9����ӻ$�1��
��о2�W_y]����}{`Lh�[+;9;�bYfS��
�-�L�K p �`'M�D���۱cf	O������z�'~���$H>2K`��X��?2��'N�����bx���x�3����1.���<�����,��t<��?�jժ�>��[7u�ԃ��a�N�<�TU�A�����|��e����G�z��֟���0��h�G������̺ꪫ�čb����I�> �I��x0\~V\i�Y8����lVf>�DF�;���岻�jA��F�ؔe��'?�E	���ٳg0����D�a�l�<w�L<��K��)֭}'��u�����L����s�[R����dD�<X�&kO�2�
1[k��)���N�E���� 	Ʀ֔v`��bU4(~���\J�w95!iq�W�q��<f~��Y�Z�+O�4�ߋc^Z��h:M)��1��	@�$�-=�$������k�����ѣG1c���'����!� ��N~�\;	�N���N 1r�Z��r�o�R|N��ӹ41�{�.���7PQ�5������0s��v�7��l��K�4*EW�;�q4�U��iv� ]����<�2bU��#����o���)"5Y=8�/�{q�A�����x��j}�8}x�Ǻ�h��q������-��űI�?HF���`FeI!�n�ep�r��ȕ�M4y��dl��pD�a��9��X��v���{�[��Hdc^s���q몕+w��z�'>���9{.}/QR��(vׇ.��������n����5s���amդ�p���سe�7��vC�c=A��O��)�P�-�V7�$5�ɫ���s{�ld�z���x�.�-�~v�-�|u9 ���B�5L1��6�Ȑ��5�'5]�*-k5���qh��(�ꂪv�3�܁�������~���Ý�T�5��{�����ٳ�C����U+%'::>���%Fb����գ��ӟ��i�F��䔪�����#���D�V�;��Լdw�+k��IL/���	�K`�Q5�ǰ(���e'gey�wܶt�R�1�mm0�ȸ����b��`��֎
�8� �=|�bU�*+ .�#3�i�R,
����x[��2<�աDb�O~�7�~{&��;y��z��T�f���@STj�%��òU(����>��4ab}����K%�CP���H%����AWٺ�'qz=.�"����D%���|������7,��=x`o"���)I�Dg�������eW]%���}�{��N���>���_v�;o�Ј�g�Z�fMwfo۶-З������m�8��ᓟ���o��_�&�J�"Fj,���g�K��co�Fv�n�D�����JȢ�Mx)4�U6�}�e� ���L�c��K|%�e�'y
;ێu��64�O$S=�ݰ�O{�׎>���~R�ر����_y�l"�կ~u��K;OuOlj��]�vo}o�~���i=nѢEN�'���=ފPYO������6����f�@S}&�7Q��w��qFS�8�����bp����}~�0�����З��D��z}���hEjI`\
��:�*�Sּ
�ᗔ�-��u���rÙ��T���d�J�S�dω����1���hrF���K�h���*����W2��6�CIaC@�B�d��d.Cn���d����ݞ��j̆?X�B��(�n�
:�*�wͯ����N|}Ym��bs�,0K:���|��bIq7Tl�d*�r;���d��*x�磳��j�@�^���\J�n(��~������cJ��I��0Fuj���B� A�6�/���"b$��hQ,��`c@hP]z2㰻z{�!^l6�����8�]c8r �Ǟe�=�*��]"A���3�<�V<6;�����n���0�'g��+�ђ\.j�Y8�FG/YP����̙ż1ؗ�xq�����j��]��v ��͙3����?n7��r�\(����O�s�=��^�n�]oW7!r���˖�}��+�{n˖-�k+	zR���2 ����$�"��+���-����O�pF1U�A
�J���4��I`gΒ	:u�*q���;x ��rS���vY��ۗ-[V;�>��x�	��?��mnn&���.�_y�ƍu���}�X+�e� ��ǀ7m���x(&谉�$���f�4"�gI7n,>����ű4��>80e��jZ����x�,�n7�i � z^y�ݻwC�[��·��8��1a\p�������Krkkk]NwgggR@pf|����kG�R�9_�x�{�9����o����׏7c{�[H�2�Pw �����^�?Y�o;��ە%�����$������	!U�	S�1P؍���K/�ϣ��L�xtxʔ)x����_=�4��ꫯ~��.^L�uk�~{�ҥ�f͂.��b�]w�u�L#��[Q1�����?<y��%K�|�[p=dq@WU�غX>���Ǘ0�V��4 ��4�"������$��3
����u���D��U��444�T�uw2�&\�b�Ŵs1ŪU���_=fd���/Ɛ�x�ܪ��;�f�����,��L:�W�;�` �֍b�;���B!�L��#�#s�����Ï�Jּ�X�"���x�]��4�\�׊���8sB2�~��_/�O��'�Uk�T��0!؊�[�u�����	Eޔ|��7��`��r%ax񢰣Qr{�y�2���0�~j���i&x�ÌJ�,2���͉Ʋ4��`9�ﰓ�.a2;ޮ�)[(�$"�t�U��6��Z��n��̴������}~
!��_��vq��^D@rZΟ��e�Q7�`���?�'(~����:�}4��� �j��kQ�)&�C�^D�hZ�����=���!c3��ʼ8�B��ů��޿��崾�}z��O�:���\شr����6���F�"�� 	�t��.)��VD�_��Y�zn�O��"('�Yu��}(2RQQ����$�"�݇>��f�w�ر��s��6��o`��<t㭷�ܽw�de�7�Sծ�:瞙��sdf��A@81�=~���(0$AQ2"I	8LL��3�s�w��[��4A�w�{��~�駧��j�7�w��[/��ʉ�Vp���C^_`���0��b��%K���k~v��ֿ�nY(D����oh��/C�|�L6ʨ��y9�M���0Dȕ�5N�<�5�@�t紈q`�1a�R��_.b�ʸ��eK!���%���4֞��CG��ߵ���S'�}ֹ����e:OP�K�Q�Ȗ�����inn��}��W^~��rC�զm߹�,9��3��^0ٶ�΅��|���������n^C��M��Sd?�U<7m���˗K������n
�+�HF�c�L0�*4AN�B�&���NOhH�����__��?;�30G�Ommm`�lf̚	0�tt��SmJ�$SxժU����t�����H{[��y�ĳK�:e��c'3�|:gxt��~q����,���}U��-B��(	{c�	4����HCc,��v���L��~]�UsS4GC������q'���,)��։(�bwz��,Kyh�W\u%&�ګ����w'<���
���K/Y�dnGG[2��'�,Y<c��oX��A+���5�-P����?0m��g��B$A�qU��
U��Pe�J��.V �����ZKm �,�2�IW��9�wp�|�mvMMf3�
6�X>�J�D_��_�e�M���#��1�w������_,+���y+��  ��IDAT�I���9�t�C�����U]Q!jeu9���5i�������:G�f͘M]�N���ڦ	Pz���e��x<944�I�1H��"�$.���I�{μ٢s��GC��4KF_�7l�d46�ũ�����KU���0ٻ	]�O������^u˴d��\���f�>h3u�g٣�3G�wS~�CJ����*��n��URT�p:O�w2]��w�a������w�^RG|6���#-GO��T����WJ�e��_t�n�]/���=�I�����.|S���!��&�lZU�|����%������X2�4�9��	]ex8��hT1��#%�;܏���Ysˉ��x^^��l�SC�7J���5�0�)ϫm�O�:_:-$CH�,f-ˤ^C�ф�ŕ�"Ɗ;��q��cdd�"&����8��ۚf;~�EU�H8A%��S�g�C���6�8��@U?��>sR_�\�ꢑ6�;0�<�B����Ŋ�����NT&�g(+Y�����?��Rqe�Q�x�:X��d�m��o~�GN�@�c�U�Pc��0�ҝ}�y?�����ާ�zj��S(=5�뮻V�yڪsV]��7�pü9s�-[6u�����0o�F۷�����a?����sO�`�P]��:�����i�K����u{\�wO�h�8N�fqN)B*YK����(�l�\��H���n�9g��>�h{!�]w�u����k׮]�l��ի16H����A�����nM��[N�~��>� ���'9r_������~�w�����ׯ_�]�*���K9㣗dR�L�.����c����8q�U���K�EY��"Ϫ�Y��v�
ñ���d�9�����
�3�;����A���۰��/��J��������S&ac'��O�����@�F�b2��&Q__�OΜ?���_��J'L�i�SxD� ������\�t1h]#â�x4*|�)+ׁi�å�>�I��8v��$mS�YR_�թd�_R��+��ٍ�566�ڵ������kq�Y�f���`�{:�_xĖ-[~��_.\����jǎ�x[|�d�i��F� "�(L�ė-�ƌ�A��x���h�Vc��I�(��r�86F�Ň3Y
�r�@Q��E��*�+2����Ȧ0lov�M�>&T$<|�Yg��o��:[��H*U���k�����8��sa�����P.�x�6����1�T:��	������]_?w�I5�������3���D�J	5�ˌ��B��2��Fy��-�Z 3pQ��A�p�ur�R���M�.!NU�:wڥT�|�&540��'�Kyx�J�YB�c��w���޽{UC�}ҙ�x�VWW7{�T���	Ǆ<
�&"�2fW���a��d�~ ���swLѮ��
�X�����/?�T�w�zHY��,㶙�_�>����/pYl��I�x<;��ύm}��`�E<��d�'�5����rQ��)��(r��nN�0��n���ql'�~��n�M�ҳOrQ���|@B� �	P-Ͽ���~Q�����W��ѻ"4�� }4'V*z�{Z�����;M[q��.>�����d5s���xj�����u��]v�e?��Oq_z�yծÊMd��]�����O}��~���Z�x�~���|��%���^{-5A��)S��<�t���yd��mMMM=�T��v͘5����r�=� hT���N��z]��H6Oy��C��k��I6TW�t�Ϛ4Q.�7c���u�b��������r�'GE�7�9
ԉ^�JަRg[j$*�[���ꍛ�lܴ5
M�1�UÑ�$�Y�b�7���HS��姤VI�kj��7k�_{�-?�	���ںzѫ�����O��k�̾����M[v���RR$	YK�#�Z�i��릖���.Ѻ����`C}]Ow������ឧ�����F�l�|3^��������+	c�D!��sz��.C���8HUUXC��kj��<�����84A��NW.Ϥ���/�n���u�}k/���{�7�`7X�������������"�l{�~���i��a��$�qt�iӦa�ǎ�`�x(�	�* S8��®s�
�%#�	b��z[_R�M�Ӵ4Dh<���`�ʟ{t͚5���Jg�������1�X"y�Eg?�m���]'[6��כo��sq?��7m�4f�"<(�̜9����F����G��d6w�Ek��ٿ�+?KЁS)�����o)����'��@�#J�L���"8�D��hb.:�n͌�)�$�>?^�f��"��@i�h�ȁ��gφN����'{z�5U���x�g`0�iԎ�S&P���-��>�@LbX���h3�5��(s���?��õ���w?F����>M�`��380�K�x!��-��C�!���h��s/8�-���'[�"%��qTZ�;l�\:��A����3����T�� ;���Q���,cRd:��nUL/W��� �
M��^M�b�u��8_�K8�to�O�t���le��t��T���c��P,��ˠ�Y��o�X��y�S�T�C
G���A�
-��p�%���pxl��H�R�Ik.�F�����Xj.��q�I���KZ'Pm%И��LP�O.TV�t��{��o�����Xv2v�5W�s�
h�U�t�x ��)��Fvo�C�C�d�����&2�eɘi2�.	��Gl
)�I#E
w�*kR��@}$^���`��R��� �Bױ)���J(�RrK��B半��L
1^wvvϙ3Gw8�̙��C����B�dNM�h6��M��K�J�Q�����I����a�O�>UM�7�3NKAC`w��Q^�r�[᷼�/
�%�fsJ *�m����U\r�%#�����+����[��SP���s<���c&'͟?���^ Ǭ��$�a׶o�>��G_6F�����Ǜ��PF�v�E߃�>+�N�a$�bǑT�4b<�W^��J���	u;F�� �����Zꑥ?qM���삄��~E0��$2�+9<~�� �`&6�m�u�wP=:F	ۙ��c�v���0�Ce�o��6�����4�kޱe�����l�[���B�*v�^X�>�I���P�w|W���0[A/S�"�h?��N�O�=��(:��[.��+V��ͷ~��caQ<K��m����������IfKV`uM%!���Q�5�� yѢw�]��
ch����}Lp- ����ϗ���Ա�cfu�`�eϬ�򩧞z���={�IBo�g<+�Ѹ8�%ʪ+�em%6g���p=1�SUS��+_��ڵku���k�����P=o�馟��]����Z�]��I�s�N�	��G?ҽ��w�*��n߽��.�8y҆�s��xnWw�ƍ[g͚��D"T�E�k*E�����?����<�G��c���ga�3Z1C���Åx�R_�AO�w!oƎ���0�����k{��_����x	��i�7��(�P�:�{�n�r�3����y�|<<<B�C&�y��D�M�3%�_$���f��R�,�Í"���� |􌢟����PD��>PTmm	F���R�R5�K���J�<%��Q�Ȝ��������N���0v��h�NPH��`	$�~v*��NN�x��i����r�K�ˡB�WWW�5�uu~��XP����j��r�_�S��-��
,Φ�8�K�,y���{G�墘@��M8-�&���bH�v��2�0�VB�S�o�"��L�߲�p	'X�#<���MM�s*�O� �Vܳ�z<V��	�9-H������yH���� tȎ=���eVN=�lTC�a�]|��?!�ߺ�bo\�+�6��iй��!Կl!�Ǫ�c�H���������Нu�f��`oRIvPQ�0C��NWYI(�u+]|�y����ضmKg�j���*"���_��SO>���]���7
����z�o�i�f~���t.�?4��e�f4��_�t����AY��;�{@s��*W08�����&hz���vr\cᘺ
�C�+!� +�e��Y��Etz�-�s�u�&�D�j����e/�y�]�;8��C�#�@0�90P^^�����	����5�#��֖K.�mv���3�,/�'�S�M�<}�O��g�z���.Z�d>ɱ���̓�?8a�d��ꊂ�fqLDB���$�M&��2�n��hWf�J'��t��p654⨨E��b<X��gX��j�!���tls3���S�nڰaӺw�Xq�=�@|���[[[=n{��Y�ē�P(TY^��#�Ǹz��^z�/yI}���=���f@��w�ZF����p�`��о}B�<K�9ݺMw��FJd+���B)��H8\_[s��gL�2edh���bݛo��h�/:N	&��u����Z�yɒ
�B%�EU2�*,:=�E%���	�z��u���믻�:��f{ 0<<<c֬m;v��	M�7o��w��/�
��iw6�5v�uƓ�?�������?7o�YUW�|�����_~�p������G&M�z�m?���*��2Tn�q���a�G_�`v:�@����k��f�V�,v�g�U6���u�]�CS$L{�v:�N�R�X%�, t�8��=tpo.��I��/~n�>�Ԥ)�,�W�����}�۽\S3t���|�s�}�ђ��bܸ1mm'KB�'N��Ir�ɻ��{��5�U�e-��0Δ�KJ��4~����6�J��k�+���.ؾ���f���<��U!h5���B�]K�2a�Q�<T�0���JT����"qv=9�5SULJ`�ws
���������=�*C�\ZJ�ș�l�U�7�&� B��TQ/��J	�v�2G�cJ�n)��Yʄة/e~xX)`C�jrAs�A;����t�#*�<���3�x�;��t

�T���'���
,2��Q?�K���'���쐵u�5���oܸ}�V~B��G������"Yy��͛w9]vS�E�ô�P�� (� ��$��>G��X��>� ���Ǡ�nB_n���gsɑ�>��VRV�� u�!�w� ����*vN�g��. -p�A����n���a��9o���Zer�N����aѹ�N�N���?�R�k�)|��|�
5����Qpʟ���3����P�X��8� �1F�Ɂ:+���|�-$�����a&J�����o�4i�dC�������`�7ޭ('��D2���*O" ɂ��ںU����0w�ܙs��J;��奄����	˸��2i�ĉx}��a<7#.�_чYQB�%1a��.�	�3��XY�V�,Ƽ�UUe_��`�oز�cSy)t�}��L�>���O�����93oS�Բ��+K�,{��W�Q�ȑ#+N]��/~�Ku}cwwwUU�����01��/^�x��)�<��~��;��m�J��#�o� U�a����\�/���Rd`G�P�&:��9�}5<*+�ꪫ�G7�x�s/���TRZ���/�˰�׭[wϽk1��>B ���܈t�Ǝ;(1-E�W�S߼y��.>ٿ�Ā0��	BWW{���	l��bb�"ɎN]�`�c� ��e�D�	������`��	�K�����FP��Z#�n����ek�_Bk��+��1<���V�ñf��-����C���K�-]�j�w�_�W6m��h�-ǎ|��/	P׵�����{#���\�l��0�9�̢QjC�\�tiV�>�u�V�&�M.�O�u��Q��hV&3��v���;2��L�?�����~z���� }T�&A�K�J��A0��_|[�a�&�[��~�@���<��L6X������B���Kv�a�!1}��z!/F�"��\�G��E5u�m>��g9��Dc�΢X��r���Ub�06-���M����!cd�O�$.�7ŷr�8��~�W8d.�?4��Y��YVV��P[v�	�R��S
�ש�i���ݎ�YVV�!T�H���ː���Eٿb��O�ɒ���b?I�L����Ì3hT�̶m��a�y�BU0Y(�PU��xw(x Ĭ���yZ�X4�-�E����P������	Ȍ��U%%�x"�xU���+�&����/��.f���EP8aD�y�-�����H��>�Y���&�wk5x�E���#X?�R_�4��%�1���iI���,���z>FI|�x���v�'�_��29�5���Vԏ4�B�L��h�+�_��淪ku�T0�J_|!���?���9��ݮ͘����^UT�r�w����E��ӹ�K_���q0&O��HM��S��{䏏�vwv�I��rͥ�^z�h�{[7C�L����ut��y���	�U߸抟����:dw���V��Ma^�|��fy�⡬���1Q����-��Mc�x���)���>a���?~���z�F���x���k*fΞ�������}�k_��w��yㆇ���<�~���_�2e�;<߸��}0�Uu@kI���q6��<5ee�@t�O1�!��,�����y�`���Н�O���i���T�?�;}�N�Q]^q`�އz��ŗ���[o��r�Ƀ���t������}���ֻ��t�.,�����U�յ�C	�w�>��w�掓m�^_`��=�.��N�fEY�Qn�[ܦ)��NΔ!l2�S�L
�(��-Z��6B��l�^x�бw�}���X,�0�,B�bё�Є����*���U�M�Ꞡ/`4X���������c��~�u�yL�L:uV���͛6Ak�����{��q��ɓ�~wӂy���o�V�;z�i¤�~��P��op�杗��ƣJW^�fl�����o~���;7��U�	(A�<ng2��l���=}jY�?�4��`�>��
f����T�{*D���K�y�B�/��k����r8�K�r��Hn(�I��B��ax���~sƌ�П�����0���o�������)�UWT����nS��@,|g�{n����:;�k�3�I����)<z<m��b��N���xR6���b_�Nׄ��Ue����Q5}_o=��p�,.'��훣:^2�a�044x��0�)���vp������+[%9c�>�k(�<��"Ѫdz��d��Ú�'�>�	a�k��G��J���)�b1gT D�8ky�fO�i��鰫
�G�i�P0TU]46aBs}}m,��!Tr0��	-lFH}��@T>�vn��/����	����5U����L֐�,����J�#>�,prL�e�w��4qzl6���T�U�ʰ��1�7@�A^t<���`��8�75Ԓ��<G&b(�ʠ�=�O�A�t&eP�t�6���6�+��;.I���dC_�U�ttt@�d �\V�aa����tx)�AVxe����򲒒 �[Yר���>�R�g{����B*�ʧ;���|K�s� Nخb0g�BI��E��XX��A��*iŃ��T�F'��F nK6��IQ�������O=z������k��\�pʔ)~��X|�7nɒ%��kk�0���o�u���������X_�򕠏��> �T���\a�#�O�6$�ւ�bm��&�6�&��8tb����RF��W� �`^`2��UZ���H"+����2u�i<��;�9s���ǹp�{*҃M�޺=�]v,cX���n�����ןq�G���d��:���A�?��Eq$h;0HP?���"�E-�t<lS���|R���E!�QřC_�!��������-[v��7C����;{�ue���7nt�]c��445㆑X�j�d������G���o���BO�x�PI�$���L��'�0E�'D?i�F!-����jk�a|H�$����;�0�����P�L{r�+�!{�~���ho+T���[VQ�/b��$���ׯ��j�fg���n�6ǘ#�pM�¬7�޼yucǾ��˼��=�؁={�<�L���������0������d���5kV [ñ|��5k�ԩS񭁁l��L`�6ۤI�p:�G������3�hC4���%@��d�eS��&�<����9�ֆϏ�0x뭷��ߏG���ol�>�C%ص9����VVW�`���w�SO=�o�ZpL�pN�LE]#�)Ed�;�N�OD_��ōᵶ�rpM�h�c˫a����c*��|
�@T���V�7�q�z}�e�~���xS���)rz)��p;��'��>���x�΋*@M�& ,c��p������Df��ݐC�8�������0M�zP�K�iR�w���ȴ�N\Y���w�� �$�#�(x3C�c*��fӆe�[O$o�@5�E5#�
fZ�'�����U,��kd�� �IF8�7L�Q.�G 
�n{N�U�a[�RLD>!�4������n�f9Y/F��l���rB���J���w�bJ�z}F��U��\�Ў����P润�|O�c�ߺ��׊H�g�y������Qx�5q�����D�%9��v��� h�G2������z�����Ԝ���`wgO_]ei�{�ޞ<a|oWo.�Ԃ�b��̪Ug��.j54<�"����a�K/�TZ]}�i�-Y�x�I���'�'2io0`w9�^���}�A�^V�8~LSmeE��-��Da�ي�CV$��D����]�̛��m�ĭ��%��;~�J�t�s���T���w�h�,+	���z���~�[ !(
Ҵ�d��zȒ������ܲy[���<X�D{���{o���;�,9��ro9�b�i＿)O�Y*�����p����^�?��(�8�9����⧼���p�1������T*����~3o�M��V�D�B�>��;�����������t��p�e����P ��P�'��MIy�ig�*-y��|��W�����яo������2������gϞ���AUI9B�$өLk�M�GÁ���m�">���}%0��q<��)B?"�� ��^;6��r9�_#�- Yf6�b��!�p6)J+�p
^��V�'&��$��b�'[K�%�-���N���/\*����[aa>��K���/���M�O�"�xeE��:��?,V�	�v�d'�'�x�#��8n����MN���� n����%^��Vu�O1��S`�&`�̜�9�4����dϳ��'�����/YX^]	��-*�;�KGg瑃��8����^,i42��dS��𞃻�'6/X����7~�{�&�`Y	UTJ� Y#���o������n�|Ųʪ���6�x�t���mhjk9i�/�$VDf����8n(	̀�`8אd��E#���Pz4�z��n�T%g5��ͨ�s�s2��Ϯè�|�tFl:c�,��4�.l	h(k�H˂���)�b�*�J�L�,׈�6P�=٩)V�55z����jkkE5\�"SN�](�\�er���j�:U��:/8,�Y��S'�}#M��rA�a=s��aѥ~ѢEсNIh�t���;��^
���ͦ�h�T��+������
���KKC=�Js�4���MΩU5|�tk�TʕL�!8ľвq �XJ�6d~�x��Y�� ,F�A�D����P"sSÑY5�K'A�B�"�.��4�ϨԇT҄��茖#:_�X#��{��,"8d��J�:��N6:��\�E��#���i��E�j�V��x;E�h ��}��͟/�`J��PW��o_&�Ѓ��OeT�L�M�k������j�qz]^oOoOyE� L���~��|�`��N����4����կ~��=����E�j��׿�u�nB�H�5�fb�h(�r���(���'ԯ���Q��u;v�X]�X�]NeL��ϣ^�fux�����oH&�
,��7ߤ^�/�����29
���C�A-��[;�t0����U75=�ܯ���/�u�]�\rI*ŝ��sQ=�)a�M�8�ˠ��'��
lQv%ҿ�����,f��R�����=cƌH,�{�����vM&�}�������>�x����BbEc����A�8D&��$��8d�v��^{��p	)[F��$�t�<-\�_��I�ґ#GDu�L�3	�a�������~1���F��R1�����9~�)`�p7g܅��ڵk�ʕn���pO���_�<f0����Ҫz���?�S�/���3� ���ܯ���$:��Ý8q"o�,-P��P���Gޚ�n��\�s�q�� ����"Z��g�{��qUK*_�kM�"i�k*�tS���͛���/��>r	J�4���ӟ{�7�����f���O3���%/pˇ^�l^,[��7�IP�Y��q��;]����8�G �Q���3g����|_Ěȣ2Y�H�4��;�"�bhtO��	
�L��W�F����%&�1�p��8ߖ�wCi�nJ��vC̊;�3��L�fv��3u�*�wp8lb�27}lP�.�T!��Ҹq�T8O~�:egrbm��7e]D�����k���L��L,����f�͑���K��WCC(ڭQ���*��{�����4V��%��=�wI�*3�u_�q1!]vE�H��א`��t��a蔹���ck��J���￘����f"�l����q��<kܗ����9�w7~�*{O��V���p�w/K�M�:q�C�p2)�W4����\^$/���A&;�$u��b��k��e���Û�'TX�ÃC���O�M%sa��Fӹ���O���6sJ*�2�ŦD�QE�*�>���	Z��q�������*LA��y.��ϟ�|��F��O<�Ě5k.\}i,��K$��ZMJHJzd��k���y��l�T�REP:6 ���E�j8BnW(Y0k�����[o�ٳG���5L�o�YQ�s�o������,i:����vde����Gb���H�b%&�"����A��#ɰ��4o���L�iom=�n��V�	�待��߼65����˺�����ox�V%�	�Ē�',/	̔tu���r�b}û����?L�8y���Ǝ��m?���Df�7�z�����5W_�lɬ���`/��\>�l,�����@����:���e?q�8��W&>���'P�7�]bj�58�##ófO��N�qt$�MJ6�͕�&[�{�,YRRV�v�����^XSY{�m�lݺ���h*�ⴕ[�~mRm��$��h�i�t���&�`N_o't��W_��#��N��<x�dǝ��S3n����j�q֩g=��S�T2s?�+-+���������v����+Kzfd8���4���f!�@[IQ�V@0M14� ���T���q�v����65�zlv*6eꦤD�n0!J�}��H�����!�͟M\Fӝ���z���n���/��o~ﻠ�ŧ��ׄ~��}c'�Y�d������;PWQ���ƭ@Æݻ���$()���b���sIN��"��I��P�o���:K���+g�G�]~���_����KX�WT��-T܀ncٌ/X*Z��v���(ٝ��e�d�l^Og&��eݝ�y�Msv��}÷�����.UF6{��N���������?��W+OY��-��e��L4��䚒
���{w���s�4毯��N�%\6W�P�SwxS�j�s���f�̉�(��������ϟΘ=���1��b�(d��`/$���+��[����F#��\Z���:��lH���;]%o{g����)z����9�'YV̌V��J}�e�C�!Ǔ6�*�{B���MdE�b�4D?�J��!izdp۰�$T I�8�l��S`<T������q���?~l�pO+TC]�F��S��.��p4)��VTL!Y���K�E�u$�Q@c�����ΓůP5+$�I�Gմ�B���P��!�CƑ�G��O�T^]�����ʱ��=ʞ�ݮ�\��$�m�gi9M�HYQk �n�N�+r)�"�V�jkJ�ێ�jfn�\E��
�F|�m��@^� F�Udcx������r��%X�穷{�W��`N�&�v�=k��?\Q�����֋��U�Px�c.��5b�)��| _�5 �	���U}]��T�{��+�������yYh�'K\�ˆ�J�a�m)��i�h�QF�R�]�>���6�{�#��E�U��<�%�8���8���@1���ו�E���ߟ1c�D.�ݮ�J�����s|w̘1MMM�6�w�T]��xS`�l�+�1��������ڡ�\�}}�XN?%۷�F8�:u��+V�����m�R��)��Ds�Y��s�|'f��E��^H� ��X��42��6n܈G\|�ż���xE��w��	>��3�L
6�ҥK��Z�`Ѡtc��4p�xk�����	#�8��u�=��'ϝ���1_<:L4H��p/4Y����M�[k�oA̰)̡}�="E<*�\m��
�a'��>f�q0��(��vc���<q�E����ϭ����[oA�7iN�=��g`ʐޠ� �An���x:{Ǐ]�[��֪U��/��:o�J�-�����'��6yʭ?��F+j͍\�Qikjj-Zt��1Mw��!0B���J1Eo2y3i�I`Ȣ��0�8���A$AφbpD��/� ��#>����i�.Y)����~�y�[�o{z ���X�n�! w9&��{� &@�`��P���H�K.il��Zmݶ��_4�Se��z�/����c�b�u�\��&F���0և FɊ�r �C㱎6�e1c;�"-�|�[V�E]�o���(a�<�L���BqC�$�M<�r��Z[[̜�B{q���'N�"�{ �{��*���jʜnM��M�R�x}}}mm�f�@�����LI@������v����x�tV3>O5��=��U\v�;*���0i�n�L�eQ�Q��8�d2�2��2}�R�?J�8���a1�e9$�t�"�����(I�����na�S;�*+���텕>ၰޱln�a0��D����uR"���
�x~¹K����+����%ѡ@.Y���ç^�'�ĩI��J�(�#9l��9/iV�&WG��o���p���4j#�<��Bޱ\LaI�1�}I4�%��R�߉������֐E���ʮ�������{��"�(gQ�bU�@@]�f1��ό���S�Z�v����%F����b�'���^v����G����̙FP|`�Ixgy|����bu��}P��*#�+������iE��
s٘Cw����#0:�`�@iY����`��t}Ƭ�A�����`��z8=��Fvye���Xk��i�Q)0)���*��eԊHD�Ă�Cb���{��g��+�g~��_̘1㦛n�<y��_�χGtrF�1r(�BI"oXCC~��rE[g��;!�������������<�5���ʚ�r�ܳg�{/��GWU֑�_�j���N�is��5Fb';�U���%^o���`�r���DKV̗30�K�&�Ě�q,&va8.)+��9p�4�][7׏i|�޵�~���_�aW��xFy��I����SD�����K�����tEE��?<2~�8Ȓ��Άq�n������5�/ZmJ�t6i�r!�+�?��	궁�^�ފ��b�(6S)�CL'/0�!�y���\�#H{3�{�aJ�P5&0N2F��*��mp��ƒjӘ��6l�Db��*�����lfۖ�cǎu���7nX�l�?׿���s�������W]s��K��l��]�vy������!�Z����ګ���sW�{��ѿoXw��!�~@u����nj�?f����s���.�3#x.�NF�0�X9���.�� $�J���M�?f����d��n��i�4U։��� �*���)/����ʊS��"�J�`�N.B�Hܿ*��&�P\��d�WUk9���=�%��Z ]s����{"L�F0uq�M�i�Ғ�B �f<�f%b1�M�\0'��C���L��_\��-��EXu�4�/��P&����mH����AMI%�C^�M���d蓣�N��
�i���`a
��b|���.ggO'�h��vy�(��1�1�?H�AnQBN^d����X&cX�f�J�SKA��c
9��{ج�3gcv�H�����/,��?���O�_\��S��L�v3��BM�"ARA<��g0U�dO�<�6�$w�h���r˻� ��x0�,�'�w�#�A!�^O�5��A��3+�%�)��p���Rld���s*8qބ�t���e�Ĝu]tڶS����@�pXZIEa��ik;�����l�G��?���I}�R����ڡk���X_�e�N���`��ei������r�W�ؖ�%թgs�Z*$��_�B�Ǽ�5�eGNvp��V�z���O��+,��:g��4�ill<p`��m۰UӧM7��`� �N��T9Csڴiс~#b��ջﾻiӦl&5w�ܕ�cxm�����Z]r<�rD$��Çc9;J�V[�,�%y"�tYѱ�L��"¶`HTf:�!��޽{�L��A/IX0x^�z��	�w�y'��� �)���7F����/�lڵcG}m��g�����]&���;�@`o��A[[�y_�<���-~�g���jB�Uo�w��:nY�F��7Flу��!m��F$r����Z���e�Ūhܜ��9��%L�����������[n�奿��{�d�0a���f�7T��vϟ?f.,ZBX�-G�i�������7lؠ�����$H��"�C�du�����߿��3��a�y;D�;O(���,�-JE�'�-*e�S�V@K�]�W_}{�]���_���!H���:�<���ql|��������aSS4*�M���9vҤI�fL_�|���N��-[��J���j"�8�?�5k(�S#D[�|�PlK̈�Q����HL�V����:�BHH�(���͙������愹;vl�Ν��58q;��:�^cj7nğ��c��e�ۘ�Lؿ�}�駃b�˪�o�θo))�	w����j<�:q�DD.������Mɲ�N��� v7{d�!���<A���N; �a�s����"_�"ǰ ���ĈD<^D�E��):+��$et�ȋ�d�32��NT&�Q�pu�DX���,�Nΰ�+�W��>L'\�P.�сs+��1y/�B+2Gu��.���Tp��}�H��]�0ߧ :�F��e'v����L$T�,����L>V80zl��)<E��^1C$A�� IR���5!�\�7���+f��"�;�zl�P��r�;_�C;�Ò4��I��l�����EX�;��3'��Q��hym�����!��,�``[�;o�ǔ����>Iݣ���J��B���hON�G#�$*�*����۴d:�����H�iE�9�v���v֬6��@�M�q%踀$�1e�i�NC�tuu?~��q��Ř}����A�.�R4L,S�sUWW�`�`(���Ύ�ӧ���n��w���;��������1�X^\7�l�hΐ \;�9�e�tI�-wJ���`�a"++�8y���q�=�̘>���Y�n]YY��W_�����կ~������.�1k&�t<A|<���]n�[��n���'u���߯�񏃇|�o��{���:; f.�W�аs�����\y��ɑ�>�x�^�Wѩݭ����w����`23���l9E��egG@J�$�v�>���s�|ʻ6��3�]r��s��|�O�h{��Ѷ䔥k����n��k��f�Eæ���c��aÃ��Qj����PϹ�F�K(�QzTҕNA���S�ɧ.��zhﮍ����<y���J�4��!���-_�������ѕ��.Z���]?[�6a
�D�Ϡ�5l��u{�t.k@�Y�T�|4�JIF��ew�} ��.�������x�?�y�\��@�9��ʅ^��?�"7{8<s��D>Kp��(�Uȶ3�����ӧO-��*L�qS)��m����`eЯUb��:�x�ԩ`��H8�J���\9H�Y��f)�B����2��_0VP&�N��Iͮ��$�LJ֑��i#�����$�*)��Uξ�\6uRt{r�:�d<���{��t��r+Ξ=����#��z�8�r���px�����7B��{��g����wPWQj�Ƴ�)G�G�+T�W@���.g�2�]��I�`O8���X�,0q	�8��"�+/0�
�w�1�BǢ��K�L�x<9<N�S�4���Ʃ�����9nrRJ��������ϙ�tB�<�%�g3�\:C����A�빼�ΉҞ�K4Zt������j4/k�b�d�r�q��ʧ�����dC�������_TLi�5�[~p*n�PQ��8S�]�Î-K&�CC��ӥ��%����O;�5_��[�����LXc��`6�?#/��{ysI=烩�(_�'8Zj����bQBK;����JKK�rU��<S�b��L.;�L�s�2M��m�A�Ş�2�����+��1<�M'�����8�&�D (Bkm�A���\~<Z���������2"�T�4�Km/*UU�azP�p���66��|1�� �?e�lb5A��"���R�.W�2���Yr 1���H"`O1T��E>:>ia�Y6I4�P�ݞ��t�����"�
t��c��x̀2��.l���]��:`+�M?����;ԇA֏i�h�#	�z�bL��[�I���T*ɱ�m$<�Nr|�'�C"�DY҇���~K�;������1��\t�E0p���w��A���*p��*a�
_��`���*wwt̝;��瞃nt�WlݺV��SW�%���|睎�.ƞ�E2�
�&�'r,`D�Rd+�06W�6�pqF�1�J6�� :�2%�Z	Ҹ3�	�V{�̙�ǣ����?<w�j<�w���vʌ0|1f�{JA� %%l�㹰�Ɍ�ȇT7�9�L�NwwowU֏�G@�=a�H3��[�P�[�,n�`�(dJcA��p�lِ�O�jJցg�D�z)�E��dS'��(j�c��+)��ꫧΞy�ş�?��OA�S�N=��PP�W�!�c�Ǐ?x���)��!�? ��N����A`)He�6��o��=�E�e	�0 P~�:�	�$�_��Åw`rFK-+�Q�V
��@Ӽ������Fڃ�!��ٳ��<��77�{v�ğX��GQl����ի_}�U���;�"?����I�'cS:::�M��HR�l�k!3f̠:҈�*�L��D�7�v���4��<�DoCa�����CXg/�)z�85a����l�a�R�b&Td�������L��&cPJ��.(`N��Na廝��99\rT�9!�C�h�Ug�JMZ�l}����+T����IjO��Ώ��G�|K�[6q�,��X�ӖK5���
��ZΗ��͕Q��o<BQѓy�*�9�K�M��Q�D���qs�(�zC���IS�5Nȸ`���]�rIɪ8�E�8L�pDR�g�D���q`^)v���ĕ�����ԕ#H�0KK}39��7�A����MS�W�{�9��Z���X�}�JKuM�(�\_nJ�hB�3��3�?�ʦSaOf��R٥&���\Ȁ�c,(C7MBN�;���`�A��} G#g�q��|�KR��3�P<n$M*����رF�?X�A'R9E�j=�X�9���@(�\����Lw�OHӿ����=t�����n���/:�֖�f��G�H<��7���m(�\�ʋ@��'�=+�*�%:*Y��I���n}"P`��c�>|(3���O�2	�w���>���Bx`�[u����kj"J�F�ÃmV�!	�	Tg���e�����4���o~�����%��x2��𡡑�=�xz��,a8����ʙt�2��=�x4�����@��V���$o{������8�.�+�9����͝�k=�yӆ���<��Gw�R��n����}��3N{����g!�.]ZUWW"�(�ץ�Ix((
�H�-V�vQ"?4$ؐ�{�T®�[�x��۫����s�|.����k���3f�k���`׾0��d2
1˦��.�V bTD�$A-	�H*�.�0��h�QK)G���J�\>�/*)���'N��w���3�?��Ѕ7l|��K���w����r��F���}�?o���xdL��G����fL���X��#��5��u���9�+���:t0v���r4VV�tdSi�M�F"�Hd��9�E��=ð����������.�1G���H�&�5S%��#�3�Ι�q�.q�$;F�tJu�s.��导�
�K��˗��|����pd����C�d-_���7߄�7v������5�O�`�-8�d*�i�iӧC^|х5�U;6�{}uU:�W��&]�T}S���̭u��������{@B*B��E#`v��	)�F�h����$d�%lJ�.	�G	�n��%6�x,�����fTnO��v�S�h�ӘL��A��r�{^�����uG����`}z<�<J����|���F�1��CASej�@�>LZ�, as�X$��ȣ��O�|����B�X����l���4�!|$Q~Y;q�d�{�S5�~k�i���(���&�\N���	�@#�K�ל�AAaD�*��bU���(@�VE�P�JP�8��'O�w�`wW��hy��9�+��2��U���I&�����84����Y�-����a�P��XOg+�xM#G=�SI����He��m�"�ޫ���� �����$�1����RQT���d�O�t_�UQ���d�"����$a�W�$'��$p�29� T� �][[˟g$T��c������SO��W�
�m����J���v6�	T�?�R�n�
�r,x��o���ys���*��]��iG�=��#��
�җ�dE�p���-Z*!{"��@��!�uZ'�!�[�$��G8!�J����R+�oJYfCf1�W�X{����1�w��	�@Ⴡ��WU��lQi)�:ȃ��ׁ�*0�8���&��SZ9m�4�d���j�&M��c�Ơ:������{ ��v��fw�}�z�0SOus����frl�s�8�N0X�v�|�b�Ć,2
9!��`���PoB�z�gJ<�P_�`�3O?����x��O?�y�f�������f`�C��v���b~	F��_�!����^�ӥ��8��Ow['�Mo�����vd��*S\�Q��޺u+�!�$͚5���!��P�,��&�2'���*�f{�
{�%��|�M7a�o�{��|��ڴ���^�fͮ]����8��֭[��a�� �`M��-��}�*QMˑ�d��� ZX�6�w*ew��٤��d@!�����Y`cS(=��8q"TI.��*s^:�V�*�R�a��`s	�Q�XBKT�4<g�x۷o_gg�m��c�� �x衇N;�e˖1x6���������k?~������|{^�qϞ=�K�~��ݠ?FJI��nx��?©�U
���2�w��J����ae ���T��п,��y�T�.�&/�m�e���L��(o��h���S ���ے�'|OK� *J����S�Z��Eq<0�v����$%����Rߒ��G���bO0L.��dsI�1߾9
^%_�c!��4�zz~�T���\��u���G���E�,��Er���̟�*��0B�����G��S�M����C�6������'q�1��l;�ݤaH���R��T���!iEFăE&|=Y�]c���d����b{��w$����j��y�bGGE�tp�Ϣ����ź0͂F�������;Ǐ�
�F��0��AʯQ�2��֮X~������8����M��_���3�p�bi��g��߮o����XpSԮV�+�ˊ�~���f� 	RUKC�k�r1�1$�����l�,|�M�8e:�;Q�d�Rؗ;�nq��F"�mm�AoPM���;�L��1���wX�>���D���@VEO6]'����G֯BH�0O�l�3�+	�4g������
H�������a�x�c��@xb&ǎ�,]��P^^�8~�$�,$�ڻ�>�3�=��]{�@�)��!�U� ���d:1��R���n��
�Czt�'%������ͥ>�����?�W2�f��[	m}����G�!���1rl�TTU�����[Օ7~��P�"��\ :ٵ}�nmu]˱�Fbx�ƍ����?ܿw/�c����1�	���d2!�K�aw�:�i?)p��S&�=4���ު�ABE#<튚��fmپ�����m�\n������<�T��#Lӗ_~� ߾�����kc/#!�hl�۶�2e>C�N�Ԡq�r0�*��'͙�0~�}��~���뾺t٢>����[������-[.]F�y�x�ֆ�c�q6n~�/���~��N�6���]S(�&�� -�+�'w�~��ǱES��I�g	8-�L�>1X[_�;<��p�g %�,���0d�*��n��E�Fg�'���Ѐ��������n��K��|~���L:�4n��h��k��jP����VCik=����\�O��r���A�{��3w�����8TR.s��o�#�3s���ϯ��k�6(�_�����ﾖ���.'�[䇫5Uե�`���TV>���](442�;���=��`��y�Y��$�!D��,��y�_7%�`o�d��@)/PTv�Cr�W0���UY�?H䫰�S���.ψ�KD�2���e�n�Z^�D����]�p*i&�ьʹ�m�4>��-6s�ӪfK�R�x.uÙ��L6�L��ܦH��K5�~�Db��d�TĐf`|� n$�ڠ�%9�N���*\Y�D.Ves�5u�3�e~�/"�R ��y�إ�B��0*��@ʌk�G�:{��j�'	h�U4�ÚD`��	����2JG*�r�좉�1q|�����H1��0��Jz6C
:���zAF�m�`�]vH�J�TI���I��'O;������L�u-rli9�
�ֲ��)
�KH���bPL���]<�%F%I�����~q�6v9�;� j�����O%mYу�n0;N��\;$��&���a@2q��@�nX���;�s&�� ��2�h�_#V�\�
U0<2�Ά|,�t��R�˕b�fM�b�e�0���:�v���p�D�>/�R'c"T�K��ƨb���Y�}���SO=���/����WlXc6%G�	+:A��D("���#�7o�
���P4�a+'������=���J���k����9��w`?$�+PF8�����FF���ٷc��ʯBc��Ǝ���yH}�+ę;�m�*���a��_ZVB�	:�"^C16X����֮���r����+KCG����ri,����]�����;x�`SS4}n�)�LԷ{h����~�ܹ/:ZNBc�=~#�	��~N4�9�:}1qCR�nq�5��]=���&a�u��r�G��L*g�����7d�IlY]�44��{�ӦM�;;�m�<�*P>�U�	�A��Ǐ�R�'�~�W�z`�$��?{�l�#�c6M���`�f6�;�\�	Kq��a��*xða��Ģ�H���Й�ӓ¯��\F0��K�mZ�
��a�hģ�<�p�I�㡈�d�w/���������������+��o~9��� h �1y��H�Q�$KZ��$Y����v)��岽k��.�E�T�J��uiK�T^R��I3j�8$f�AF#u����������������X�-L�������w���?ŷ>���al�~��q/��5A���ǟz����PF�x�	&���G,B���'x�!��!�>����o�y��B�/���syp��I�T�E��ie�uQ���V�Cb�%@��u��4])��?TxG��m�G�p�R���.��9GVf�[�%ge)����X>Z*��ԽD�{�gI�.�����h�t��L��^�zs�3yWj�����N~��k�)[�c�3}��9������ϥ�?��&��I-�����W׃m���y�C,�
�|��c��Ju����΁�TkEf�`��	�ށ&��jY��Pk�-��.&��B<F�@��'�29��<(��j�_��K'�=7�ԫ-N�V�rG�P���
q�<9QW,^��C=�"�8�q�~������vŦd_|�ࠂ^�8��so_���ih��n֞`�c��<���7Z���!P��(V�W9��-U����	/{��w>���N|���zkm}c["�q��[oժ�)�0���m�>#C`O��۠�Օ�B��������e!�#'3�	�xY#'[��2�y5���k=L�݉�?)~�B1�S�3����94�ҥ���w?����?.����*��`p�JM�Ry����@�3?�7���{��W^?�|�P���\��ȏ��O}�C�FCK�űQc�lD�}��a�๘����C1*�Nawc�nͩ��g�~���t��Gz���-ݺq�˯�~��|�B�|۷}������W>��=z�慭h����������W�[�]<�Kv;�.���7o_����_klCQ[[�E��ѣ�'��j�����up
��ha���%���5'Ꝯ�.lwvY� ���PP&�ſ�g����{}���~{�Z��r���ve�ڱ�<���z��҉��7 ��ˋ ��+����ϯ������O��w}���;p��Ͻ�[���������?޺y�L�ܰ+ޯ�-�*��IT����_�����Ԑ�Wgb+j�;N)�Y\l-,l��� �z�����aX1Ѩ4���U�A�9J�nvv�d<�kgk��5���$��	�e��#�?�7Q�[�h�n��~��>�O������܏]�V���G�,�ׇ���5h�t,s&yP�~�&��j���?������sϽ�8v��_��s�.�=� ���fCכM�����n�tn�m\�q}�ם?4�x<I�pWYA<�lm92E�����ݬxX���`\���x<,��ZtP��'����"* �8���-(�+;k��n��y�T��^`�E[�{�֯Ǖ�=����n{7�=<Е��[��f�Tʮ�o�{�!tt������n$�Y1�z�ȉ���I~M��;n�L�Y^����fͱL�f���^{�������[����DY�A!cE��O�*��p�[4�Ѯ�Z�b���������¡��IHM����M��T�H^؞��f��B_p0hܷ�[-l�;35�kk{1Ѫ�d1G���m�A�b��#�*B޸}��qsg��;D���J��X-����F���C��@y5a�H
�$f�{��$���I}Q6��J9ոIy�n�:.N�� g�{�K�>�$���AP������D��3Ua�)� lh�8��o���ٳg�z�	3��>)�)ٜ㭲ң�v��{Z���kۑ��`_޼y�2�"�>p��"~���s'tKW��j;lMX3<>�4ZP���(���~� �R��ѣ44Ce�̺W��A��d.�����	�Jw0��D��]�1r����0qm����6^���SҒ�13�С��G?�����]���?�hԠ��+�b0^%����N�7<T�4GI���Sx�{��/|[K�I9�z�z�h��$l�k�%?8q�ă�>��=��#��pgL'|qq�q�x���D �����w�k3��6��q�`Kanݺ�Z8,}J�W,��;��{��{{����|]�#��X��������@i��c�TD������c��a��k���'&'���`ʕd��eIw����Z�?����+XdK[�Cy�� 21�;��9y������7����չ��l�8�(��h�xcC� �|P�<��Y�����⽀�C6} /S�V��|�OSͺ�
�E=ˮ)�4��6��>�䓟�ԧ �?��?���������w���������X(��w}�w������� �c���A���������5����O4Bi���#�$/�XM �ؾ0�]3h�:�ML�1�X��k�7��mg}/��8V{��a��8��6=��"��RkZ��q����I��;�������Z��Ys�;<����ÄqN6ċi�}-5��;�¢�>+���0�;�'�m}����~5��ӭ,	���9�X=�E>TE!H�ۃ���`�����@kt��gF�v/�r��(HI�R�+/�l�!�4T�W֊�z!���ŷqϝ]�sr�������w�WO7�>�r�q_r�W�����R�7X�'�ϖ��"��N'E �����N������wQ�i��c�	�Xk���8�F9Z��p�B%q8�1��QTP��r�}A��hk[�@}I�)k�W����ͭ-��k�R߉��5�dҏ�1����ۛ欺%������g��7�:�#�H��ӚhU����U�|s�*�i5�6��`(�c��.a�/^V?j�����AH%X�g8��<q��;��ࡎz�����N��mm����jI,9<�=��+gϞvz�II����V�'��z����N�T����x��G��s3B�n__��G�:�
������vwg�~��/�}�?�t2��J�N��2���D���`cj=8t�gjr�����I�tl����R�2;)�o���>!.�zS�]*�k˷:����S���{�_�6��Վ�r������=��=rD%(Z�0���G����Ǳ_�p���3����.�g��''�^]mo����pw��6�����@Q�Vuc
ׯ_Ǒ����&VHso0� �5K����������*~�Ds�H � �1��"ؑ��Uk���y����q}yye�6�����;��/��G�y�g?������pxt��3O>�K?�������o����=^� q��953�,���6o]�8�w���c	4$�?ѨŅ`ug{ms{���"���5,�(S�g:^)E��θ���X[-�<�8g��+ނZ���z�I'(�b�V��(0�Qk����O���<��ß���a��zP���&����NW8�v{Wz�4�����h4�-�ţ� �W/]z��O�>�C�~{m��C����Q8���d�`���G۝]�T��[�q��^�94�x�K�8�	��NB�a�쎳���4��b�%�/Jv�g78�	�?�+���@A�� ������������[�o�lE�7�l�J��� V4�H�
����p4���Zn,�?����[k��p���|s�+#���hyQ�%�-C�b�.����b����¥:�����2/5i�Q$�a�f9P ��^�t%-��Y�A�ifO�[6�|,����a馫�/e'�C��v�Zi����Щ��=�ꗻi��QD�P=��%0+@���`o���N�v���o�˓�c�;[�j�/;ɍ[�n__�v6�8��Z-MN�W���)K4���&�V_v�\+��]�~���&����N����L��xΩB�-�$6���;6�jU��֣��`�L"�(!k$\)��
W��xY����_�� ��Q�붺
��g1k�%��U�va�!c��-��k3
C�i�5D��a�&��*��4�إ���G[pn~�)l�8)�����G����T��J3�A�/��-�w��m�?A�A�@�x�7f��aSӞ������i��$��c>H��_��_��HK��?�9p��x�`��݆�e�DX+�	s��p1��^z	�������	�«H\��`Ϙ�3�<������G^��/~��@�~���C�����M�3�����tuH���'@#�Ӄ>LC[KQ�fg�o��:y�䣧Naп�5�!�՛o^�U��+�*�����Υ���W~��Q���@���
+��/�'N�~��2�O��?���anw�\S��8����R�r����s���4�aOK㺸m}��Gܼvm��O�/���pwK�(~�2�j��}lm51�����S����O��߇:us�>��?��Z�5-�$��߀�-��H�x�ş�ɟ�G?�J<6,o�|P���^�7ku���a�4��	��ԥ>s��=��CǏIR�ү�Y�ʤ�����C�h��[��]�AQ?��?�E����z�w�z���_�/O<�����ak�u>��2�V�@B�R�k[{6C��,	
nl�����^:�ycE��2�V�P���X�K&a�q�C�HHq�����ռ�0�9�\���~`J�[Mހ(��o,~/�h��4�/�/�vj���\W�6��lf�������h�p�x"L��;��+o�[�VZw��hkM������&���o9�G��N�F�)���w�	�!���,�` P.�/�L4��r�u��Jk%p1��a�vw~����`�i�f:8Զ'�U[��[��g�u}�+��ղ�1ǂ�#j�`��I�RWM�j8Mz 0�Q�촪"a���/��'�$A4��N�~,�z�'��J��"�03�������Hw����0��D���
:�S@��� u��>{>��X�[���
�X�L ������Ql=���/�����ƾ�*�&��k7V<;V:h�O\���g�W�є$��(��;�Zckk"G1|@�B�)���j�Hb<�R�^\)V��4�j��Y�F���'%om�?�p�Q������l�ɦ~/��0��'V���ٌwGN?�������n�9=�\*����n{���K86Z�3���e�9���c���]�K�#��:ێ�$=q<�;���=v�;��w|���u�.�}.�֎]z�'���wc�o�����t�����ϟ?�5a"�H�����g��=�裒%T�ڭf��i��%���/.M���v�x�h�/��p�7��|�}�B�\�~��/��>�!�q١G@��§,����%.Di�H��X�<D��Z��ܧ?s���P3S��kŎ/>� V8I��Z,��ο�ǟ�K_����ѽ�@u_ɸl��\�2۬�'�;	.���
y9������~��Q���H���o�����Ͷ��W6VDwQ��{��͘���+���gO��A0�r��@~Wڑ9�Ϝ9�Bl�_F�m��������᲋ڧ���V��詈{�;7.\���`���&��bZ<"��h֡M���{쩧�:n���&[ӒyW.�}�M�1�W��67k��:Wp0}s�V���[��"0��H����*u��ƭ�7nA5u�`ks����~��~H��*�����u�+�f�AG�����ͪ��#NS�R-MM�����ͥ��n޸�ޯi�m�n�#��H�D�/�h}sazַ�R�>�ԓʄh�=�2艂?bʎ��nWhaf��͛�v�{��	����ag C��b�n{sk��MA+����+��3%�}D�H�޴��c�:&pc�9IJ��K ,A�hC����� &~l��j1T\	1�� >��ɡ�e\�2#j6`��&�&g�777��6���$OV�'��.Xi8������;�z�pcU2%/L0�]� ]����N�B66ۖt�v�q���5w�Ӌ�^�V�|�Ր��p�H���&E-]���hP���Bi�"�9��	E��D�R?�>���I}F���%��T��:Q��c�y��/��v��o3/D9���J�F�5'n�P��6�+�=�y��wi?��/bX��d�wY�\���Ԉ{j1����`�ۇHa��"T�P��eQ5S���0eL���gtm)��gu�eY&���EL.E�,�̀j� �j��(��Dr8��� �Ә��p�,��7֤�y��}�O�no�����<�ԳX����Iiֲ�{S�����$�,����"F�T,j��H��4�7���.#�W/]��'>cJ��?<��1�S�<���x{�	?,;n�_��1'��9�����v���������זWVV`�����=��Fh�5���t��:�0S+$'_+��n»�{ �,��vdY+�іT��`�'N����O��ή��K{0�+��>��K����{n���K/����T�?� �a(������|�M��h����?dNP���P�4R
��x��5q
"�wz]�g������)2�?�={����0���ʫ�Bn?~Rze�Q
1�L�����}��}���_|�ŏ�㷷7E0w$����Z.K��������3�h~���#���g&[S�����[o��F�"8�o�>���cG@9P)@N�;�Z"���ϳ�g񬕫�I9 ��*����%J���~��~���<|m���O~˷|��x��������]�J[�8�8�-zY)��c�r���� s��o]��q�&_~���x$H8?�	Z$ _l���I*��G��nE���0k�h�;�"h��S��M�S�&{�o���-HA �5����W'���lw�v��=�L�cSF [�-�iҲg�U���}��~�xt��^�<��!�3kP2�ԧ����
�v� jV�"�mI�*�=��M�h�+�lJ�����#��f���0!WÏ!;i�t��|!Iru�"~�q_�bD��}�T��%g�
M�E�����h�$w7*��R_mD$��r�������5vh���uH�p��\���Ao ��o����ޠ�zs]�4S�Ib��#mA�8,pl���F�`R���w8�J���[�����8l�� Um�9��&�f���=�C��|��/hl�X���0@j��p�6�o��І;�zc��]*v����F�8�.8$~X�"���`'�Ѡ?�U�U�m�7���N�@�Yf�ğ\�	�AH�6���L:���!ޔ8�Z ��ޮ`�k�`"k7n�6��S���;v�����W���v}mb@����l�^/ܼ}me�[��r
˯�lu�^���p+����ݞ��mv�)TH�1�o\�Up����n�\u��eqQc�&8f�����}�''�оh]�J���{�����%L�Q�ԼS�N���NJO'�hHTkլ�!�&W.
:»j�������{�|�X������Woo����?^�r��V�X1��@����	�LO�
�K���0}�}g�9��4
�(�5�9���_9w��z����*�4'���ȲSҺJoss��?�K/|�_{��g��Aw[S[�Z�ȡ���lA{�y�{�����dXx.�s�._�Ζt��o�.���`���}+�dukKj��q#�[���q�V���ys�}m�ʭ���p4�p���&iV��K�d�|���*Lr��Bq�1�O��ڡ�\XR؀4UsB^�0*��a;`���������o�8���t2twnw�������_<���"�O��>��3�	&܁Ա}j�W�a7o�h���;7��`��ܑ�-῅��*��c�W���XjD�ʹ3W��_�<a�0������Օ���,µ�[�鷼�[����	D�iM]d�����M��7n�@���v�\[�jK�M�����p�ڍ��t��d�Q���#�w�����0��bg�~wk�;ؾ��f�&ck���'�?�3#��K~�^ߺ�Cq����n`�?si{��ܣ�GPt��VgvǏ��q������V�����vSR�Ұ;�U�t)����qWR��D�v(���^?���V/k�������eq��{8Ђ?�%�Y��(f~�u��#G��f�`_v�Hv�0؎F�tp�������w��E�^W._k6&g�w:C�y�&ⵕ�O(x���Ǳ���h�t���fHǀ$vm�B�\��$҆/��xq���W;�pc�|�`�&���ڔ6j��$�hDh�Ų4_la��� ����(��x%�w�cY]�E���鯔K�kW/�7����*
������U����ԡ��ӿj}_�W�p8R�b�(K����G�HT[U�Z��)*y�Z����A](��3�)%��y��Dku��o���r1������fR�:����ˢ}+~�dK2�JE�A]O��bU���n�}���_Ը���j^3�D�J�󡧽8M �7���>��ߞ�����t���A,Q�-����-�������d�̇أ1$O��

�i�[V�b��b,�`���ĖH��zmM�:˜G��0��Ec��{0$"k>���vZ$�|�b�u���%���ϫ7�Z��)��F� �j�Q�a���&$Yכh�	������)�+�Gi���,YQ�U YWVj�$}�<	�� �JNꅉ`�,>���No��~���&;Ea5 ɮ]����3��<�q\7l�w�)�������5ɒ�]�I��q�8	�[A���lBW$��zGv)*�� P�R���!�=��`����_�݅e�/����v�?�-z�X,�u��D��^A�ժ��z��ǿ�Y�H0�/~�̌�xQY�5̈��Ғt�l��M,2X�㋖�b��--�cL	�R��h}9�E֬,�_�}sM9l�6����6�X;2��	�xC"�I�yQ���eI>�?<�;�+�	��.��\]�v;3RSSqd1�~`e]9 �H�p�����u&��V<��T�1T�GC��o����)�v�:j�jD��C,{�:�q�ՍB���RuŌ9��U/�P+K�,�M���k��ϱ@�Py���W�V�ĕ�`lS�İ�h����AB�r�����,�_�Է2J�蠶e�����_�bz�P�SK���*p�CM6q�,�ӳm��/x�d�5W�"�q�ֺ�rI�|� Aؑ+
odg}`�������*��;{G({S�`��	/���3(j�����%:��o�q�w�ԼCVe�F[T�M	��+�u��1������k뫫�o=���s�3�>@C�q��f&)�._�XY�9�j��M�mHW�M��ͥ��)@�fvaj̠��vz)c����� R��SV�f.>_\e�����Iܛe�RJ>�>3?SmT�X'f'�q�Z�0M���mI�P���;Q��&f`V$)߾;s����k�f*���C�c�y�ɘ���QRl	��Ai	��UsD��W��IW)0��� �/y��/B/�j�1���k�d���$A�4]�v����^OL5�gIv�;��;��/�Xk���ðߚn�+�䲭o�ѣ�>~�Б�.b�;�݋�/m��'Ղ@<�b�������
�1��ܢ	AͭdD	?��ܟ�z
3�
`?6����_}��J��x�1��(YA��W�
Ug�l�N��.����<��R�zS@�����4eVƹ֕BG��ӧOOO-<���W._��o6'XϦ��̓����!(��j(o�HL�d#I����h��K�x�T�a&5�A�f�tY�%�j�r�v�-`�K�=�m7
'�ba����;�}�
Iyz6�
%|A��C�gk�����t����rwk�*�"����X2*I�����O4Zӳb�UZ(a�K_[��$�؈���u���I}�,����Bɢ_z�)�y��}��2��K7c�n
Oy���v"ϗ=ǭ�Rq⾓�v�W�^u�©S�jE0�%eN��Y��K��"�ۉ�7������*�v@�K�J}��ԣ<�������I�V�CEI�u��k�%�����=-,ȵN�Ke<��T���RߨN,������ȃ|a��οN.�ꪏ��� �$�b�x(�փ�TY���y���Rw1a�WPuñ��N���;k�A="��͡(�I�`�}~OE�$��{@���YpaP�`�%���R0"��N �	�xfҦ����_f^yU��ʄՅ���-���(��'Np�y���eD���n�`�G*ѭ[�خ���лYXO�������_���N�nr�hn�=5�D�	3~���Y���99~���ԈO�I��q���x�ѯ���x�6_۩fD�u����S�������}������
��d���,�2�GcF�GB�Ka�C�����Ӽ˻\cNp��);]�oc#���t��m�jX^E�|��͆��mmm��M�G��|IDu_�� �4���u|���KB���R@��+ɑXY���yrI�n4=$`K�K�ڣ%�Y�Eh�9��V����9'ˎu&��VH)�E(Tjm�w��tbia��z��_���_z�%ےz���i���'[\��̂{DO��6H�&F�YS�a�%��1�9R"|�
%�T���${w��X��	&r�A�J?���q���� ��VWd:_ � d��|�̙��/`g�u|r8>|x� ����il��Ţ���h���@�}�E����6�9~����z��$Ю���=�yo�&9|�Ph9V�@��y�[�(�d�� �(֪X^MZ$��N����������\�����f�6��{Ew�R��'q����������(������N_�r�:�Ur�?�j��(��&��q!hK;.MJr�?E=��aYmevBOH��a��5i&�N�0P7�|���7Lf�J��xPann��Bbx1��T��,Or�7�G.Y�`�R[#�+����J�p��j��z��5tk@�Π?GǕV>s���95v���bk9���D�Eqڒ�QW��۔����&4__cH���i� ���ݝ����d��vv�_���$�Xp=��Qtli�=�hzz�X,9j'�Oss�����V���˗.]b�[���@;�\,�$w�3�G��A�0a��&�:Z!L���
I��¡4S��3�QA�Cf׵�4�������\����@��xb8��K �n(J�7�|3��`jn>ǷV�_!&<m_��Q�/K��Z��"����q�]����\qY�]P�B�Y5[���v�苚2o�Jx�X��^}���G�Jq��lnކ����̲�hA��b���Ą�#M��c5�,_�|���'� ��,_�>�Kً�i�J���a����V��hZ��2I���CC��[����P���\���c�<z�ƭ���D���avXjG�~b	W����i��%��@0t*�MCucl��x��:=l�ڝY8�0�ӇA���戽�	�#��%]ҥ˻ot�,Ͷ��q�oJ>��ƕ�8q�ǂ�KՈ�4㱣M����BJLg��|�����=�j; 	Ƒ��N���kS��э�8B�vD�:�9�l7�U!fW�Á� .�E=ޔ|�񍕹B���'%��*����z�j ���r�懁L�s=�a�J���i*�ACº�|"1
%5|�)�:a%@65�`��x[;���F�	���v6qS^\v���9�:Q҃Ѯ���D�졪�G�z�����Ξ=�� �Ž�4�k<Yl,-j�Y``1�_�òq��f��=[1?_ҹ�잝E�'ذ��]O��dv66oNs��&��b4՛e?��۷o�n1�~��?��7󱳜m+�%��o���D��qO_Y�(��Q~��H5�S#�yUqV�i�5z+/����=f��)���j�ֆV��[�����>����u�>��� ~ƙ���yP���*z,�-'
�$��f��d@�]�+�ȓl:���l���$F�)Im�
�Ej�-���V��[�L^�Ų���n�N	���A;Ɗ�kT�|��)A��p�l)z�٨��!ga|��F4��jf����9��M̅���1�(v Υ;���`�'N�>���1����6���+�"v��v$i�{�!hŢ�P��)�^�٤r@�>ΐ5��,�0xJ�����.&ص�v6m;��3(�i����КR�3:���fi�(�6�!`Oª�D|��_|�0��[oa�l���#��T�[�bkJ� ���u�OnK�E�ʤf����,/�%ŘGN���R��ó��L�
U/�"��A��v@�bk��1f��zT�X��ַ������*�X��3�PǢ�a�%=S���ŎکR2��$��.��Rpj��H��X�����&��(&��+xа�!�A(�_2�sJ;^r���Cj������٢3-&����`�C#���
0���S�СÏ?�x��A	��A����O�0��`}r�Rr4��i2G,30����'�Ǆ��\�z��9����u��MS��p������GY� ����Џ_-���'��Go����������"��.���@A��3b��8��{"����)��;�&qb��K�&y�U$Uf��RDۀ��=b#XX��g���T����z��нo��j�M�%�M<?�))��ʃ(Ӣ��N��7���Q٬:�[�ꫯ��}/�tg`d�@u'��vV�7��15��w /A��P���[4,>P�t��z���R!xjF��F�(dR���X'ג��\�P
�����32��cS6��B���4���U|���S�t���iS15�����ر��tu������'�
[ʛ������	ܜµZ��z���B&%"��3b ��K,vmm��J�qA!���$�|�059�զ�����T�7'j�%�͕[o~!�E���Oq�$�mm�UU��)�w�cg����5���$y]��Q�W}�{+�;ik�ɒ�~�N�(�	ܐ����*��[t���u�q�,� �-8��0�>S4����x��^+�a�5�	�r�h�
5�~s�V�ߝ����ޚ��^���[��f��{}H���*�����[�$Y���Q���mT7j�x��������^��(jN������t��#����WN����3��[`�mD���GN����*��;;mh���O��25��ƩɕҼ#�˝����z��	�Zֶؖ���1��Pа�%�J��%r�8�� ` �I	N�"��:B��h����榛'��぀�Fc���'����ѣ�� N\'ѳ����Z�ґ�`�%I��J�Dqѫ	j�'�e��Xώd=mq��:Z����iN���v��ĴK�N8�v�U@��=/� �*%u�0�]gO��2���l�]Q���H��`ѻie�C!`�OC���Փ��/�b����[�{>8�����S��-ĉ�VR����v�ڵk�zC@�Je���`����ȩ�f9ZWkD��ӭ��7��s	��QU2�NH�*��tX�J:^��q�����'7�g���5>(���l@�CRvo!�g�����ېa��,�|ҕ�R���.��V���j�)k}k3Q��D;��k������q���E��y�����ej��_��vw��UM��"2DJvC����X]0/�ミ4��I�/T��/��:�U�/_�|���V��OMMz��޸3>��M��q������䥾1��͗�Q��4'�Gv��g?�]w��ZE�X��"6PP��5� �f���:<pO���TWW�M.��*����r�I��r����	�\���6T�~
��2����ߠ�m�a��aWr�!�{R�'~���y��3��V��T��ˌ�r��������jH�]�_kM>��c�����+o��&�{>�h�3lDA�\��\����^������{Nf�e�x�����t���_�v�s��1�s�Y�{�0���~��ٳx�L�����E�#i0X���z{��i��?R���z
BW'ƾ���Mm�i�t�p��i���fk-�^w@S���~q��������!���$��>�MA�0㰕̖'�൉����+&��G�5��y:�+��O��fS�J���A�@�R�jNh�$uҏ�RM�.kb�t'ۓVR���`i;J�[8<�a��S��{XgL��F$��)bތ�� �vYr:;;�
�)�/_~��@�l˺����|~�X�h���$�W;��H;�tG{Z�Fl�[))��6(J?ê�W���������&1Ѵ��QF��x7å�~1R�q�8�6�R�cj'y�WGǣߍBq���b00�/�������N�Ps�3"k�DiW���Q����C��*ƱJ�����7T�L�^���0����ՠ�pv�c��+g~���"����Ϥ��׃�7�F�իW�����j��u��C�8�35���Lhvb.h .(L�� �����e_��.O/4�no�J"h����տ��t[Ⴝ����������'8�ۃ������t�9�3h���e!��Z�J����
����17���7�rL��ɓ'A��5�?Ym���C�x��J�ݘ$ũ�J�z�Ȓ���P�.]~�/?����90x�P*�a�, ���_Q�	*�N/6�?��,�,����$���N���vjk%�{=��Op0�<�/(�9/�S��n�t�2f�7W�'9�2$���lc1�������W�{�!^��#�1[oN�3�R���W�p�t�덚-�ӠP��B�Z+����n��' l�p�r�
]��m=w��+OJ� d�����������N�$E�G����ss����_,---Iv��Zգb���ъ���y�?�;�����b4���c��j���dO��mB9��~�x��x��/}���C�o�T�+�11�ʐ?��;��,��b��֖�4NM���� �$��5�a����6Q�ݭw}��,��\�y�Gq���RìL}ܸ���Ov���fsǎ/�p1%�z6��nK�����J�.�r�\�0m�^�R/�<����+0_S�c0����P�Ȑ�޸3���QP��|������Gg�g�����"�\���>&8�Ɖ��q���cG+�g���!�[庫p���Iu�ݽz�jk^�B�;�43]�:R��Ƒ���W����T�v��"����%}+�t�6ݱc�Š�h�RXp-w/��H_���O�O�X�dIU�$鹶]���"���	�g-������AP��t��D�)���Q?�\�L�#b��:2B?(h��!]g~v�v�����'?�5qq�fK�foM`�ö�=�Z�Hї���q���O���&�8T=�8W�,WD>sn�8��e;^�^�#Wo%A.�_$�J���Gϋe������S&~�c�%wD��,�)�_Ņ�����*A�Kt��>�sސ�ɖ2	��7�}�Ϭ�v{������&�g`�aG�ƣn���ǔ�C�_�����=��DD372:]F�������H^��Vv���C��\0���U��J�y%�ee�)���~���Ϳ�7Ǐ�4��~�ఔ��J�k��F�j*4�\�h��d0���?~�r��4@��i��HX!-�Iʏ$���вQ��fz��GT�5��%V��+W�$��S.���`�#7�J�aH[�ơ���v���@��� �[���aF��J#���g�l�I)�T�p}}��W_�%J[�na�W^�Q7kgM��q�D7rd�E_<��"u���D�t�β^Ԁ'������V��Ab] ���:7�� 5�S�M0q|����)���5W7BU�B!Z����V�Zΐ1X���$��=ƺAV�0���9�s��G�6s�A,�?�E_%V�U�%X)(-ǼE�U�'D��s.)�z�/�R�0���[��L��4~Q���X�\.p^`�����1��#� �Hi�I�#;u����}Ko�H����8��H;��(�=5Z��/��и��t�;�+-A/Q������g�����$�ߺכ���gét/ҥ��7[�,M�R�&g��Mb�����Y����=�xZ�D�q�@����t?�\�0�,n����wrX��*#0@����|T'^�?�B�&2ZDN�|mQ�od��UΓ��q�nS��}񪩾6��ih�z�0�87� iK��T��ov4�EPը�F$@KV�c�&8 N���bE�A�^��Z���ѣ�S*�B����H6M�4	F
�+��yIQ4�f����2_�٢D����?%;U}�[��k�X����D�G?�_萀����F�N��zn��`3y�L������Xzd)�/�h������7��� �P�[��N����d9ML��č�ו�蜓|�$� g�e���[��{��_>~|Q��w�����;/H�$C.��ᓐ[mq�Z
��:W �[G��tz��>���K��J��R^��Gi��?�*V�=W��\a�rv�7do��̹K�`<���`�V*^����gr��|�ʮ�u.��o�1-�4�0*��B0�?cKG�ӧ%�>�[���оe&͹�L8��B�|�	o9��o�5me~f8P�[�E��9z���#>�js
�H.�̔�$)C�������by@WZ,׍o�<:�y�����1_z.DY�xVI�E7Il�'+sY��
I�� ѽ�d��ۘWrߵ��� U�L�߱;f��k��j��k�n�=�T��:����T��w2GL���|�1VZ���aAl bW�CBzdD�/���N3���#=�F> u������Jx����(��HD����2��C�<>V��k�u����jc�n��E*��@�r��_��EC׳�U��l����������1i�4%U�3����4y^��h�*��~[�R�&��`-��z1�VO�N|*�)Xj8��*��8���j�g_��q��#K ��\���_߰R��,i,�4k���6���R�U@VV��ԏ5_,�KB���;��ݢfM-L���K��cv���;
�ni9e�(ʒ����>r�^W���>vb89�1Gt���o!SK�T���*z)�(*��a�/�5'�ص�mA�i%qB�ȸ[ͯ�f�����}a���"�q��ĤY)&T��$�aq�aɎ3�aj�P+KK2[_�*��6����z{L�4��r��}�c����O�8��B���u�r�l���%ޙh�b�֤������|�M��q���Ih�-�x�gΜ�t����L�᜷�%1p}��K��Z��u`�6�*���:�_0�](
1������ۋGI%�j`���x��k&]�0,���2�îF��4���N�'>�	�P��W���ND)���kȌ�����X�G�hL�-��x`>�������h0LY�de����:�X�3a_�k�?����
��n'�.g5�M�	Q��^�xߑ#�����2c{�8K�4����S�vI�?S�I�>V)8jXk�gL	$�655��������x���O<�T8�*Tհ���qI�N��h�3�?�+���Xxb��稸�ÞZ�F�4���VZ�L�]u�(ϊ����L�k��~�� I߉_b�Q�P�ײ�& �k��c��Q?�/�qvū���ڀ���?�0��ٳg�<�'''���Ky
dQ���^��a�3�d,2��xT.�z�%ie�|1T��U<M���1rr����a����Rkw��-[�nb��j�R�و�k��KC�Q7�5SXL����)7�/2ќ����R�R�Z?�4m!(��֦�%r�%�C�p�{��VY9��lyb����:�F��A��d;ӵ��k���"�S��8�Ç_�p��%�A����\�T6�V�T3)��2}�N�շL%d�m���-�ͩ6�H�e�ْ�"�׉�U+ZQ�P.%�?����t�w�p�6e�ܩr�(��X1T�h��F�=���-���NNN�L�be��u��w:�J�ζ!,�����CH̜�>��])�Mbr*�ʒ<Q��w5����j��v�wtJf�A��=���ׯ�D'��
������`g�\.�����_����g�pA���_ҹ+0/%#�HETX��>�غI�b�h�ӹ[�(�[ۻЪ����0Ȉ0hB3�j${�A�d�a ��	�V��\n��?U�e�J�ZM������o�����N�"li�g֐���:�W�9�Ь%��`��Y*]#�gh�~��`�q(O��Z-�閌��ֶeX|�hn�)�Jr�Pb���@8Vʌ��Iq��V�vfff؃�N4�];Č�N���gN�{��Wp�g�y�s����dK�4��V|
Kӂ`�e�j�'[��f(F(� >A��%�E�J����1]����������ΐɸk"�Z�1������f�w�����Zl�0#O"�	���%���-0;�^�9���ӗF�T׷Sd�w�j
$nFc�R��?v��l��t����ϭ�덉&d���\Q�o�*��>�v���j���҂)c'�g6M]�r��N���n�LC�pK���۝")҉PK�J���
����wg=p}#K�򘇊��$IzK6��|RA4�P��t[n"eu�K��6ٜQ��\����,�\m��~>�M`���N�������-E��F<e	tI� ��"x���Up�etx�,�E��V�:
{J}�)	��9~w����ٝ&�5� f;�e�}���c�VN�0kE�@N��(����aS�mj��9WvVC���U&�+`�2��,5�s�e�d�oXFڅČ#��t���������)H��G[m}�z��AY�Hq4�Ĉ�hIQ{44�@��O��0ȳ(��$Y��?��y�S`d*�In޺�+��+a,�z[mqx.���Ґ�Ҏ��x�8q¬���J�u%��e���2`i� �$�-F�l�SKb��vw�\P&��Y���.��7�ZƯ�d!6-�+3��4�U(���������H��j��`�����,6l.�3�9x�t���+LU�b5l��h1��:GOB�B����a��#�;��ց�ŨfG��'�:�
;m10
4����[o<�]�l����Smc��v��kb�$�;����<��!,!�/��8*�-�¨̣� c:�(adS��X�ns�œ��#״5�ʩ��h�Q$���0������N�� {����^Z���w5����'�;8��x��FbV�U��0�077w��U��?h��ކ&��"�q.i��H��;�k◘����y���e�@m��Bh�T����1���+����5T��J��dN�DA��(@�վ��Z�����y�������5��E���!�2
��|�qXQ^�����1�����2�d}}�R�d���L-�g\�uD����F���B�gͺ�([�4tDD����j�d�ҷ���Nzz��U�����,�+i�\ ���X���)�tz�Vs�L9Qz�=�f�<���4�B2��ĀLVFj�mS�s�d�q����E�ݨ	�Y�L���+P"#a|��������e����5={�b���~��pe�YemP�]�,�'՟P.U��l��[�}�qgkg�UI��H;gQ� ���۷�\[	yf�G�S%vнND�����f�1i�ǡ$}CÑ��Hv�&��+�هi����-3聼�%�h&�>��tAL�f��K�0���8$H_���KX���b�u׏Mh�C�Y O������X]]�]\����Urd���'�'��$C`7nݴ�ZAff`������LHS���p��u�����ٚhٙv��kc��*�$֋-Iì��>��Є~I��D�JEp�r�Y*6��ݷN_���kQ���B[ "�;X���o���?v��g�yff�%�q�(�%�p7-͟��=TiV]����ci黊(5�P7X-Z�Q0%-q�T
���g���'Q��S���$�1�&9�t�U����~�P`�9���h#���Q%K��	<_�tL���nѱ��K���*P|�R!�<w8�5�����J�m�}�⅋W.OM�DMM(�Q)9�����o�1N��Z ΐ�z�g�h,\b�?ñ���s��lϬC��?i n��_�~sq�*���P�k{�Ȧ�~����d�;я�, /]�+r?k�d��n�p������aϽ~��D�<��jYc6`bOz�&j���=:!��[��g	�����$Oaඉ��BZ�p�0��	.8���n�՝�3��q\2����H����Z-�Ƭ1�(�Y��m�?�je�Zl5Oܒ��8�.;��S�&+�Kae�B�E�f�(�Z���%a�֞ˑq�+<������!U:��,AL�GL�К@��B}Oy�=����\4���h�p|��F�QD�
�2�ZQ�1 e�x�n��Tv�M��c���g�q����h���\ć�]_&�aI.�ġX�`k�_-��Ϛ��	X����34;�"hc��mtz�MF�lA���
p�e�b����^n����4΢7�s==�pd�?l;�GĹ+��-.��ɩ��%�PR���L�X/sR�,X��B�J�Z�,�;�R'��S�v6�/_�p႐w V��ж#Zȷ���8q���Vx����%>���$������v��N�X�XL�T��R��t8���4�X��I�dT��Sf��Qu��wct�����7��=���ǚ�o����E�C���do�xB͆qD$f)|8zT:�ܼ��u�K5�f�l�2�����#��b9{aA~���H:)���5���H}!���C�I�֭-:��:�bv���Huw]�oX�o8%Wv��i<���t��`g�xip��_)kIF��j���玣p0z�
��=���q�Q"�c1DN�V�6�#М�V� �͎�H�� )���CO�ܱі�V�*9�z��:j��N�ؑ6�QΝh'�D�\n�D�p�`��ʑ%�$�^R	���ԁ��+MO�u:]��*���ǑT����-9�@Rc��ד����I��P��GC(���(D��������/��.�Z�}f�������f+�it!�?i�[������i�Hn���+�A�r�]e�ҷ�Xp��W��\�PJ3��㊝��^Z�c[Q"�u�\���l%�>�7o��J{�3ǉL �p�Эոbs����ߨhƺ[n��������a'X]�Q��O�~�^e�"jb����}���^��B����.<���U��'��&?5��))��Y6k8;�`/[;�8�Z��H�
� Lg&G�J	D.µ^�,}�]h�&F�x0�W땡�Ē%j��N�\[]Yu�Z�V\*���ӡ��O;�+	<|��AG�u����bG�fc	j���Y-�9Fä=ر���p�,��Jw9��K�t!������u-���jy00�-���+�@`���D$\��Ag4�T͈��Xg�A&�ʃѸ��R���xLXh �_�we�=��V��/̔��N+�8?��U����C��A��zI	����s54@�aa�U������_�3Lۘ5i���ތ�|�Ù�+�F+r�7Z�'T�8�d��aľ�%'�d�[�K%^�	I$N�hA\beBZ<��:��͈ā�S��l�41qxbb~i	��E/���A:�� �G-�!Z*$ͺ�v�r�V��M6�,�ĉj�סM���&hW
U	n�2y�������vc}c9th~jjF�a��XA�I�b��."�V��ʫ�\���N��V�b2�bh�l��>�tV���2V\�-7>p�&:�ŶS,���7����ُ������5/1�&�4����/�e|���*���齾XiuEc5�y���f!�"��ٽ���C�\ϷR߳�����m�14��T��*��5q�5Y��
��E����I��a��ݥ/D��$/hӊ�;�n�:�~k�K�W�:I�\v��:K����u�á�m��W�B����b1^o߾}��!�qL��'�{C���L�X3N�z{�PY�x`0�@�!�ScK��f:��tHZe
��)��b�1�Ui`!"U�f��=!���8Y�P1�-W𯈨�T�Z�-�J����9�Y����"�Ұ,ɝZ�u��c�g�g�D��g�;�\�H�����T���c�=��tf@�c�{��`8:��6oнy@oˏ��&
����寻��a��&��$ɚt�y�/��^i�/4�i[�dZC���A�C���+a��w���X{Y�8���8���c���:{}�_!�} `)G�az�`wx��o��!Q-yE@9�.����(�~ �`F��q���f�#E���"��t�ڵK��q.�ff|M��*H�7���_�0Ɔ�|?Ʌ��\ew{ľ������q�2�T�hI�d���ރǛ�;������y0͓,��*�\�!�<�TI�d��[��G"�9�e��ך�7�MD�^�PI��>�����i�3��搸�b-�Z�t��1�lgH�\����͑#��r��y��� �̾��A\������	[�l�.�����.�L�h��ʓM�}ˆl̇�{��7�"O�V�0��C�������H�F��q�R���v�[�d����f�:�[(��e��eCV.>E�]��߁�ʋ2�rΈO[3����<lᦖ��7N8f��5U�5E%S@'�P���Z�+�p�כ�,��r�^&MPw���L0.���7�Ĝt�&�ʈ���z��4�-�E���F
�!��K��%�j]�i������0�3�1��(+lq�BJ�K�C�������� �;�NNP�8í2{f��	Jy�3�+���z��Vf˚u0fƝ�f��m�Ə�81�����{6�h#�ٝW�����8���t}�
$�����lI����*�qש�9r+���w���1#S�B����<�v�0��p6��v�GD�,㕫��X��J'�0-�&��<��"(�,�كG�����Fx��͛7�7��	��߰R�ޯe[��[�U��0[��j���8C�d�^��<� �ǝ�J�i8�^�x&S���Ȃq��{T�O�1Cʫ�d�����x�R���������677WVV5�A��k�:X.+����U���B`Wz2�,L?*��e�Q�K��\���:NRyc�7��*o�E��r�#��r���%[Bp{�� ��@��4zJ#�AHJ�`*�����������ʴ��I��Hs�k�m&n���|�k{*1��8iԬ7��f�\�[�d�8+�s[�c���o�����(�L4:�fԒ�K����(��+�H�����b�{=�Е�� �2AȈ�Qe��
}u&���� F\�,q��*����$��je�������� ����Ix���7��f���Vj��T.!�ÐbL'R�+��γw�L����u���uw�?�0���4��zC��O��5#Cl�J��t^qn�^~���%��3Ҽ�Ď�c�.�͗V������7��OGxO�F��+I}�~���i5Pbk��ռ�ߌ��Ѫ}'���A�;%�բh�՚�̊ȟ>yṒF�p�|=�n���k(ַ��|�~��\YY�s5cq�L?�a|Q)�'�C��0HDX��=����?���d���x�uxcO���
�ce4�,OP�����	]3����iվy'β@���H��%������իW+�2sŢ$���yJzP0��g��nloNLԦ���B���6�3o���8-����>sL�g;�ڨX�E�'���D]&���v�c�X7o�\�u�ikD��S�Xa�0/�|�X�dERڕ�S��ុ��i))ݕ�R���o�� I,�<�$駒�T���l^���=��FyeA�ۗ�X��7HF�gJo8��(��]����A�v��r�S��?/V��X"KM�5���������eqF���2M�u#[�3�����e����E��&5&;������ᰄJ5T���scL��A]���ixa�k،�!>,fˡ@�ie�}��\���9����
�I^�e��<�]5Z������้�"��׌���gɖE�F�.`nA2�KZ�(��gu����@{���@���K�o�Zi����?��׳�k��{�J���uܡ�)%�+���C�cHO�]�<|�̳cn(�G]'�������Q��!�N���mo��� ��ʿH�&;s:ĭϝ�{���+� �81g;=v�w���C�f=�<c��FINh�t=�-����]�j��8mΤ1,;�-������{����Y5�j]R��z}�dU���wbǾ���.��a�2[vv�ܹsV�%,�7�-�����&��U����]X��>���?r�'Fv�/~JM�;���慽�9���t��G?z��e(��$DD��|���԰8K��<~�8^�B�R�ϐU^;1�����r"$�\�����$��q��>&�:�B�{Z��9 e���ä�~��8��-�.��"40����e�p�T��Ӕ�s
y�*���o〲���m��<�ه�z�"x��1���nӦioo#!� ��<M��`̾��V�Sbg��O"��N����*����.k�C��I���L���F�e���3[�2	�����<Q�Mb��'��^+'��x��fem��Sf��m`v*�_wJ����IZ�n�z;��9Ym�i���8Yjwv1��I�=m�O}��/��W�s�����;?/k՚h�Q�Ȇa�S���J��Pk/|�{�R��o�M{IXFus�������le���C�a�g�s��ݞ�O� �Rה�5c9���)�������Uo����X���X333ν{n������q�ؑ/�!�]M�e�T��3u�;�U*L�L>��<x�W9b�3*�w=��{����@h�PR�]�o\�.xw�`7�/�+T4b. �ޜ��`����D6V�Q}衇��-�񳁞�M�:j(���F��2x2���֎��Ir����`��K�~�~ǲ����k��z�8�tU��lJ�(źرsS|O��dv�<��f��y�Mv������>-v_��<&�d��y$�آl��x�=���b��"%���L6��s��9��0怶�W��x�:M����N�$G�<��Tl�Ѣ2�V�!��IЦگmUG���� �9����i�[�4�h��Z�����k��ono!C3T�=6�����1�L�[���jQx�)[߼��J��P�Y?���&��!�,={���i�E���ܤ��=@EjGhr�%�"d����+���ņ� �����#�}jH�e����A)�&[l�\�:��b��Sg�@Vr٥��U��W�[����i:�Sr.����-<L"�Eo�����s�va`�%�c�ɪ.��{nMƦ�w谮��9#J<�,�����fc��ע�{F�\9?wHǪv'n'V�.�Ӻ�ؤ����!�_$e��P�����O;P	[_Ț�L�1�֎��F��xC^ �D����*M�Gۍ�[���5��\�qgN>� d[�5?T��.G�1�k��N�[�(���9���od�"x�����߼y��`��"��0�?�X�4A������[Y��}pJޣ��=�гRs���"�� n��{*Q��U�<lW ���� �	ȽF�� t1�dh�y�DG�@W���Ԩ�~gvCV_+�s�B� ���������%�r(�֞>k����!-���WWWX⛪�KY)�ϱޚ��BO��8�,oG�1��P̗���`�� -4�yH����_~�%��� -�ܾͯ}��?&VbLLlb@I�
&�%�Mb�Z�z�*��0 {s���g`Lg�AtW2�}s=���&f{{�dޓ'O`��Z-e!õ��F��N���o��@��x�+����0��eD�K"��T@3s_a8�<�)+����0����2�W����"R��I���IX4�(���sO3��<�hִۆSս�k�i'D>t�^9��i��؝.M��$N$#�qE�s 4nCW]����x`䎁�h�<���_G�����������Z�����4�@WA��e�#Ͻz�{N���{�}����|�L
bF�c�~6�Cy2"��~��G���;�7�y�Fd��}L~��EӤ��"e���y�,}��(ɿ^o��x��d�?~���Ww���k�!1 �ݸ���w�������lݑ���V7��k]���͉Y���c?E��{߫\5�[T�1��m�y�j��l�a��C�h,�ZO:��o��/4���q��Df��尋�V8_hu��$���&��V�t��e����?��g��VWW�pS8�/��:���>����zx�;H� ���՞�ZRǍ&�q��(�� ���.5w�q��t�\S�Z��y���=z�6��8E������|��K���{[��[�:�\۾��͍h"��] +���މK���ҙ/�[@gd��7Vq�P��时������BHa��d��<��Rt2ù��޹s�����\�3�ZQ:T���tn�4�o �<D�D�A�Ӌ��5k�~�E8����w&d�*�'���JʂG4>n��N���壉֯������7D����wJo������֭[����t=)����x�-�����q����K/�D_��S�T�/��K�,���~������H��#�
�ٷ�ܸq��ݻ�"I�l������8�)����C!�d�s<Sz_!��ؔ0��;��#��Ό��ǵ�+g���pv7I����~�;!���ʦp^<UR]J^�8U���A��N�����mM��K�5�J�j8}�����ÐEЁ(�+�ݎ��W"v�t���~�駀q�S�'��PV��X�8n�d��d������Ñ�3���Lp��$���������@�cZ��r��F�����GW��C��R ��k��̺�#�pc�p����Ǎ>jr�Q���h�Qߝ�������/��կ�]t(]9�/�:	�Y�.��� i��:hh�=8���tmu�w�G������������\�Yw!������ߺu�Ν�R� �呮��z�|�B��Ϩ��#�Wp;�e�^��j��q�
��`8$�9ұ -�*���:�8��铿�k��kr6���a��п��z��\��$���Rݯ֪�A��\mT�`2�L���	����"B��uLg�!�ӳˮ��/Jj�5~S��F"D��?�+]���M8i�8���?��m����o�yhD�
-�7�-\��hɏp3&�Fh�>��Z�UkI�B����{���w�}������P���s8߸�t�c�0�`�(���*n��T�1��`D 棓^��ݎ#+�1��!˨���N��H�mI8,�ԭ)�5��=��}��;b<�΀Q�h���%G�C_�3��WN�ϫg��FX\$��g�>�@�W�@8�6v*ca���6"r�6Y����0�M4��]ҵ�!6Q�l1��ܔU�!e�����#k��T� ���k�z����Yj���19�5Aih�8��;[��ظ�lX����4���5j�KR��pl��u�VV����?����?@�v	n�͛7o2e8 ���o��j
=3emGڒL��M|7���W���xa�������oiM���"}(� ���q��s+xz~�8U؄�U���*X�G��.e�×�l���}�W$��Z%��Q��z���}c{{{w�ktv:���讜ԟ[�e6�#�4Q!O6N��ٳ����*�N[��]@�L�B���3q6��<�h�	CQ���QEܪRp�n� ��K�|��ƌ�{��ع�������7�;\%��dUOk�g$�������5�l�8����@�։��`KGr�6�=:��
��N{<�;	�t��'+Z�p���a1�M�Y��f�)�����5?T��������駟^y����qn�[�qސ[-:����Jݫ�Өpq|��\��Q�PMDR�U�\�w��|����"X���V���%e}}}kk�����;��EU&����Ʋ�V��\�u�P�4�?Է�)�?E�a^��(O{��뤍GЙ$�N�������V� ��"��i+�P��CR�^��*��A��D�qs�A�j�_���h�ۣ��Ⱥ����Կ(�(i�H� H}�D9|� N#֖hVy��}4��&1�߽��̉�����GIS⬭��8O>䔩m^��/��������_.u��HtI2���z���+��c�o�.	�+P���w!�v"]&�,Bjp�B{^�y���;��/y���ߺuK�'�  ۢ�d<�(�N��T$�a�U���#&��,={�looyCQ�~}=N���/�p�I�p��1��a
W�(��T+���Ηo����3�՝a�!�ń����	��U��F��^�~���O?�}ʪKQ)��&�܌�U8�.)�um9�j�y�#����*��G+�2���P��Pi��yi�R��Xa�c+������!(4�=[��%D�0M�P)����-u�'7�N ��:]߇��͛~��7I"��h,7z�1|6���j�67�SØ�Z.x��j��L2���T��y�E"f�XKvp��A[ð��x๼�v^��O�ioO7}V��	VX����2<%�d�?�����
�>��{4���	�V�'Y�&~��egAN�nmm�.���%����}���@����+�h���u���-�	����oĘ�L���C;����)2
-o{^��	��鿅S�����GY(%�����Y�R�B����J�Y��	{:���Iw�Ǜ�'K���s�|DӉ�"2F���;��2.2O�&T����7��� l���k���B�?��:�.I.<rm�q��a8v�jX���ќ�ل��L"_����]��+qnnn���A��q��穫��	fذa�X�g;�
6Ih���8�'��e|�	�Q�gJ!��G��
ZG����H#:���"��uv�z5�#V�\Bփb
 �d��Ъ�ekW(���=.S֕�����k�y��@����[o��l6�`9�Rw�h�۸0dd��~z�[r���E�%;�k=�~�,)5�+���vWS�ޘf�J+��^�����0��3���p�^��;�_VE�v��PY�����+�0h�"�A����)�ĥ�Ҟ��[��:��5W���E�"ǁ37"Jz��������820�R6��N�&�*�u�P.�9aN�H����5&F7	fI����*��D���Ф)�h��.�g;U,�U���\�CT���G���ڬ1e��<�ʜ?�_�	��Љ�K26�Tݏ2���O�#��d�=k E6}j�fo���,^���G�A*b���w�_��"|���ȴL,K�����;,�醙�#�v,��TCPZ���s�z�'+"�˯Ȩ� ov��>^3�^}T����pe0���l4\�kw:��j~����^��/��d����p��=>�j��݉��j�����z����ŭ�tt�������Ke<_<ҨU�l!��!8�מ��Ⱦ�㭽��n�:���P�VJ�FSf4��g�����E�Ȉ%u��eQ�L<=%�দ �&�3�kf���rK:�NnN��K:yBE)"���ޛ�Kq='T��8M��������By��5�J��h��̉k����#ѤƜ%���Ѽw1����O���`*���S�ڒ�y'hp!T���@2n�0�L�I���ڍҔ���k׮���7�n�[J��H2޼3�)�#�G��3��O�lQ��M.��B�<�-��f��J��h~I�v)�ϖ���)�(�d��f��I������o��g���j<^)�K:y��˧#�ŧ�'�+��Yd �h�R'�Xd��V=E1���+K�hb�i��V�^�4 T�BZ�#��'% �.@e��%�ð�3c��;��Ĺa�?ﰋ:��*U���|�3�"J�|��9��|�����DȂ�)��Q���Uw�2r�IJ�Š��[���I&!��>J9���Q���Q\�:�f��Rꗴx*e%��K�&����#�r�%Af���A��B�f���Q�G��+������J�R���s��l���8o^�y�H'5�9�/��/j���S��S��"4�˧��O�8.���=�#_|��}d|e��/m�K@@�q�~�����z���ӧOIꋨ8��Q��pt��9�/�~I%]9:5�_3.���)�h`��>	~��I���F.�~I%]EJ��/
�Y��5�t�ϒN��R�Lkkk�~������ޣ�J����^J��N�.7��rЉZ��ĕT��	�$=Y��w�MJsμ���3��~r5��    IEND�B`�PK
     w�O\4	sj�i  �i  /   images/5c3bf32d-6880-4472-891e-2d4d904f1ad6.png�PNG

   IHDR   d   u   7
�=   	pHYs       O%��  i�IDATx��u�\e�6z\˵�5��8Qb@BHР�� 3�0��6h`p��HBܵ�]�����ݧ*a��o�{����*�����9�����~������!�������Gi�$������(J��ƒR/�$/�UQU�0��(

/�CE/�����?����\|����A.����v��Z����?ᅢX"�ԍ�=:
nF� �W����a�CEUpKY'�SM�,��=��u�i4ô��gk�7/��.�&������/����a����>
������7Ջ��!�������Fp���+��?"Kr2�2��0V��ߦZw1nXMB��c)�N�k�R*X>�P�1SݬpBETM?	��+����F�5e�K��m����E�M�OQd���<���᧖:$�����>#�*�m�G?J�K���'mk8�����B��s��&G���$)�ʰ��������0�蔃�oXG�Op��)�$~�������J�Qꮵ��5aB0Wtۨ��	��]M��řH���Σ��e�_�ӂ�\�z���_ӷ��8a���ٗ�*E����b�p�#i�WA�����C���D	�b1���
��(ࢱ�Ѩ"�f���m,}Jq�c�_'���� ���yKÙ����)q�@R!��QUI��DQ�J����?T�<m��nL�O�4J�	�M��k�'O�EڕRNgA�HjlZzR��p<�3*M3�$� EY�	,=Gp�2����8	F���`�P(�ۉ����Ν۶�uW�0w�p����b�N�w4W�M�6� ��-8����7�T��M+���b<���ϳZ�XLQE0N������¸���;	����������t�V�+
�E	�)�1�!��0�0ܔ�"pAI��0<�E����t����8I�`�-�+�����0,~��Д���0�)���a�p�qJ�-�L�$%}����g�&�f?�`sO_������L0�D���Q;�������늋k"1��S?9�S�а�`�����������ޞ�m۶F#q�gå뮻}�9��$��ӧO�?��������V\;e��xj<�Hh��m[�~�𲅳�.(+!��K��c�COmݢ�	Ւ&R��vu����N��^TR�&DA4�\��O�:�&}�/_I��*�a4́=��ύ�N�>�58��8�8@R2�?y��Ҋ�6WI"��P�-I2�4���I��H����UR\VWwف�;���Ns�5W�1v�� �HH��]���O�z��}���WH��)���AI:���6>��S��_�4G1C�<qx��u����W����=�>�v76�(Ws��'��|���C}�,G����We�U�yf�/^oo?�)2E�_m��9}x�������i:v�����?vuO�1��8ߘh���z����v��W��~��AF{O�>�i�)�?�P5an~Y-d)�R�Щ��s���d�/3����%ͪ�b�* %�X\�$v�X,�A�$��>����4�]��y��ب�(���|V�iRy- �[(װD,�!�(&���j耜���ǂ�!@�x<���8�:�A4RJvw��ݝ�c�=GB�D�Oi����O��������Q����pNAuM]��3gC�e9�H����7�rG����}=奕F6%}#=��Խ���Y�_}����6o�{>B��Iw����D����|S
u��������/= ���� &3y�)�ewfNE�����f�"�<��k����q��Z�A�j�%7� ��*� N$K���9���
�P<���1��49r&TTD3�(���¢��H�d�����̞�.$���M\��lV�es��TA��p�EF���b�TC��f�'6L��qJ�Q?��(���TT^O�f�af�DY8�f��f�2<�0Y��1�
F&'�C2���� �DT���%4�L�S���� ���0,���r��jM�*�$� hF
R�ɂ*cp	� �L�R�")�<(C�K�t��ɱ``V�\���9�F�8� $݃����0Hg��	D<�a�2�6��$��2�C��-8ɚIV�/����Ь�UBY	�"�\O�����78j�Z��prA��&��CQEXap��IB�PH?1!�j:�H�0B��d���ыDe	��J�U���x8�%����3$°�ܢ����͂󉂜Tɜ���E�$���%B�p&`/�"��WV� ʤ�1<��?4
��.�+��e��9#b�EaJB��5���#������P4���41s	ͪZ"*P&�ba�A��Rհpp��1��Y��� �8o�d���������$&ȴ�Pun��H�eM�$H��HTU#��7�tY�&A���1��.i�!�8�IRD���������g��#�g�\�+��Zw]w����ùy3�.���|���I�����ء�N��d2M�[QVQ����x�� ����##S��^��V�����4o�u��'ϝ��y#��j��e+�����+��ǟDÁP��4g�/�,(��z���O��EH�DӴ�&M�㜿`ᷟ�?��ɳ4x�Ց�h�:��̜��'OQ���X"�,��ً��	�XP1;�k��$JU��R��DBb���� 10r���1aܔƪ��`)��J�N�c�T��ƚ>}:�?��u��t���TC�E��M��Ι �������;� �o��{6ݝY0��ң�>�����iӯ�\}MV��`�S]3{Ǯ][�{�g��s֬�6���ĉ��L�%+�g�mmj�`�Z�^�~޼y�~�iVV��ի/\h�����6��G����'���2O�Y�iԩ�Ǻ�:fϝ��'��q��N�5o�e���x�g�-\���8s��W�7nR�U�n�����	X5w����]�㑲�Yy%�>�hK����Y��X�Ap�5󵳯4[c�v�x�I��/jA<�/����m����{� =#��12���޽{g̘���[~ڷ��l��Ѩ���/;q���?{��3�<{��YP�|�����Nn���Ҳ���q�O-fS]m��矘�h�ڵ7n����S'#�P0���_�|���6n���<��#���E#Փ�z�q�f�Yxp��s�=248t��ީSf,[s�eKWj��������h$pp��%+�\�����(�Bw��]_�1<�K�t��<c��	��'�	����|����ݱ�֪Is��-���*�ƆB� ��(�ϲY�vQ(�B�/�"fAx�kiiL���@�onmho�W5�Z,f]ĤT/��ݝ]^�������r2 `��;6<<T=cLˑ#�8���hko�K�426�l��O>�B��H�'�f ��/����~��G�X2����J����dwМs��-<o��b����=�ޏ�F����������,�49;zhW[��ǅ�G����@eE9��������N�����o<��$
��I��m�����',�����h�]�i2*�HB@��1-!kZ"���{�X��V��_{������RkKg��,��Һ���MI' �  �+k�J�qȯ�
˲)ՆE"5,��tï,Ì��_�<�]�����rP�Ŋ�I"��g�3F�5����(�ţ�IJE����М�N�/�R8�	0B1���Q�����p�BqU�#j�ay\W8���Qith`�T��4Fa���ۺ�\۸i�����X<	|r*qI�깳���bq��nA&&ᤠ��&KZ�(�+a�.�e��E��- �.eEAW� �)U���K�z	@�ΐH&#�hz8*���uY�B��x�����F���:��H��v��(�>�X��3�~�v�q��dq���*�4Iut����@,G�Yn�#5SJpWT)a�`�M��HrR7/!�;09.���9���v7�DC�P8�rF6+	�0U��G��(��%%pf钥�u��y��K� � H�y����䔖����#��A뎍�\.gAA��f����"�����8L������L�O�U�� ( a5��2Y.P��a�Ģ������0��\w����"wc|$)�Ue�@;a*�TE'�L��X\�/̊D���p.Y��:%YA	<eʄB3K�b�Q�d�V�_��8,�k]V�!�AX��lI�<�Z����.lۧ!��Y9�fj߀g۶���u����������I�V��r��ymm-��\�����^v��s�ͽ������Y�{��g�y�	8���z�U믽:��>��S/���ݻ��EP�-����5���{�:ubwg�џv�3���Q2e��Q�H$M��aO+E�A�{Ys�����*:~��o�=7�.)�"���S4��6����&FÑD(�7�����=����v����n�
UW���-(����/�ʠ����Y�=[���0��Χ�t6���=��M<�5�U�D"���[>ҫN���������|���3��B�<���={�v�����[o|��7��Y3g�����>�Ey�}/�빽{�555�x���(���KǏ_�������>���+��b欺���>�p]u��6�
�F+��.�A��C�f�O1[
�[��b��gWN��nI��O�4kMVi����.��8�t�[Μ:�����?^��Ͽ���͸j���9�y=�]�}֌������O��)-)��-�M���'9y�uY� �8XIy�x3�C�XE��74֓�/�~v��7�����c!��`%Ay�-^��{7���m�v;D��l�F��<��e���w���������ͩ���#���O���ŋ���[[>�������'���˯~��^xndd�믿���@-?��;>�{����K�H��8}����3��wY��څy�s�����?:�x��i�p<�x괚U����l���;�UKK���+�����L��3����|?����5R5i�¥��5�Ccޒ�g����_h�?g��q�J���UN�5D�!��HI�z~K|ii��!����D�K�!�$&]��32�233u�衃G�G��'O2�$� {>w�a���}v�ܙ�W�p�!�n���ؾ��eK�����pȶ�B�|�|����{���k����a,,KQX�W/*����_��"$�� �kv��w_�|詧Qw֞7^0$%�1�Rld����@��}����Q���������{��?��fE�%��:|���s���r�M%�>���W_~�0�T^��y:��ϑ;Ş=�&�H�bIE�TI?���������qU�x��<�d8�q�����c�
�&�#P-7���v�@A����[�$9�x�Xc����8D/q0�'�'����%n�P}}�, q��P����>080cR��vVEC�"&�Lsh2���d0�i�s��^Eū'U�A�"	=m�B"f�@Qh>_�h�ZZ;��XoW���@E�M�H\@}#gN��7���~덷]��	��.���p7]0Eu*�����&0��4��s}Y�Q7�ԩS�C6�S]{�q���s|wwvf&xd8���i�=]6�R=�^\�R��\M겕����`�A���Tm>�z��$�\�|0]V�?�n��yB���j�X�p�W��o�9W-k�gy�?/�H`�EQ3�,Bey+I!9�Ԩ�p�l+a('p���i)(��Ugf�Q6�IHV���r3L6�պV�������D�/�+Vp�N�xzz�n\�8F~�Xz���]3sNn^&˘|~el�47�A�]{�Z�����A� ��tZ��۝p�pېN!{�#�^���XZ�3>��f)�H�iD�͒�����>���4�@E!Q��Z��p�Z�#p
����|��{jUAa�vg@��c�xO���قTb�oH��j���O͟S�b�j��8�AhE-�c1��\��y�[>i���X,`M�p�2UqJUi�LE���J���D���Ӧ�@e~VM�p����m�u�W��OŤPY5��[7��Uwu�=���w��~�����$�2x��w��W��XM�v��� �`^���k����S}��O?
���hd��ݷ�`0�[ͧ�~�ċB�����g���Q�a�ސ��F2���1�ܼ�z{����7!~g�]e���Zc'��d11NIR�I�r��U�=;���]3���fT�M(�i�K�3G��l���9���=�1����-�TDQeP=�=��z��!L�e��ZSEe9�1����>��;��־`ѕ��^1}��֖��K^�аi������/޴iӔ)��l�l���ee�@Ķn������{�2e��zw�r��;EI��_�
�B���o^z��z$��7������ݯ���u�]���ޱc��;�/Yy���S$��KOO�Q}�c�ʑz�/$GyG-Q9�ļf�6���_�����T=����n���=s���b��7_=sv_Nvֵ�^7o�����ܼ�%W���_���/<ݴ������`R_`e��rO<ք3|��%9Ñ0E� , ��K��z�FolHy�RiIŹ�g�����poO���Ƴ{~�s����.Y�����q/p_�_n�z���{����ٱc������IRTww���'o����81��?�$���n8}��k��v�mw3��_777�ñ3gέX�����/Zl��������ޡ����&L_��N��G1d�:shUz���ƕ>���#ޑ�&�ݻ��?����o��)���7/��ھ�'����7^���w�99��s��?t���H��֛gf����Jr4���E��J�;���Sc5s�=gB���О1A��J�. ��]}��],Ѥ��jcKs��SV#@81a�)�N�<�q���݅�z%�!����k�����AC}�7EN�I��g�y��������_�8.%!q�o�����7�t�� ���yQ퓏�hk�x�՗����{v�'��2��ԩ#�\t;[!Ƽ���b�G�ǆ�~9e�d������dP4���Ç��eÍ=��{o���7�8����O����+���f���8���2g�rj+C�KJǭhn8�ݱ] N]N����Q�\D���%o=���.UT����ػ��-�yI�{z�Y���Ȅas��(�)��� ����XjQ<7��p$aX#xh(��~ .,I��j��i�I�7�l�9b�ÙM�l,!SE���M�'�3��X��P��L ʔAY�_�|��c���������~Fu��Y54J�=z� =�*h����c
�1�#����̞57�w5|�jiq~�x�BQ1�!�%��R�D�@2\np��?*���-h�(����5|�)��|�as�&��̬rH���1B��v@�q�X0����F��{���$&�n�7�%�Ν���7[�h�!���E����<00`sdF#1��f���~#q<:��q-)J�������Bp<X/;����O�2��Ywl�CA�D#dF5"K�*�����W^�1]����<ށh(�_�ط�̋/�\��q�6�X!�0���:���
�99��1��W����zՄ晋 �!H"U���9�������B�tffe�[9ݙ�d��� ꦨ�=�f��!H|$Ņ"1$�H��KB������a(��@ ��%�ܱX'���a�t$�׫MjyW�$��<��/GAG5	��T�	�jY^Ÿ		�1�Ê��8�_@0#Nۀ^��n�b��N����D�~�7���~b�CY	QЋ>ZBR���Gپ���LG~������!Mo� dI�H�I�-�6;CJ��9��*�w��WY,NUA�{��_z�Ё�*��ꫮ���ۀz��W����G��=`pU�3/_����,7;/��7�N�e`�.Zu�*��r��9r@"@e�p�,�d�UW��������B��L��a����(�6�" z/��H<.S�����<�G�Dju�?��񂆀��:��_ IH����"��s�Y$$Am��*foKR��(�P�.��W=�b�����L��_n��(���}��ͻ�g�X�f�lom~��#��u7���sO��ÇA�/..|���?��3�
�=�������V�+;?��BW�i����#�::��[N�+�UV�g綴�j�0�v��Yu��}�_�Ά����]S4;�㓅�͜3���_�;��K���w��A!;��3]�&�f��88V����ڠ��
b�,cxH՘`��c%����8�!�P$���~rlԗ�7��_<M2��Q�P��(�Q��~{����+�c|E�a9ޒgp��J��?��XI{���f���p$; �Ï<2������{�I���,_|����������;n�i�;�xo ����]�|�ƍ�fͺ265�EF ���ց������+�W�;�s��g=��;����oߺ�;�k"Bp�/?�n�y|�^�����ȟ�[�


��a-�Sf)��X�����	C)�r�p^n� ��Z�"���bI$�qg�x4f�[�c�+C�F�P�X�����s��ڱX>�����$UuY�>�j��>�ϿX���'���J�X�;��唆�� �be�X����f766��o����������윬�u5Y�N�K��M۶m]�r���_O*��M�UTd�������������ςOY��3}��7T3{m<=y�K�w�����|�o�m��������DG��BPs���ڋ'Ϟ���:qhǡ}��|c�L����́���h$��RjE�b��\���� ����A�9��q��8j�b~���E���%	�VE�������c�BY&��a��C�pGo�'[�,[�}E�� [R51�Pz���e2��6$���!��ӧ�0&���G�h`@�=~H�(K^�؄�3DI�h�t�q	�a&��
=�C \áHkK����c�u� QȒʱH8�{� x��T;}Œ����R�S�
3]�~Ox���4͈� Ā��[�.Msj�0
�8NcH�LٌF'L3�Ɉ6�c^�%Q�NeRݖ"�2d�C�s�Fiz@SMIf���e��~ޔ%)�=*�Q�h��O���.ey`������,����7�M8v��F�T�agV�\8�P��klL�uoE��xj2�4u�E1����`hkG	@xw���;����j�Ǳ> 8�F�ȉ3�NSI��``X�FU��i%�n��B���}B����B�fk	��X��^�(m�*�q
Ì������jf���fi��O����T# �hvh���]Z7 ;��3�Q�(�[m�t�����*F����� H��$Q,��l������8Iv�i�n; Ĵޢ��x�n�L�|QIw�BRb�0p}N��vz[_7��##A .9�N�$Rm�*XP1A�x^��#� �I��8�4$��I�A�kIђ�ɺyz�R�z3��c81A����7_�7nr��7W8���8^��� `I�iFѨ�Q�b���> ���
BRR%!1T����f�E���ucy��ή�qUU`��+W3���fNAA���G~:x6O�{˭n�p��d�w��w�}l��l�y���X�haOo�`� |�]����j`�^�h^^qK�q�ӡX`yi�;�f��S�P�32��77��Y��g�b�4�"h��Q<��0����LOO7��`�4e�E����eͭ��Z�{���Τ��hE��\�@8,�����g8��@�`BL%(�cR"� 	U�/6AkZJ�+pz��E��H$"��($��<�_��7�֮�y񒕍M]@���������|��-Z���^=}��5�Y�l)d�����+V���K۾��ɧ�fgg�s�=ӧM۹c[vn�G_|���o~��mAD&N_>Ɋ`���o����s�:Z��J����&���/�m��09w���VU�9kԇƓqD��$7O�r���;��dde����\Ӆ�������+#�����X4L�<o��u���$��i��4)B�BǮ_��ȷO-B@�����/�b��z/�Ū���.))>���ݻ��Y��{G���C3�,x��O����Ï/��bGg���'���?�[P������[��2����7o�p�]w�_� ;+��ٳW\����S&u�����-]�D�v�#;G��$o͙�`uqiE$���-
��O}��}#=���A��ļ���j$5����K�{y&4�).*�(lxhx�7V^Qi�Tgdf_���"��G!��gw8�5<2�����##"yY��F��bF�ΪJ��foru�75��L�1��4�B/a���?"],�u��8|���U��1�������ά���o����6�s^��J
���sG�n����{WgOy�x�(8��}a|�������s�5{wo���wN���[<�ɻOh���X"�?|JM�M�]�U0���α��p8b�X�`�d�f��b�.��fI=�ˌ��h(��`2[Y��q���@P���ё�l���L�m_B��Y##�0��l�f�(bM���@���(�1��aω��K����F��$�,M_�H�'Н�?ee�������c�2FŲFHg� ��6�8�x��)@nA�FƕB�JrB���_)�VE���-
wwu��f��	���Ix�=���n�,D��6��Oz<�����"�pG,����I��n6r43�]CbbTA�����x8#�I�%3�t��F<�D�a��QLY�:I��%݋�Z�P�V0._�iz�?�
S��a�st�G���ev��h,�A���*�3s��-���\ʆ�g��r��H��(PZRJB�h,((�d��0r ʐ�}�:6��R�!��u��4�������
�����(���PA�D�����1���VÄi���P�e�h\:������5-��@P�Ԭ����9r�b^L5�J�0e��(89�h�R���vJg ��QExah� G;ͣ�2����&
C��?zes���i�D(2��WI%A�B<��r��H�7;�)���.7ñ}C�BQ��Ac[���A�c���������@'%Kq��R!���,��^�0T4!(4�a3RD��s���@V)fpEBQA�#L$��{���bd%J;mv�^tSe�&��☬��"t�izwYE%�j��F�ca:6#�}W(��Y7YR�a�Z�{�(�R�ӻ�U�(�"Q��q$o՗���U���<I�%ݳ`�#��qp9)�բQ�U}�f��+@��_��p��ɓ�&S$.)��|��ӹ`��#�v���o8!��͜kwXf�T�� c)����/,,�LC��Y���ͽ���2J�8��Y̲F57wgfd4u�b4�BI���Ѓ�gJm� ���&a�>b��"�/��I�ŀ����0�ri�0MEO�z2�t�H+Ł��0z9���(�RԀ�a� 55��������To:w�\mm͕��Z|ߏ;gT�\�b��b}�\n��/>��guz�UW^5k������p�Ё}O<�ȁCG�z����ݛ�7������у7o�~��e��^�S��M����;��xv�u��S�}$v�+6��ϰ�,��E�/?���m�}��{��g��@��P43KH��g&�G�)��8���8f52���(J2zjGcB���q�xB����a8D���O��9�c�(�_�)�"�	CI�WsZ��'��U�l(��#av��-N�BDKoQ�X��x>ڲ%3õb�򕫮�����o����];����|�Ms�U�?p���h$�����yMa�at.^���Ͽ��7nܾ];O��mLIw7d�U<��{~������tm~��]���l����ꇗ�՞��ɕ��.44?�ǯz[6�q͚�7VM�u����Sj���ݮ6EƼ��Ĩ����M��SE����c��	�q������q�r\�?��ܚ��-��h�>�b�PV�M־��)`w���z�� �rZ�W��K�ķ�E��I%�sv"�?v��8~�sss�̞����Ï{���;~������h�f�NU�Om����;'����z�#欬Mx�x��TS��_��ç������%�WUU����?L�1���s׮m��uKSc��	����?��ig�ԃ�wy��N�>E�L�x{o�ѷ:/,_{�M��{��F��b�4l��z�5$���j7�	P�d�6\���Qo�/���hAa?C��L|<��x\�=����s,��ĭH4�Lz����l���F� �Ǵ���4��隵��F�(�&E}cGZ�V�/�tc��IRR������I/P N���g�����4&����H:��hMk�8�Q"L6���l:��FB���r�'	2� .)���x=G���)�ϥPt�k8nU�=���Mw;{rP�	�0)BE!x��.wF�?���ʅ��u���U�K�!��B 8Q�u������
f�70��Mq��EB�Nw'
`�9T�Ф��g{[�--�d`Yo��E�d1:��a:#��bSe�tSCg��kݕ�E�XR�4��IH;TZ���0YvvnvN6���0� <O&5��43�H�r�FgIٔ�I�%p���pV���L,>c|n����"[DDDH�,LN$c���h��DA�mf����pP�tz(�X�Р�	,/'?�4 ��x��[�i���ċ0+A�8BX��#M�f ¥W�ZO��Jͱ(�;4��fM��^qc��@�X$8����A�89ld�382��X�ԞP�Ҧ��E���b�Q�zu@S�^(a'#�p��g�1��ޭ�D(�2�PƊJ_y�h�i��H���rd�__�� �MJ��7����7�cacL�9YR1.
���2L�Yf����X�L�@��r?���"�޹�p�A�$��gqԄj6D g�}�xzs5��/�!�f����M��#�V�͉a�Vy�AH�
+/�sFG�P�BR�@uk���+�0�2�%�Ko������L\yYU{ǐ��h�&+�Q?�gͭP�(at겕����[V�ߖ�mE1�c���-++�ț(�b�L�I�zf4�)F\f̒ScGz)ax�ĳ2�{�_^Q �
��1t��P5��t��BP\�EqXTߤL!�A*"�"(i���9�G	�-	fE0E��z9	1�SW|�-�z48�9Q*�v��4�-z]O�rT�D{i�n���������������jķ}�)P����~��g6#�2|�u��og=N�m�{x�U�eZ�@C��M*ND���܏ڍP�4y�]o���P0�G�**|��h�����˿���"���ӏ����U�#$�a�0m~��5��.[uÑ�hj�%	�_Ql�@�/ j�Й%�4��8K"�zF%x8f��(��Ao��T.��=!�	q��T߬�WI[R4���cYʄ�1�Y���[�.w�I������O.m�G���|���������7���t����ٺrպ�o�)`���G��\�὘��l�FK�	��"��ﺀ�����I�-/_vxxDN_a1����-�-0�y�e˖����%�JV��=���Y��ͺ)���¶o��45���{s2�[�w��N_s��U�O���XΨ׈����P����%Y���B>_P�:�&����z�c?EI�D��(��Rq�8:��'L�,���3V�TV���~=�HXf����������l�P$-ݷ�ֆ��ש�)�ggg�O�?p��Ͽ`���h����?����/�����H���7J�8�T���n�Z��X$펷��gw�ϟ{�cҺM�5�ܙ����kH'�*�ع������3��Թ�߽��@[B���_��xͲ��W���;Z����x���\[k�ő�d�5��b��v��La�ƻ�No�ܱ�����9#�����TIB!�l�u�8*��/�J&�	�e��M�>�$s1�� ���a��*
��츈L�Y͚2��c�&ɉ[F9$
୩��~��O�m�\3k��l>	
�AY���8ZLT�7')�`%q�U@0Q!��(�F��ao")c�����W6g�RttH�����(�>���U�מ=�?ֶ�SPc5�}p�W��U�'���}�&�X4�CCǖ]���K�,�2�*<�����׿����^;|p�[o�F8�$Uno�@�����������0E�AXjI�<{����u7�ZX�w�;Q}��KvӀ�	��c��|[��r](K�G;���d�䌙�g% ~A�!?��c��& 2��q����L;	�@��O��#��)u���ߏ�BPV���'�c����9k�h���
���3xr��� F��9Y�hg(M՜6����;��#q�H$�YZ�
FJ
�����l"P���C)����P)�Qx~I���3_xa���#��g��y_8�?�g��
pT��������G�-�S��c>)D�^�ב� ��ӊ���5�]!��ðtTx���kr���Q���]*�蛁��xD����x�2b2IS�"��Q��wɋ������X5�	��N�k�i�>q�C{*�qP�zE�8�I`H� g�����8��0�{t,�Q��H 1,Kü��̬p<j�������w�bx"��l�D��a-I���XR�v�JX ި��p����)��c��%%�,�Q��"ɩ���za"��J���l5� )�ሆD;Gˊ��T��%
r�A�AёQ%EA���DkK��i�-f3܆�3g ^3�d|���r�u�+��?|��;8�����B[�gu0�������y��Z���B�Ar8�@a��`$q��&ȱ�0�-���3���%c��j� ��JIZ,��Ĥّ��K���P�$h�ňPL������D�fi��N���SX�FC�x�iK2&�RzC�F��MJ��@1)�;T�DU�Ԩ�k�����_�Ԛ��<3<<���˟]3��	_SskAQ���-X ����t�M��2�4�#F{����}�Onv[��Y�v�:�qۍY]��fm��Z�DAᔚ�9���"T�����v��6�Fk����1��}�^����-w�T�_�ܓ:�}_UU��]��ɚ���y�"��d3(A4}���k攗���a���qeA#`(��GeuN����d����HG�IMR�B)!r�����aQ��%� {T�J&�8%O( f��.+�QzY�H���s��675����^�|���'�_�p�&�{�}������c��������WL�t`ߞ�＃`�;�����_�o������^���/N�:S5����o�޽����[q��+��������?��?n��+��w5卖��3!ꇺ·i�z�eEe�Z�����x��"u��qw�'�ify��dD��6������bA���9,cMƓ9c��H1Z�1���<�q� ���� ��{|.I1�L8Fp5���}���dX��3�v��E%��Ω�S��S$�
�WgQ�a���t=����h2F���6�5w��5k�?���u����������7�����>�`cc����t��ɾ��������;w�mw�ʰ�[�|������H"�哯����'��Ӈ���Ѵ��=m�P,𪂷b��e7���֦�m�G	Dr8�!Aimͼ5ɸ ������|dJ�U�4�V3w�r��%$���Ã]{��N�_9~ڪp�P���M_[�>�#b	k�*fO�C�X�����1M��E��U1�/@�u�_8{tx(�t��K�no�
�T�	�z����J�dFF� >''��v�N|�������'�����Z�W^^<��>u���o��jժ�;��.*�1�mѨ����������j���c���ѷ��m~��U������@��"����r����w���`���������a|c�P �*&�sdN|��g��Z�8z�/Ir0�i{k��wl���?�����n'EHz޾k�o�[4x����==K�4C��ٺg��9'�t�P�qZ���;�&N�7{��ޑ�]ۿ<{�Ap�;cǎ]y�ų��,�4'�b�a��{?�������;����b6� K �v��5��i�h�d�f�U��	�	'���L��!O�*baYF!�����p��H`teYN���I�C`����@��~(�e(��FCq��Q�z�zz��x�F⊑�-Nc�`W����Gp#k�7{.I32J������I�p�F,V+�0N�<��v��UD�z�3N@��%&ܩo���Ձ��g�bx�34ǘz�z���?�	�M��ϕ��x��Oy�$.R(����4��C0c~�DH4c �E�Ee�U&	Hy�t�K��8�菞�8�5\�
(+�������s�<yF�lDV��O$*vtT@��q�lfI!EU"�ynО�	�tC���^��r�sg�溭`\{V�����'j��#�F�8I���`�=@�Vџ8E��08h~�$���?�D�hR��;[(�&���T��7Z��/j���}H�/!7��l��՗L�����4���f�m������0}����C)I��� Gꏦ�X\���B�p)�����
�b1��ɤ �O��j�h����r<�(�T����GڻGI6��U�.�'雪�p,�M�E�Ӧ�y�Cm���}W0"�9L��!�6H��}���<���جF��"�OQ��N����0��+�X���A�d�͏Hw4�u<m�t����~��aA��״I�2�N�海����'.�{)KKKV�\a�Z֬�� ������-]�h���p�ŋ�ٳ'�o>#��DNN�W�4�mKV���o�$J1���)y�Si�fs'�U�8��e����H<Y7kNq�$�1��h��ĩ6O@����*
� q���py
8��tiq�,�f�k�I��U�;ÚU��b�@�	���R{�d ˲�P�cIP��39�0n���׫7��%�S���i/>zMo�M&���7m�����-�}���~��֭������-�l����#G����S�N�f��ښ�?���p.[v9���Ϸ����bդ��}�cdddٲ��f�?v��Mw�|�m{���{�>�����ɳ��(éSG'O��9�O޻�K�qL�[�p՚�������W�����-*�tX,6K,��p�2�L�e19:�c��W�F�D"��_���۾������
���,Y�����n����}��N��I�͖1}ƼP82o�Y�O=���x�%�����v*���,���z�@��uQHϞ=p�����{�1�UX���o�=�����~��ߝ9s��=���2cx�ȩSgW�^��#���v�����N�Ц��E��p�z�����+���՗_$C��N�[~����5�z�($�{������%���.�r�ĩ����_�?�}	x�f��}�[�ԭ[�%[F����`��Lvw��<l�$H2لL2���af�$@��	$3��\���|[�-떺[R�G�QU����U�13�g+~�%wW�����~����?=�q�Xx��i�~����L���D2����F����	W_m�Z|���=+V�m޺��o������T|��������>	oںk�w4���ںe������sFK���{o�\��{�-f9���9�.t���ݠ3��t�����;%t�H�V� ���#N�u�����C�^�������3s�b�B�VG�����w��/�"�D\pW0��^z�c�+V�x���	�8�ň��՗����|��G��8��B�<}�l����<��oN�������.��#V��Ν>�ٵ�����|�4�A^���T��t&��'��MOϩ��tQ�����y�"6uG"����5|��G�I�w�}��pӊM[���M\:�3�l���wtjj|����? Aǣ��f��/.�]8W�mp:�Ru��s��u�uRBh8�7�N�zۣ�8K��ɯ��J8�"%J��2�I�&KR�U@��ob9���MN�(��S�ݢ�����hhb�����9:���x>\�tDgR�d$a���,%�*����n6�ѽ�l2�t�j�4��.?v��\v���K��y.��y6X���j�F��G���憎g��Xx�j��j�c�y�͚���)�ASQYf2'&�P��1&��x�ť�e��kv�����,5�{'Sr������PE�)�Jv�
�
�j��&)�\��\�$_�'s:�36� ���G��mm����&��,�����M�H���a;J�mg>:�L��T��;�755�gsY�����D�nk�1�,���r��òj���o ϲ:$;�"LUF��VC�i�^5;�N�O�,�z�A�S$��d�Rr�R����I���r������I\�&芐�.�dr���b�k˻�E�� �Jf�Y�%�K�	d5����y�+a�� t�\�E��g�T�����X&���8t:��Ȥ^����(d�t*Ue��"��lt:���Zu"�½���.������~1�H)$��rS,��^��P	�a�j���H��3ad�%v��f� ��XJJx(�[&�G5֗���c�sdbI+Ag�oJ�"�!���%���R�XD��B_~6�b��@��d���i�q�N��u���ߟ_\\�htP2��p���n�������ghp�H&,���u���<��}��&�
2�e
{��(����WTU^�^��|>N��U(�J��X	 ���\*��F�������|3�\᝷����Ųa�L&{�m{���T"��1�
| �� &��9�Q�Vh��u0F	p/�]�679��0��`R�Ӑ����|^Ou�P��nބ�nd�~��G�YèUJ�������o��x��x4�uϞ��[D$v˾}k:;�}�����:��`UUn������?<t����=ϲ9����v�n>��gO���c�	δ���㞯64�b���pUx���/�'�X캻��_����K�9Y����}�O�=��ˍ]6o�a�V�X����+��O}�`���%�ںM���ro]k�`��R�6g�Z�zM;��؜گ��w_y�?.�6z����eUm�i�oj�����7v�'�
�rS�`w��W�G-#/�PTWU���I+م-l���)a�����X���҆���j$�\n����<x�^�˵��%VC�޳e�&R�+u�A�e��Gսe[}C���|{{�	��TQ������~u���RMe8&O���^�i���)�+�4W�E���*�����rE���躍[zk:�!��Uh;ve�h�TU��C}0����---o�q8��v�[E2EKy^����x��]{��Guu-]�6c��lh�-7ϵ�|�x��}�v`.�r9�)��2�ZZ�.���3/QRde��1�6�^SS���P"��H̓�^H��9�lI&�8�O��W���6���t<���h-Rخ���$Rd��2��p�cn�����
�+��yҲ�@�ml�D��3;1Y��R��RIݾ���r<��R"�R޺��5-��T*�p���UU��<HB�Z-�*�� �2F�������W�H���?�%&m����ઑ+H���D]X�&\O2��8Ja�R���E |E/J^ �"k.K���(|X�DLMʾb�DX�*"��CT"�	�"���_��oB�-���$���,�)t0@kLFB�Fp"II@|�
�@d� �{ܜ�-).K��?SZ�T��{�U����OI��^�_��*�L[,+�.U�?��E�R Dx)(E�_\p���a�DT�U39�b�D#Q�1���C�xe���;o�����Z�F�P�~�NW[[k��GFG���T�m"7�(voAqC�KX4�s�Z
���HEy)_��K�HQE��I�	�1�0`n8��N�R�T&��E��̈$�7��pL!��mV�B@:5B�u�����h�d2x�h��l��TO�����uUu%^���q�ƍx��ʪ
ߜ�����b�����K��N��{z s���K������+V �޶���`���C�a��b�	M�7��?�����L$�	�����~%D�H����yK*4��tʈX12��x0�l&M��2�̈��<��VA�86W���?�U	��:3o-�Q&�H�V�aylQAG5F3Ee�r�mA��_��"�ϕ8�v+�o1�gf��z��~td~��Y� ����+W���dR�T�۰ojiE�
�z}6M�>�H&<u��$�_���G" ��h<��FY�����F� ��������}핗��_ h I���(�o4[;;��������J�S���f�����HL[�0�NtFp�"��u.�_^m�k����n�@��Ļ"/��rF�,+UR�H$�fRH��n��6�a�l�Fm���{L&s4njn"�*R���B�0�;�2�
E0�+��@�U�^�wP����P0��ԤV����~5�ie�57�0<4�.s��81��X��}��2~�����;\�c�"������M�,����xF�o�41��D,
�B& �_/�uH�éi�(*Y�]*�vJ��̦t:1�_4��k∾�4-p��tZ�?L�ŋ�/�V+���3��e�b���p8���h��$l�X�T
;�[=�4 N�d6cz!w���wΓ�b��z1�\�%�����&�ov�:����۰I�������d������g�Ti�r!��ع3ǰb8&U���:|]/x3����q�o����w5E��{���O74&�lہ����>{�sp���L����A��;~nvzdx8���4���O*35����]��]}��Р�l��� n�z�WF���7�!��F^a����������hDb�IAa/^8��� }�C.luF���-^g(q�|>ː@��A��T
/fw�S����9>�S������Э��F	��ߞ��W^|q�ޛ�0�Q:_㩱;l�P�����x?h�/����j4�����Q�?:KJ&�nU�R_�3H�)E��Ґ{mmA|A-H��d�T�S����di�[A)c��bu8K�l�А�M�\�r`zȇ����V���F�9�I�C�u���'<7
f���<�0I������~���v�槯c|�����ψ?���/���c�~��
�J�� ���:��/}���-�S[�
��	�-i�JMf��j��#"ㅂ�pUU�x��ٙi|^�Tss3CP��A�\:��0J	x��� $ NR�C��Z�}����$d�K.]��Ё��k�M��7��o��z�����}�{_{��˞�s}}7��axpx���6�M��/ճ>GR�`_���僅fgf�������]�ܻc�nᔎ<4o�h���&�+��TO" 	�㱘�7|�p�(� ��a�|����8���G4$�L��}���q,�K�3��
��{��dR�҇M`=��Ϥ3Sӓ�	���I���G'�*Y(�0��ߵv=������k�Ν�GF�^~��:�N�q���?8޽yn�,q66� E�Q�8��Hؿ>�k��ï�v��8pe�e��--�Τ�##t�nl[�RiR��v6�#�a�����X<;q�RK��Ѷbeiy���4a�P�mvF�^V�I���0� ݽu;O��P1X�����T.���@������y��)Ku5	�����{��[���K/�gy����V�΀�O���\��ӧ��5�������3�:�y�M8��ǎfh��ɞ��W�<�t,�T�5B����c��_;w�~��7���_�z�m;���m�[�q�O��w��ֶ�UZ
��L&��y��tyE%!ig���~P���0+
�_�Y��.I����US3��H�g����f��lY����
-GFGv�ك[9]%J��J8�6ř-�X$��ˁ���=�;o�Z\H%c�R�3�MMO]�F��z6�_�����n۹]��q�1�8��4�%������-�(+�b��E�(����.L,p�w��/?���n�Z�w��׿~��W�~�pcc���"�Hm]���� �!`$��4W%�h�l.'K���;v�k���$�mJJ\��MRB�d�*��h6y�ut:m�h��&�B^��!���Q �ڬ6`�h$BNP*�o����r,CĠ�����0��_�_@>PU]�;8m�2�S�&�٪U����W�qǁ�CCC�=���������A�t���R�ka�BR }~rA��nO��V �s�/�d�������{n� �� �#���������RGI푚���À�W1��B��,�!�l6�$2�ޠ��jeG�L�'M_p��e�PI��Q�ܥ�AL���s�d*����	�H�H��+ƇD2�����K_�r������_���z����;�ϟ�{�7-f�\X:�8�s�[W']��<͂G ����>�����,��z�W�c�eAY`2��� ����kM�����`�\2%�thp9�U!6s
��r�7�.��7.�$T0��%��]]ds=�k�cW�tt��,U�����z�� r���Z����A.%j�?0��7	G�H������aI�Y��U�W��/�zϟo[ٮ���%9�욳���/~���~� [��'kA.\<��������`z�/I#�5�m�t�ԩ���ƽ7ɖwKV^�'ʓ�D����"_ذq��/*1�,6��zC@����$n�X���C�.���n+vT�⑥q����ק/`��Ǐ��t�u˰�(�0��{v�Z5>v��>�E��<T% q��UII�����cpE#��:�UIID
�k��o�z�S[�w����F�ٌR�>gx.@���*-,, v�no>0A�]��l�(,-�>����F��-�v����[r=⊛F��`�۾x�݄�T�^Ҹ��gΉWCC}����^{�B�p�3v�*u���e��W(~�>k֬&2�,n�r�G��n� ���b�Õ�Kan�ETUV�L�=Ҁ�~@��X�%⋐���
�x!9B6+Ҩ(�$�e]b���R������ٌ���B�� �	O|q��B�ݞH&�B�R��^��"I4�]Ib�)��!nF$͕Ü �Q�$�*�D\,��^o�ij�g��	�/��p"�А,+��!�����*٢���Io]��TQ����{D�
.\��.��uD� ���ãǀ�^!�۹sϑ#���X���r��g���Ɔ��T�z�W(�4�j��F��+2�,�'돰�"�e	�2a���J�</xf`B��"|v��*�[$S	<&�TR"�Tx})9����4��pB^��E�#���
Rﬨ���N_rĜ?@)EXN �B��	��
�H^<w���Y<.���
Yy��:v����/�]ܽg��˃�>�{��
�����ۚ,F��|h��࣏>:>1�s����?��O�2�]yI�JkH��R_��{�<��<��CN��˙�o�ش�`��2ɖ�؅˗�|�m:�.�̶P4b��H�XR@J����ꚾ�!�͢Wi����d*/7���t���2F���0S�+J�ـ d
�)Ɠ��j��
���e
,�[m&G�)%�R��+� عOl�����ѩ��G�O��ӧ����#��'��z}jfi��dE����ѣ�}��|���7�z�����g}OeYEY���8���'��W������_���޻}3�I!����ϟ�cx�[��T�.$��^8x���`h>���K���W�55��#>v�x�Ӻ}ۖ���ZK'M��"�A�C_�-U��DT�x�Lhzv�����X�A2��P$N��j��ɤ�no��}e|*0�i$�]K���TX�\�w��ü�ON�)��5�_��nw�#0� �ѽ��烡H,���]:����w�w왛^��������G��+tJ�!S���k��u��������)�fkd1D��k6%;}i�sæo�SG^���z��w�Je6�)���r�|`!�f����t �&�m�Z��,��Y����c,�)�3j�F���Q��pT�a��V� �gy�6�*�Ӿ�lE���_�R��F�Lʗ�7��k��*�����Q@��DXB�#��$G_��~��mٲ�wO=5:��ź7l��t(Nf	O9�N����N��NO��f��:��Y�Ŗ�`p[$@���㣉H�n3k�Z�e��c9N�@He�"�g�����m���J���p�z.�*UZ���E�{�o��Hx��������s���3���2霟q��N�Z����ʊ\[K%˱��f׍�O��������dr�W2�+)��L�S�T�YUj��i�a�j�F��-�,��#v���e��/)9��)��~��P�ފ�����b.w��?�鿂Iq��b1��l�LLE�2*I�����)T7�o����cO��#�8<Yq1��nkE0B&5)��޺��9�逴{Kw�����8]2)R�l���f�>w�`6�J�N���v�ˊxG�xY:��k����"�%�$[�Z� YSc����ʥ0O�V#���c}<����.���r>	��|Fht���br��٠�y�r�h����:�Bq�[N_�m_ӹ~�ޞ�B-�vn\;6�H�h�V�?���'N���~#0;�f�+�������]�*P4��M�{�/��җ'�O�<��HA1w����h��ĥS��}۷l���~;9�CH
��z�ZkJ�,����t&�ܸm���(��w��;0��z�4j�H��c0@��C�+U�Ÿ\rr.yi��*pgJ8;3��O~p� /��p8��%#QL��*���77QS�(�+�Î?[X:�V�T$)���	#��67�`s���ӓ�{vn�Z�>=�?����4�X�pJ^����hh���/<�|Ksæ�JR��R�Tb��R>���~�W�=������V��_��%<����j�7�o�x"t:�-d�����p}���/u�8v��?y�?>f0�檣�ݱ�e1�̇���Г���t��*3� ��:}��0�o��*#`�P���jߵ{��So������x�Kg.��:Z,��+[�9����^_[�L�6�f�z#�$�1�ݹ��\�XI�T��u5�d��_?Q$��J���[�֌�O������mMg��b���L� #wMMyﹳƭ[��i���ˮL�RJ5���h�޻Ko4D��Қ���ڏ�0te`>6����m����
 ��Z���tC�grd4��:J콗��tMe��b�!b�C�Z^��y���Eҽ��� h�]eeE&@�\���؀�����l2��(J?nf[��n��x��Ey89��L�R�����O�֠7������H����&}a�W9&;48�����澯|%����K����K��+/-�-c�?�ԃ����[B��p����59rLo0��1Şˣ��Ѡ'�lfҧ�j�֮;u�����L�Q�Eig�d�oP��47�^�ڸ���>�S�p�1��a�KU
�>�*�6mA˧rV�����J�VjԹlF���=�/TWU���g2��k�fg�γ��S㦤H1�*ɟ�,�ҧ���Z�A���RJ��OL�����y��I.����B����%Ȇ���È')x	�a�:��Y�o�^��H�5K:E	Z�3��GG��;���|����Y���׎���\�f��\�:s�¦�]jX�N�N��ȉs�3�\� �
��J��7X,ez�B� �l��:m���P�j�B����'ɛM��F�/@��mju��A�f$k�q���l�}BX��gXe
	�an&��Sg?��D��2��	��z����UJ�?��w�~�i!�,
Y'гV8�ޣ���������U����$žr�"Ei5�'��-rcKK.��|ZF6�
;>��N_�5����bقZ7,�w_0[����T&��գR�(r����^���脌O�"�W%������Ǽ?�ar�{��B31�T�ʬj����k/J'�|!U��O�H�Hv�rM���~ARp��J��_��l�U(�|�g�|�#'���`)��5��)�b���؜6����e،�i3����Ɂ�	���juj��)O�xQO?�<�Z"d㸏NO�C�Bw���ڵn�M�\,`�b%�K��L�]n�.�k�C&�v�W5�Ig8���L&�a��uE���/��S��?�S.ǘ���ښ�|�_���gw�֥r�R]Fh�J����Z0�p�ཀV"M���J���E@����9���0��<�|A8�(=��N���܏\�A'��d4�7t��J�D�U*�"�8�d�A�J�Ti�7�%J,ҟ�Dh+n37,W� y���$�@`�(�˄cinn�L	풼P���رSx ��`��7��o�]�o^�sLv.H%"�[�s�}��_��m�n�5_�,FZ]����6�E"�쵻�k�<p+�t���א.�|<X�L��r���oN�Cr���7���2����E�ᖇ&����/��Ҷ�uy��K�$��"��S�U&��\�K��x�R��i}�%X�vb�Z���(�� ��9���B�������
�b�B�����V����[    IEND�B`�PK
     w�O\	��} } /   images/bbfae99c-8036-4c5e-89fd-a87441410720.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs     ��   tIME�#Պ�  � IDATx���{�m[���Ƙs����8��GսU���袍�i�4��A�("�q�6'9�Dq��E�HEVd��HX�d���&�Н��g=��n�}����ךs��?Ɯs����{����f�J������k�5�x��p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8��}�𵂪 ʳwQʄRZ����k��{�Lǁ�%O�h	*T�J�`011@��#�QD
*B)�@ FI�"4"L�Db4��L[�>T	
4AU0����11��*��J���N�L� ��m��l@�(`\m.@aW��7W�G�|������%���<�Ç?���p8��h��@K�J���s�H��K���EFi��_j��R�kh�,A	P@	`   �jQb���!f(PA�U{�B8��W? � �FE}E��z�T�0b��P�t�>��1�yPr�P)[��7���I�����>P�+��T�hT ��ۻL���J��ui� ��5%Nd?#��z�vH
U�w�[��}��rV)R�""�%' ��f�v�U!�bs�!lJ���x�/.��Σ�~�S�����G����7 xD������%b~�]  A�=��~l�,!	"bz���
�*�E �
$S�
t�Nb�Z�L�WaEM����DՀ�Ĭ
�h�AU���!7�(���?��˯���1(��a��%�۽�����]���$���}i8���U�5�ժ��T�[T�GE�C-�J��eC�����	d�VE�RM��F���dQ�liO~M�?'0�w^d^�b�Op�x<��L�$����3x� T"��q���/@%B���w���w��ڄ����k��3o������k�q����:Eӯӳ� e�n|�Z��	U�M"�7h�Yr��((W���� D��@U�����y��䟽��� �6� ���X��D%"H�T�(�R��0+���	|KLO�x��8L����m.��>��m.@aa�]�%����P��/  �Sm/�J��eM�7h.�SD��J�$_+t�RM��
 ن^X�f��@�aJ��QS�t��k��纽o>c8y�l�BqĻx<������{MH��sF����J�v�������U�v�+��K�������]^\��^��������ԟ��|�^�/�-�p����; t�0�>]=����_.���FD�[%���P�)	R
b�K)PUÀq� ̦���2���_�+t�;������2{��W�~N�D�DF���k��q( �fB8�g���90��2�d�����q��o}a�X	�@�>�G�ᗍ�VU����n�./��'�����/%�n���Z�K*%��Pɦ�T d�ά��H��Du�Z�9��yeӕ�����}N�]�v�W-�~��;?��c|���	s)(���QJA�fB�C`036�`6q��F��,��j�@�.�q�}�_o��v�y�~���g��W~Ƌ��Ǉ��q�`ڿ�_�o~��-������<�Β�o�o��V�|����D2��\!���!F\]_#�(Q�W�Y7ƽ˧3]oqǕ�\`S���"ZM"�� J�jTM1+���y����M`��P���ϙ�gƟ��~�Ke�q�1^\!��1��,���;�������/b�]�����U��HI�Z2 ��"	���`^yۨ�j���l&��mH:��@��l�
^P]���u�{	@��9��s��{<��s�7��.���L@��i��%c��؍6���1b�<b�#��E�0�+l����U�_�������b|�_n���7^^���, "���~����g~�G_�2��W����O�����%�v��7�i��|8n��[���R@*��PJC��`�!9���E��^z�U쮯�(��RU����� p� )�z�5���5ki_2����&�5���5�Ye.1WEO�����9
�'����e~������3������1ݾ��}�������o����!����?��9�.��T��9���I�"')�
�慢�B{�g�Z{�^IU��mt�Y�8��ieٮ����$��qԮ�0Q���.~a�9|*���ÌL���9�((#cF�P��BDĆFly����.�<`Ѐ�p��Kx��|}��[����/�~���T�O@)������W�������~�ǿ��y��/a�yʘ��b�]���o�Ͼ��2r�~��p��3,����4�P) ./v�$ bLsƓ�^z��x�ʫ��
� "���ӅA<�t����<���])U��kH��Wy��P��]��� �r��G��C�U�/J?�!�(��#���,o�M���#���#��p}�����u�П���|�G�|���������e��_�|+��*�Z��BHU��(t�ͧg}	yK���*3
�U](y%@hM߯��@���a�y��`��s����N_�8�@IAA���`F �!�b�
��1�6<"P t�J@���p�勏��W�`xTv���8?I<��ƿ�H���4��.��C   �7��+��4�i�p�x�xx<D
�:�ߖ�߭i��A��8o���� � �3��Md�H���#��9g�./����g�N	�^~��������Č@=Q�z�I��;:_���LV6�^�l��H���_׾6	�<vQ q�P��@���Y���q�� �o�D7x�c����@�P���/�*��A_�����폐����_�^�����Ayz�� � �J�h�V���c��S�w�Vν~I5!�)t�j�/%]š� 뤸��P���x=@B"��%Ct��@Q2��j�H1�Z��JI#2fd8!% `@�� 	!d��������F��:��?����R/�t�{C�o���6=~��v��o�~�qw����AU�RP��Bd�p�:s)�ó�?V4��9�ߍi���p��·m)�I��{H:@JB �%�'H�(iF>�Q�H4(�>�@cA�	�M7�i��;()D �%oz����q�9t�:W�dg�o�;��#����u��I�%�X�a���|����(�߮y�#!���@o}���8~vs���[_�N
��~$�}�y��޲,� �Q*��9�%��kXӀ2A҄��4�z�P���oYY����aJ�E�*��j_�*�cYXk�PN��l-(/4;��.�S*7����S�����	��IZ
� H�H�.� K-��"
5�d0�6؅+\�x�W.���xix	�0"`Ѡa��4���g���e��2���x��p����-!����n��K�u����9��3 �����͗���o�*2��O�\~_��o���O�i��N��y"�3Ho�Z 2!�#JN`"��9!��r�0�nn )!��8D��r��E@q���5~�۰���FFV3#R0Yc���Q�.DW��ޛĉ�~��P3	j��6��*s{ͪ���O�u�y�T�����UM�0(�X
�'a:��C�i�ݏ�{|����Ȓp������/	_W��/}�!l>���(�Z��-��D'@Dg�(D$��I�\��%�-h�Ӿ_|�U�v7Zy��1o��B������״}��;��"�ܴMȋ�iT�b B$�j�,�JBT�[J�A�X���B� �غ �H ��`@)B�6(��3o��4��4 �	�kL�c�O��g���8�0��s�Ͱ�~i������w1lw��t-����@��m�$�9���M<|囯5��۫W?6�~�j���K���U��n�O!�-�dYfhI�r��-E��	I,^.9!oq�y
��0n�u����3�4�c��ͣ�-bܘ�#��a�K�J��J�S���$�U�ng9��޳�R_T�9�h�EƂ�@�����OՒ�J�I9D����)㯕0��D�ߺ�<�����~������������O|�ʬ����O�ւ�Z��!�㿡e�(�)G�r�j2[���T�<s��qن�R�T;�Ψ*t���F��9��z�Z&'銢jT�4*���-���9��ւ�Y�]D@PD
�H%�&����Q�VC��H*�b�#Ka�]"�Lϰ��pF��~ʀ(
�y�&��M��7s���Y���t��1�� ~!����g_�t�3�C ¸�Ї��43�3���/�ٳ=��
WWeh���u0����#��̀�rP@b-}�j%A���BH�L@mX����D���Iָ���Z�X�K���jZ����1�}��p�b��`@IJ�A��AT0� Ί�2f�vD���q����Q��0E�t�c���
����v���}����;�y�%��j`���A����o��I_�"��>z=ݾ��*�E�'E��Z�5D8���h�C��	�@��|DIGS� H.ȹ@0�	ДQ�#�t � C���05���uw��"_? �&[T$K||�7�ӄ@������u�{��KoΏ9\����%/D��=����f_tN��;EJ�֛R7J_#�@uF)�e��{�O�����~����~�w~�w�����V���u��o��|���W�|��K�H���"G�L�2�lJ�%ͫn��1F��Ϊ
��w�yL��M����E)��z�ž6^O�:��׾�aU �Z"@�lB��;��,O�@����z!�$(J��ށ ���l���p0R�Ť���3bQ\L��-�����A� ��RB�v������5���������3S��8��"z�oso!�o�?�O?���q(1��%��f�tv"�w��T�Բk�a � J�s�a�q���	L#�iF�G�M3�:Z2r���<�������}��ʟ���G�q���D��2LE��FG�b�c`��B���L��	, )�M��`bb��Y��I ��H�tr��7�>½�
�����_R�U�Fji����P��
U"����V!�K��R]
E� n�b#��:�Ah�t�����p!P �����^������ 8>y��h
n�S� xh+�Q
�60C�~a�.�J�s�JB��g�o��}�f�g��]4b��� )�����/�9^
�Hy@�!��H�q���7��oW�߂r|]U^*%_�f�P�W�Vb�%��@�y�e>"�(ǣy���-e���'@b��%c:� D�4�e����!�@nn��gL9B9X)Z) ��oN��%�T��G�ÛR&��!��Xe�$��nғ�A+��.R�m�e���Ξ-�K��%�i3 c)lT�D@��H��)�''�o.����nz���O��#���a_+|���f-�a�0o����5_)�R�Ũ'�H-+SA˃T]�oQ�a���g�8M�X�jU�X�6ֹ-���s��2�kѩ
Z)�wR��G�؅["D�Ь(�0A� 6A�(g(B��g��#B�dU*`Q����)^C�
�hA��43��A�!��A�^�^"���{�BxF����D�%����ox� �q����ՌF��� r�0��N����N3�W��z���y `_��"����.
D>����d�"ø9��IidC�qP�AJ� �1�C��n�	1��R؍X�S�4A ��(TsE��*7�\5s���C��L꒮oZP�7�7T�/IAbJ]�i*UΩ�Y�(DETUE��Q��q��THJ	�E��,Y@9�EU���PJ�&*��"���T�\��-�˂�-Ƃq,�~�_�9�B�R����٫Z��*���l��r�^�3=��C�<�������`�hH�޽P�E�#��HyՇy��\i�;���9�ΐ־Y�'ת
J� �(%[-�<��#��M	�fS�R ()4%d�ӌ4O��0#猔R�P#�b�R��0����f�� sg8툩9�M�5[���Kύ& ���K�{}��$ԭ����ԍ�ƪ��ηváv�_=]��p�b� �d�I�oU%��w�VDE�n��2��ܼ�i\����zV��*�ӻ�'{�q�M���/i�sH�G(gh��V�V2���>���@��L�QSƴl�N�t^~��۷}JQ{]/1��Q�&�v���^N� ���M^[�f��FR�`l8��#v�E�2CHl�Q��I�d���I�zp�`��DDe	 &&��Tn��u�b@s���\KE2�L��  03�Ja$#��� V�P�C��8&���(4�(QS&��L���U���(I��+���� ����k����v
�<;��T�i�����a���2���(��r�BsR��H�L��HDL̡*_��i`Bd!��͆i�/]1^}i
�U�K��q�u�V�����û��|Խ�6L+MD$���Ｔ}L_՚����R/n�7o+%Y6qVe) e0���([�DDC9BDTPP�([P�P	[`���P���VG��"�%�HI��R��Ǵ���V�!T�T�c֜7�������Z�̌�{5Z�v<UHUI�����V��b��*K� RX�0����b^}�P�*��g��S�Ħ�i�q	e>�oQ��d�Ϥ-�Rl��������
���cJ8���%��ْ�b b4�:M{H� �S�-iM�@cS���YS���3=]<4e�L��&��7��D]Q�2<f-��w�n.�~��G5�,"�mb%S� ����Cx5���k���n��4r�x��O��Z����~��C\~��雟�m�������'PI֛Xg@��=��F"�j��V��w~" O��~M��S4����z�}�,���歯�f͆��ڇ�d��fc5/{TƆ��BϬPeX�2��Q�D��p���� +#h@�!����!?E. �ƂѕD���huRTC��� �"�z��`G�� ��o�����Z�&�Qz�w��y��CUf�<eL���O�xrTd,�X2B����$b�:
�xf�<�3{�D*}K1�ĀAB���0!h��̀a�������D!�����жt����M޻��o�[}����F�,��'����ͻć��ď*A���Rt�-^V��$��%b�p��[HA<a�`� ���tܢ�K��щ�P��-!l*1AF��lbM����l�=Y���
{?�x�=Y��k�
h1o��Ĭυ4�C(�"E���T{OT�ԩf])tj��u{#I���|����) �֬�~��j��|D"R��<�8���8D���M�l"B$��ʼ� ��7S�(�i>�϶լ^�n�ﲹ�l]���{��*���F��* �:�et�볰<+2O�b芚���ĕ(�Q	Py���P��}������ȳ�O��)<x�[�aǇV��~����@���4���n��*�
��5Ͻy�B���4��*���{����z73׍ghq������K������������E1[���
2�P��  ���
��b,�F:� E�Rz�A+0p(��\`��y
(]Yk5����C#��jV��!�׃V�q���#�g*w�ξ(�/pW�j���1�$I @�3n�7�`�@����D�;WDP�@T0�	%[�b)&l+8�b76RT�	��U�h�\�	~'��}����N�25�6��~��	Z�"�	"]��l�
�{��)T��!@��t��i��#Xf��`�
@cy��4@C��-hs�v�n�p�{_�U=4�¼(��8�2�M�[S�XN?�m�(s�5	x.�5>�3��j�I�z�K���O�,=f�{���'��=@5�\�]q�P�#����JNV]R�0��V�V�3BP�t�����^_B&3��R�t ������ߢ��h��t%��2�O����T��^/�k �Tma��0�����?{�J�KM�CϷ��r�若�E�� ������������'���{�	�|�Sx��oy�g���R��޾�gሇ�UM���K:��G�̖"�f�Ve^�~	��!7�l�n[��%�ӂ�-J����ן�)z�+��O7�J�wLZ{Rj���5�X���ʜ �2�H
��N
S�\@�M�Aњ�7Ȥ"(�}ge5�t�@��r�1�A��`�8T��湒V:��}�*�%j�ΐ�E���m�"H���:��`�ύjڽ���D[̀�� �#O�,RD�l1gV�@��5r.�sF))���!R�e�0�-."a`���UjhדX�3���=(*x>V���-LY��u�� ��=�u4� pT&�NвM7
SX��0���vL3(O�<�'j���J�TD  <��:o �%�`�ov ���^rZ�U��Ր�5-mMZ�ЪL�p��Mq��g�n��[Bz��֥��m�h͏��_H}F�Xy�-��׽�O�}��)��a��$	��L77fP��
�����mă�s��2w�v�n��Q&���	6�U�!��o�N�Jj�u5��]�r���5[��ht�ʘj\���AlD���^�Q�2�~�*��~`�L3�j�Q���`���69W`{��$
�����O�G�+����`��e|X�S�
���ޔ|�'$�T�<hIF�kF��PG��r�V�V�̓v.+ֶ�Im���'V���wS�k�ܳ[�u�z�<��/[�]ey�)��ԪI�l���w&�v�@m��d0g(�*��%����6�%P�Q����4`�r�$3����л���ٵ��^&*�W�*ШUi��P�,lM�����Oj��w��(W�kJc�͆ ���Cf�"(U�81B��� �\��{�V0P�Zl��-×a��|Ļ���u��
H��O��T�C��]�rQ�͋�=����v��(��b�.�`���.��9�ƺrD��L��Ϫ	(
� �	�� %�����T "0,��T�2�)��!� V�._�� ���M�	b��GX6�+��:ٻ��5m�*��Z7�6���S�|��β(������h�Z={ċqQ=z�RKK�2��,Dl}�I��,N���9�!0(0r��b��#f�-V"I���`I��7�f���ۍ�<�?`:$�3dN����z��
�:٫��{�����5��x�M�wơ1w"+�[��`�G�����\�3���}4̌��OU�#֌�z�a	J�������9=���G���'�����q��gq�!m@�S�7��T���%����%�XӒ�e��l-=�]����+���f�����j��$��Ic�٬R:�컀&+D�F�¼��,����*�C5Fd@i�DA����2�b�'�f5+�Փ-( R$�FիoP��(2�5��Q��/#c/��2n�G�A���vo����Rf�;2\@� ���l�r�@�Ӣś����O�\ʲ2wj���k=1�B�l@R0b�u��	9<�f(P�le�2Z�p$F(&���d����Lur�Ֆ�R��
�12�����x0(X'�&�-���.���[����J	P�o�Jm�tU�띪�ꋵQz��-g�R�N_Dd���	:�V#���Wg��
��`L�,IrU�TD���*
���n!�-�b��PF 5�����B���O#�-�e	^�@lFT���<'�6N�5׵Z�ֈ��贌����3�L�Z�ZmHͣ�&�+����o�
o��vT((�e!OG�)a�8B�`�7�W�����O�<��֔��|�s�LG��"6q�V�K����YyY�nJ����^��:��*p���T���85�~�4�3�<�ET_������J *5�*˥�v3���k�$9�/!��O����ç�K/�>T
}z�H��'�|�Ki>|���:!�)	��lJڒF�4�Tzh���Bk1�"[�R��tE�uO��V+�����oS�M6,}�[}d}��x��
��!PH=�k%�����(��`�)�X��>6�	!��MHP��D	3� �z�,G� ݮ����,c�f-�|q�5�u*���m�cB��5���+/H� �������Ѽ��x-$R�9�T���9�Br�� 8��ԗ	`A���
)3�
���2z��@�R���RlT-�R0� S��`?r��y�]>�k���ݵߴ=q�e6�Z���<�~��{j��mˡV���Ȧ�+���6*����D���̥� %�L�3�c�j�V��?GS�f`�	 {!*��C@k¤�A��^I2&��0)jߘ�%le�w2�K�C<�<볳ؿ���[;�K<[����V���.��*!��m+��Y0�*aD
D[WHE)���h��!"�3?~�9M�\I�a`!������./���/DH�1����iF�%3�焠-n^�U(��Da��O7_Ջ���׶6'������ڴ��pL��idJ��.o��oK�]�����M��`�Ř��>��9zB� ��o�7_��v����[��/�>����Q誊��/!�Ã��͟+����<�J2�\l�o+�`�D¢Z�E� 5~��$�d�F�-�k�}+v]�D7VX2�W^�J�T����i{�	�槣�!U2�bk��Z'��`�[v��kw�~�%2� n�>�{�8ҌIf$(PM�#�f0pD�4� &�����܎$t��Q^)iՓ�5������Z�t�i�a=�R�P.��	�2$)����<!���JѶ��1FcD@�hID)�T��"P��{�Rޥ*-�K�=�z������(�^�VN��BJ�F�<�u��'5�AD�O���[�q[y{FEP������PB������ws�fԁ��B$���0K56YH� P��8��1�8�ᵕAB�~i��s^���^'���w��DO�ZU��_�.��B^����!��?tf�����0*~=DJ%�>���Ŝ��[�yBN	77Oq�&�֫���k��/�q��BDPR��`���'����'8�(s��4M� ��j�����@M�yW������BS��o���3�(���Bn����\������nșaѪs �_Z��%�ތ\�1�������O��;�����]|v�o5�&|(����������9������<�ђ[R�1b��%�Y\1KY-~�g�7ũ?���@��y��Q�%�ף�(zvh���3!��n�;�@�����7b�線�F���J�Lv�"@z�0{�v@Ĕe��$�P�g5�V"w(3&9b�	%�`W�}��j�����#@JFN�QJ�`��P��r �լ����h�"�(�F�׷�>k��F��Z%�2 �)f��~5\��@�i&���y�R�#�1 F�u����"�!�keA�sQ�T�Ů?FFL� �ϧ�q'˵�H盡��]��8`�ce���4�e��1&K�9��
϶΀e��ʘ��a�:im�|ʼP�T��R7��{U�x ��h� T�ʆ�5T�/D@f�<IP	�o�������c)��%~�i�n�/K��C��nG�V`(j������k�gM�=�S���I�Z:o�v�TK�<"BQ��������equ��d�>}�y*H�#R�8�v�ǓgO��l0������)%��<�\
�	����Gf��%l���7u�,,�%�ô$�َ'9K�@�r����:�җ�3Q��6�h5Z�:;-����)z�LY�u�2]�r=� ��2�������Q��|y���ǃ�+>,����"����]|�o��S����<}ea6��՚��I
�-~���Xr1�doz~d�z���������j-a�3�W��X��L�L��1*#��e���5_]p��aM�5�A{G&�L`����Q2a�#2f�Z
 B�� ;$��5�02�x��F��x����0F�U����W��r�%	���,KZ�v���߮�sk�c	�F�.��j��S�-	�Z7S��pn}�T�JAI�s.AB�H� �(IPf+�4`�ڎA�%F����m��J�5o�HWR��{�'�����e�`�t��S^�g���JʟP��fL'��d��`��ք�Z��e��["�P5LXZ�F��s�X�n{E������9ke+��u�v�1��Q^+�sZ:A��.9�gJ�mW��E�����]��wj���/	5����p���J�Q����R�tx�iNl//��G^�~������ FJO�1��r��a�ʌ�xDJ	Zex�)�sO}���a]���㥯�k�;"��Ȩ��\^c��V��$����z�S�W����I�z�^#3$��6B���?���/������}��O��cߌ>p��������7�v�돤��?U���J:�%�D!ɐ�{2��R��s��r�~��K&o#�j�2 �z-6Ӕ���9x�ڼ�x�h���z�,����|�r-be(b����q,��2n�P��0}��S��j�6���%aFƬ3�L�2c���l�!�pG�C�ц�l ��xF�R���,�z!��OX])t�$����x�,�{_�V��1w�J�
��� �1a@ҌP
B�Z��X )c.Y3rJ��>�gD�F���E)+R*`hQ�ڞ�4�*������S_���5��[h�y��������0+����e"��Q�EiA��iz�7&2Mlg�$��0��T#+t���Ĭ-�ь 5�Ό.!K�5�l�n.�����ڪ�_)�x�ٛAsj ��v��
���F��I�7���W�S_��("]�o���9\Փ�����QE�d�C q@*�<g�R.8'l6#�FpQ�qy}��|�u���x�����}�� �i�8L38D[����	i^�,����3��s���Qp�F��$c���oxnI���J�\�{j5�:+��8n=1L�����\�e ��L	N��
I>�����0=}��}o���x�o��T���%���ax���(��G�|T&�Z��6�	4Z��K?�Lړ��k��S�Qd�� K���Xka���Xv�2?��Kq��/8��V�t��=ʿ%C�6��"F���������ѫޓ�:oAT�X�M��Fւ$3�L]�[�j��z�bε�e�vW���8>@���:C9#�Yp�����S6���εRWt��}�L��n��lb1�w `�)،f�
��֖��c{(KY�KR��X�%�eA��`�C�hQxUkKlԟ�n�?m��
��;Վr���G-�g�hԽ�h�*���! %,^��>FcQ�GҌ[��5-�7�޲��%���q�8�&�ڡ�@�Pڹm
�Ң���[(Gc+Dj��T���E�:/����K�����װ��Y{R�H���3��(��#pzx{�W���2o�C7ԛ���3*�[�@ss@�qq�4g\]]���#���8N3�d#T_{�%�~�d)x��cd���T0�qs{���{�a
��rFN�ĠYd��lRks��t���8Y�;����K���:�������H#���ۺ�I�Z���~���B[�f	�"��A(vn�:m?rI b��t�^��/��>���;�>��ۿ|`
]U������_���{~����h>��2A$�g#����	�j<]!@� �Z��&&�-�D;�5i:��d�V�D�P������e��k���y�H�b:������;�[Љ
;�Ӈ:�KA1��0b[�Q��)����ژT�@�2*�n�aP����lY�(�R$HP䈩�"˄P�B	�C�Ad��$A�%=����!�xe�j�!<d�Bt���&a�1)���u��{+���E��qq���ŦTJ�BEj��"�pE�����焒	4bX:X��Ա�@$BΊTj�
� I	b`��`?�΄cV0�d=�j��P�h�0�e:��I��v% +ͣ�̖��R
��.���?ۗllPh	�U�	`LK)(Z :!ȡ6	1!�4����$"����JMk_]�F&k-j]�
��l����������4�����	����E�֑ �)YIT��ֹ'���ւ����v�m[v�,�Ѣc"]�-L�:�gevF~�>5�n�Y��+;��i�����w�l/����ݣ+l6�4�����f��^������	�b��<���,'�x8����r�m�{5M���#'
�}y���vΔ�q����L���g'���t9 �o�u]����C뫯'��Z~�U�؜�j�$��I~�������������߂����|�o�-�������=���I���t� 5���,Ѥ��-q2B�Y�u�A��ن�W]j��.�`��O(������W5��w�Z���|�$윾�Y��\� ���7}A���[�U-.W։)�M�b���,����f9X'�b���-CY��?:���@��:C���L��E��������� $�Z�o����,ٺ
�nNUa��ߝ%�����D�c�E���m$"d�q��fQ2�T�p HY�&�D"D��`���5z*�\�X7-����o=S<>�K대dzZ�*ζ:XNH�ԖF��=��c��Z9���a��\�Jw�)Ag��^"E! J1_�,fK����rWB����Lw��(�Evk76Hm?��[	(��a����e�`�|v�������a�Ӄ�&�E�5�Q��f��J. �}�j� h�H�S�f8�Q��q����z�-sga�Z�jkKZR��i\ (6�t6`ETPJF�'����#����a�-B���RJ��v��	2�9c�#a�ݠd`;��n�SB��)8��)M�P%�J�!�,,sKe��{�x>I�<Y�;G�����z���c��3���Fw�c/_���>
����:�	l���a.�24-�D"�%A�d��_���y�}+�>�<.}>0�>=~��똏��W��GJ:��Ɇ���#���T�]J��Z��5�^��K�.ٱ���ߟv�[���`
y�1�f�)�=v}rg_��(],����p
�u� m�.�bD`
��jrגd�(�H�ſ�P���EfZj�U�u���Z�EY��U�	a�#�	*���H�,�ea������DKM�Z���0Е!Ж��0�H(�\=j�GV@R��j�s�&��J�zܘ�$"g˼�LP@����Aр���@V�����L���18��ߺ�qCN�����CS>��;���@Kz����q��ǵ�U ���mF�V�3C�2їw_�Gv^�a}�hM;��Ty���"���d"Y�Bɦ���-=y���=�P��� ��"+O�5�i}�W�\=c�)�O�w�V���*I֝�t�m?\��f1�g��i��[_��&@5A���^�j� ˄i>b�#�`�MeZ.���߁����A�f3"��'X�RPJ�dWǨRs�Ob�f��f��}u�V�ק�)�ޟ��q�峽�����Ým��xr�r"_t]]�Ƽ
 *���=.�2�1���O�g���?|�����	�������UzH4g�o�B��$�w�:9M{)Z������dP9��E���U��Xj?������[��7�*rfMU���ݤ����sZ�Z2%���0%�Ɇ���&�B7Nl���i$��5��דs��SR˜O��:#�D��#����<�;ͳ5��d�&�N�������`j�nBAd�z��^/�s�B*�lXw[k�o����[���L�o�m��a� �%�Υ�Bd����T���U��CR׮������x��w��?���Q�]� �����s��vJe�X������֙��������J�+b�!��i��[+�:e��#v-���K^Rm���/�ql�^�:U�
ъ�4/{CZ��v����7BNAulks�AK|v	�-�	�>9�X��*��_���-�R\
3n��|#����)��A�@ ������vLs�������^sr��@���%��n�#�<M�ӌ� ��<�w��u��{KM}ϟ�����-���'��:z�*���V�ja=TÔ5�Xȥ�L�Kӌ m��@Hy�.�����|��o���>�m��'�s5�Z��+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs����|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�f:���E�s�.�L����)������@��w��{n�<��D�^K6�md�c�pcs��yN���I]�$�����i�!�����9�x��=���b��ko@�[��E�S��y�a1�F�bf���W|��	�64졻V�#���޵_���d���є\[���0�h��9N�	���N�!�2�}���2c��?�ߝ��
���{��HI��z$��W}����7S��o=�|ֶ�����]b4�3R. f$ʠ̠\@egJ��%�Ȼ=�T�4�h��]�8T7�1�j�{ȷ#�i���f^���=�d�w=ܲ
	�1Hg�|_��O�Zb#��cE-cm����>AXj��T M�Z�iF��3ي{o�GE�z�E�8c�v�7�n�6��e��I-����#qs��F{J��w`f,�y+ �׽S��=Ӵ���Í�����WV��H7h�!�kO��6վT�#��N�l�N�E��O�2��e9~-�����!�xS�U�׾�19��?W��NH�w�ȥ�"��x{a�p����Zĺn���|r�j������!,}��}cu��o�2�T�6�;�n���1tKY�&�!{��1��]�}zߺ�F��t�*���ER;�H�t����ǯ����z��d�a��x��iW��Hcx��-`�*c�&�b�ns�z$�o�g�{/E$\#>����ЅQ��HIM����+$'�4AZ2O~� ��yM]#�ߌxn���%���L�ځ��ہ�̣��c @�b^�l��1.��cch��}=��&4��ƒD+oB�#��G=t�b��O�Jid�m������>uʫ��C��i�&�T+n%+n圁��){4���g�$��J��kB����ͥ��V�ƃ;�:�J]]w��{�X�?�:�&���=��������O�m�j���*V�����*C�=,�!���*č{��UD��������ݣ��q�=M�\���58.ɚw�iY{���tG����U�-��~���7�O�o~�e���� �il0�C��Ъ��m-r�� {�sB*;P�~�S���� ����x��:П}�{���9 ���r~+��H�X��ԭ4���}�o�@j�#]�^�*$ [KR+�#��W���s�Ƭqtݱ��m�|�6�]�ݲ$�|zYh[=�=��{zQ���f`�{CX��]cX=
�եz�e��i* 5�¾Ag"$����LDA}L����vA��!�Vo��t�2vۤ�o����j���ĭ>�s�����Jk��\,fqO:5+�Y@�����`�083L��&1���e0+r��guU(ߚ=�/��N(d1���WG�1!� �wX��̽���z�ͷ�kߓ�XQ�d�:x����I�H#W޽Y#)���:M̢���t�܈+�$K�d�f�]��D&I^�h9��� M٢>�w-���ugQ��������[�˼`�ŵ��ͫ��}{{���F?n����%��m�4����>��	�s귕��WHպt K���S����TPe��Ċ�#�ہ�Z3!g��tlW}k�Մ,�c��xh^Dp��Hy�Ϙ�)\ER-Z'	@�>Q�ڣ5↳�BU��?��7�������a����^{3D��m#�2ڂ\�������$"�w��;��9�8A�
��r��\ (�N`ڻQ[@y��Ȼ?��?�7�����?�7Ձ �����_�9,K��n�JOr��ip��0���P��NԚ�x!ء�:*K{���G�������c����_���pc����YĲ	k�Yi�L��M�0i�>�O7�77������ɼ,�l{H�7�Q�L�F&��5ܷ�R��0�> �c}����5�%��� 6���m8�/�Nv�j�$~	��A]<a�:s#\WEU=������hJ��-R��y�x>�Ɋ���p�4N���*�f�kǆ��q�'�:G˩E⑏��5�QJ��E��k;������0<�/tv�ֲ�"�PuHޓ��i�l�����'���f�71�:�^��)!!�Y�F�i��^��̮�X.���R�.��*VX^�6�Zl�^X��t�Ϭ�$C}r�n�I-��g�����]��^�W����X�����ӫ\k`�f
p̌R\��>�4�h�v�UR��5ۏjkX*0�Z{V6�͕dG� �_�{���P�u9�I��E���5r3��#�Q���-b7�"]���=j�Q�d��^6��SF*djp�<d�X�4y�������t����w�Agq�����~��K���7~���NzE~�HY���h2�7���rZ=��a�]�o�2�����,k���m�cV9�߬�'76Y�hm.pϫ��Pݶ*�o`�y>���r��e%�y�͐t%� �V�:B�6�I|��9#�y���@N	3^T}x��i; ų�ÓD����5�{�!�l��彘,�^$�)2Ī�uV�M�M� r[<�A�J��`��ŕK������J������@�N	�^��
4��Sww��3�^[/���ӄ=�8��I���Z�:�����������>+�X�����:�^�u[���՝t�+�48�b�/��	>�N���SO�)�&9�5�~h+e0'��m��R�C1��ٌͨ0���z��A��g�y��������@"t��q���z�7�\\��Ū��Vḧ́�ך�_l{�=�$�ު���j\�J���r7������f`8@�V�	)OÐ�V��d3�ن�����u]�P<m)^i,zlp]��v��{Iלޮ�n�l��gA�m+���Kߺt��"������ϻ<��2��	x% R�(�<�ly#�I=�)!BJ�א��s����2�^���A��xS� P���o{���?��~�����|K%��M~W�̓���0��F�Эƞ�j��e{�����@�l��l����]e<�}'H.[�19{xh�gW�z_���
�0�y1��؄�Z�W�ZG����f.���X7��X3#b҂ H�$s�x�i&{���3k��!^?K�ٔi��@���u���:�6a��#^6�x[�sU y�V`n ��y�P������h��=�f���\�b���m��	˲@!�rBNdS����̣*��|�K��]$�W�����f׍y�z�c�S&�������خ_���[���ӱ��f=�����}� aW��e1/�<$��{�잒��!�Ecm�׾�\���@+�2��<	��$���,�v_�쨧��K�6�MX�/����ֵ�][�_;����@�/k�}���~��x�ǟ��vcٌ�_����o�=K e��6�~Y��� MpCI��n͢�Sbp���^Y,(@"F���ڈ��LP�H �)��M�3�،G�{(6?\1�q[�G�H��U�p��9ҿ�h�����8�8��=j�w����!�c��E� W��8O�#�8'(gP��T�<�R�0=��~2��+ǫ{�=���Q�y����~��﨟�9�����Ͽ��?�����"G4,X����C���IA ��۵J�ԇ���R�^/���O�6w��鮘�mB�:�D-�	�.�V>�sQ�Jzh+���R�2]�!�ILloߋglZP?_��IU��b��EO*�����t �4r��mU�g�{}�ȉ�h۞���?��26�5f�!Cү
�MR�Q�Rd�3��n��{���K2V�,��V\^6<)�L��Vۨ�ruh�S �U�d�3 ���խg�!e3D̨i,:��յ���޻�cܧ�g���ՙ��z�F�9��SztC��9z����~���M�A ͞̳�1r�������WkU�|4e@���zw�}-[�;�-���}
��]�2�Ț 9����ģX�0���y�\�|���q�����#i��n?-g��=6�k=��n�z��X��kU���4��"�%'L�	9%;�`�L
挤�T9	@�l�Fk�4r��CY��
z���M�B܈�\�H٣~�������zQ�p��������7�����zU�Yn����n���zU���{�*m�ל���@��(Д�����7�\��mJ{ ����ɟh��}���aqޤ�it"�~����Ư��q�����OO	��1�H��֦�^A����e�B�aH����#T�k�]M���C�7��ƚ�G��.[WF�yzŪ=�ݳ{�_�(Z��Z�V��Y�_���'Q�VJ�D��Z����3�0��t�6v�����"����)ﯕ֜��ٕ�n�9n����X�g�W�ۡ�s�.w+�:Q�M��s���e��+\���-S�n�qy!x��@� R=�n��j/SL)#1#�Aa�2RS�g��L4[;���抔3���L�\@<�6����h��q2���zR�b���M�j�7����Gd���{�CZe�EٚK6.b�֘�(2sF��BW[ߍ�
2�L�T��y���!����sF+tqt�.��y��@/�Z��wz�Q<�]O���zM����Y@���U6��d�{�Q�p��l�x3 s:o�!o����{�Z��li��~�4M`2�k��b�dbO�JV1�'�ͧ�l�*���*cؑ�v9EWEi���O���Q5�e��`|@�����ݯ�*�D7��X�vO��,cF�f�z=Ł�ߏܻ/w.�^�z:]�L}w6c���{p��yO{����0s��e������ `�(~���ެ�it CB�s�(�|]./~��<x����0��ݽ�q�k7�M!��湨����z��u������X���æ�lv�&44���%��t�9��#��4<�ѿO�屛��L�������y�Խi �40��v��`$O(��K��;�m�%v��IM>��=3*(�9�++	�������ٟ{� �:Q�W�JU���QEէn	�������Z�
hJ�1-G\��oy�Ɗ��ZQ[C�L���PB.�zf��y����&X��V@����ē`i���PJ��eƝ�~���W��&�9�f�mk�p�)*�zlN{t	MҪ7��w�Ev������aHٌoej���v;�a�r�l:�P�6��&���N;H���A@*;�i�@��'s�tq	=��.�8����Ji�n��a3�'7�ӣo�`$�\9��#���l���#2�kH�+���p�ѝ��Þ+��I�^���}�Wd��[=���m���b��n����N>��B�x��-��V/n�����G�9m���\�\zAl�
jd����å�>i�H�!��G��,����U~�������H�)Rqs�~�	�ŏk�EG�f��;@��kDJ��C��Ɣ����2퐦�T&�r���i�������S�����7���M�M}�w����s�(>����������K*�	Q����˧���9���e�ՕP��=r`�ʔ,TBCAZ�^�Yվ S?�W�����z�h-�R�ԳC
O���Gچ�\�]�F�����Ⱦ �(�a��B��@�)���j���[�	9�0Q�!gܚv��.pQ�8�=&-��9!��vJ�>'�Z��ۃ��d�ѣ��MW�z���am�{# *r�P�̌&�|D�'���l��{��	g���A����V.�Z��ǓU�i��3�
�Q���a���	mO(��e^���b��dnD*NMq���'2���t+cAc=�t1��}3|��^�E���t�Ve�*���E�x��;��}^wJ}F��NH��9���=\��&{b��кN�y<�i�`KM`�ВВ��!*�߃�'!w��g0JbdΞN�ϚR�y�<��7d��(�ի����U�&��[����Nڣ?�Ag uY0��=?SA��K��郡l*[�N�
�� M7��6�<��#�,H�L�`ڡ���&�,�V�'IR�tEj{��p<][$*O�i�z��CS,�tid�r;��?�z�9���"M�������[Ov�)�S�Z��E�v��6y�.��3aҸX#�}��+Fl_�}��
'���#�����-��:X��D�+�?��2A��\,���`���:�>ޖk��G����S�7�o��C�3�0n������^~��9ܯi��+𣤺K������|�%՞�@nM{ۅ􇗺����V����V�@�W��X���K��m����xo9a��Dmآ�E���ƿ�W;���	9��5�o]�@2#%�BJ�����[�`���T�����3i�e������%v(v%SvO P����=����U��>%�BA���H�_o�̬Tv�DBDJ�oӴS����'䴳��4�ݑ[���Z��¢�V�dJzJl=����`�k(�C��&�s<����&03��Ќ�)�J.���-|�Kh�Q���D6��� �	�+�d��'2�'�����б�������Ƴ�j����ѾǤ;����/xލa߽)����?�+T��n#]6�\lP���*H:���(B"�5���R&P�x�M�4�����m*����S�˧�r@&'�V��o&���5ZU��`���Ƭ AM�A�H9�%e&eb]�E[�*M�*n����������N|�����M�D���'�UIDIUHd�Jċܴ��}��.��0�X�R�)_�̱��� ��?y;��3)Ӕ��_@�p�X�()�	cވ�Z_����dެx�@�!���RaKM�}��M$��IU��u5�!d�(�5�;F��(���F��7������7�S'=`�=#��h��SA�%���r�;�:��ns�3���j�������\��|Ͽ�����?1�2: ����_�ٟ��˸������{�=��$���酪���k��+���q�����f�KI���ja\/"���zC8b�=4z��r{@������G����xiKtE'�zPTm85A�#�d�c����>)I�"��gMH�(^�iyfFJJ9`��\pk���t�|�|@!k� '$0)Zv�>�����������S#JU�-��DG"����> ½�t���!�'�{<pՓ�^K[qF������
9��*�*�T�lҞiwU���v��}-�:�'ngpR�Xt�@p�GiIN��2��e�t\x8N[D��v�D�����E#B*��pk���-­���.����yL��X r��k�ivD�2���MWA���vf����^�E���Y�U@�!��. d*����
��Ҿ��4%�\4��!�"������3v���O@�L��K��'�O�佧��̤��&�ĩ1s#BUEm�.�<SJs���r:��� >NJ�>щ���隠G �rﵓ��"h'-j�,`���W��(���p��C�])�n�����>�|	�U=�&��-mr)��փjۋ�I[+R[��L��$���"�T��HZPX�XG�\���).��)��@�KL��Φ�ժh�J��Ac�>TB����H��nl,��&P����=� �
�V�Aɮ��;�ױH����}���I5��u�g���)#�؝��*S�g���X�H��{��}�E)�K��7��v~��,�Q���w�9���G?���
~���=�f��˷ԁ ������+��q���_hy����m���<1��k�/Q�"%ki�&Hb�0i�N�:���*&X�ܛ��x=��hxI8������V7�U�C&`l �U`Q�PSA&��V�'�W ~�0)R�P�ȔL�L2�0�f1QA��r��i�;�ܙ�`���<!���VA[`�ښ��Y����T���<�Ӄ������5f�� }�2^d�<����h͉+���ݾ*s��n���ҔX.�����2��r��Sʍ�y.Rk���&�eB]
8=U�߯����wcW���������T�E�ITx�j���P�'n)�4/x���Ǚ�JΦ���	9eH3)K&����S�>+n���pkG�mFW"D���+����}��6̨��m�.o�J]ꛣ�^�lm�Ex���~��Z�.���. �Z�����	uf�(�H�V��݄S�q:	��)���gԚ���%��ٕJ�n/|�����S��#_3�Cb<,�����_�į xE��,*ߨN/��[.��[ޕ�)7�,�rc��D¹4"m��kd�e�&Mx7)�De�k�,�jEz�Qr��m�@��r}dL�y*iJ�K�Xu�mn	@Zj˵�,�%�9Km���V淋���R���|�H}mym~B��Vkˡ-ׅuIB�mAʌ�����q��i�����B�N��]ɸ�`\��КE2
d)�vB����hb:]��HPP]Еۈ H��u�Ż+]�����dE�"����Q�;��'�#u�BDS�;oM�{爌Z�q&�a>�@0{�>���>xe�R�#O{�2]q�-�������������R�9�-x�v���Ox���_�{��Oѯ�ҿ���A^�E�� -&�)&<Cb櫶il��R����D��dZ��\���lz�{��f����!���&N��@2AQA3�넂v���z�����+de
��M�1MH�=�N9{�3�JW�c���].pw�w����z*C9!��Ҥ�,Dt��&ί���Μ��S�\N�O	��*��9O'N��ʇ%]ޞ?�3?]�|��r��R3���֟Ih�J���n(������-���Vlr�js�L��'���������9\\�5��Y�q}��YQ�KD�[k���i>��c��[A*Y/��P8=��J��e��yλ]�23@���5��ä�ĉh_wD�/3������?����²]KοNە�9���D�`P���F�1Е�[�pV(�GE�B��:V��� �MՆt:i�_B�	����Δ���K�Zv;�ۇ��R�I��x�s�j��P%���y��SO�r��xI�o�i�Uʻ_W�/���
PK�%���VJie�qj<q�����7e��[,�"��y+��v��	�fc�T2���tЗ#�X��'kgj3P��5�S�L�z���Pv�L��Ί4�EZ�5H���P����"�a������u��Xj�3Z�2�_��m^^���h�۲�g��nk�����T��z(:CeA[ԥ�-���e9��#)���.�*{Bk��:5��m� ���־�D6��SS��' $Ӽ��l�J�#��vng�k)��0A��}��1 h����n<EYi7587"<%��Z,�;��R��xJ;K#��W����^*��J���.>��[�����-w��K���>���4�˸n����?$*���/u~{�si���fH�!��0���n۵b-�=�
�<�����L7��^ �ʱb���߱�l	�W�pya��������+�
����`E6jU��.�֐S�R2�2!sƄl����1+ Ta�
�|�C����%����gO�6����v�2	8w�_Ki����/�gSΟL)����IR�s޵��V=<�T��'>����z[3CiBK�' �g�y�o�z��W�
 �ZѤbYf���=�����^�ƽ|��5?|�Wi̜H[�Z+��L�-;�tGTo�����E�u߄wJ�������rI�3Cs��I�LXTY]S��'��Ki��T�%����z,,`�jR�["�*-��GA��L{�`�-�z/�C�T�R��fPv�RR�uG�}k=�ѓ�Px�&�U�[U�U����Y��ki���R[b�K[�R�)�:/u��~��ݾ�P3�ք_���|Yr������?�z�g����4?q[�p!�ť�|K ��}�SH�ۨ8y����l5����5���?���x~���  �IK���eF���!��m/����y��Nz���г�������;�����<�xWP��@��Y󤏧X�+d�RL�XeW��Rk*��tD=^��%��i����������R���f7�Y�t���A�0N��st���6C��P<r�3�X�\� `��X���/�6ʀ���ƞ���P&Fd��N6��],���H��i�������N����������Oķ� ���G��w��~	iaҧ����.˿�d����&�TZ;B<N*�y7��f�M���G�X��+?Yŧƞ]�.�^A�!�⣴�͏Tتe��ײ�ի������z}�Wu����
h"̲`>��Dؗɫ��r�dNإ	S*&/��g�j�(�w8L�qQ.q�p�������S�Ň��ʴ�r�ʧ	��=�_�����WN��i*{-��|���~���r�0��	���	w��^�w�RI8=8�x\p}\���}������Z�ڽ{�ݿ�w�S��,���=,�	��D��,hMH�uB�ɋM�D�o\1e��.�rb�2A�k�+Q����c�i��~�wW�ֻ���-�N��d�x޷$i�95��Ě�sK��wAV��&a�=0�o�{�M�7\!�*)TD�6�(�q�nr�n�r�ׯ<���8����^�_k�
�gk��.tw�6P��2��O��/t~�{��S�[O���3�[���ew@��HE��}�F��7z������~�+XN�X���f`>bz�I��5˼�\�$e��I�i�z�b�E}7P���4�ҔT�����j|k�C�j}�&�,G���ꅔq<U\_/&*����4pݴ��6�c�F}*�����T� �#&��Z�u��Zunqs[|C
ٍK�Q�H�����5�m��
ǽ��vS!T�^�m�ZJ�۾�T.>���.��?�����C�,���#o�R�'�[�@���/�P2�_��SU����j�ai�;[��&kaZ���R����pk5�9Ϗ�$x.�+m?��O���#޾����6�ի�{�+|���k�W���Ҁ�r�um�>�S�������*6PD�]���p�i��~qUP+ �q��;�{�$��}Wn_�zpk��������y7}\���~��_�}��اtwH�����l��t���^���Ջ#ꬸ���)�N`͠�P�x��5�EЈQ�RFk%��u�_b�9����6L��z���X��^~���p��C���ⷿ�{s�U��g>j��`��p�O?�=}j��km~?D_$�}����\?�;�F�|��x�,f8���"g�����Ԅ�i�i^��+�
���r��;>&�%&y\=�]�pm{��u-�+�P�yʜ���M�Ȥ/{�ڏ�o�~��P8%3+��J�B����bG)#s��8�\v���)���xˋ|���?5���Η>�1(	��5�O?��?�aY�����I����iE�I[��XߢV�0�}h�o�ӽ���X#U" �/���i�-��ke�"�
WU������#��W��'�bC)���QR���(�$L����!>�b`�&ȑӄ[��ؕ���jŔn#c�D	�/���~�ٯ=y��������n�����ҧ_���$4��sϾѷ4��B?�a���{
����an3Z[px�����{���%Ǉ/��J��K��Z�k���bAkC&��^�M	�
�B8͋�N'@��i3/W�Zsx�����F%\�I���+���'�9#%B���d����)���pLލB��Z�l#Y}��	 2��4ٰ�4������k9��J�WA����>���8��-��7�������@�/|�ؽ�i\��h�G�y�����^�N��wf�ߩ�h�����Ui{�Z �Td��^��G��7mܫ��#��f���a�
}������J׆������,*�#� jC|��I��WhRQ�u�K���%d6�f���i���U����\���w��;O�}�c��̻>��/}�ݓ�s����p���7�6A ��_�E �VA�3�y��镯���t�.>Ȍ�6ײ���{ҖI*�r�2� ���s�>m�P���ٔ7��@��xS����]�>�
U�b5�UKIu�����e�i�GǞ�2��qA�x��y+RE`���{ΩW��(/�r?O��r��/Q��H��r��;���/E����=�;��O���`y������SO�vz[m�gAx*ߣ��Է�ջ"� �C2IUXUX��h��d5�㒮��R���Ůq4%+a����{�}�EM`B\���� �����MLPb7MP.>�E-4�4�\�����������������O��,������e���[Z��?��O �^�����>�j~��[o� <xG=]�u��
�>��{���і;m^��T8^�Z5u����54��mmV5�&�'o
�v�k�z#�����3!�U���(q#2��ܵ!o(��p�˔�g��I�.�,̩��2_'N��k����?���?���^�� ��}��F���t~��[��?�ҳ��P��׸x�S}����[h�Ro�N"����P}Z���[*8a�������խ����c_q��
���7�.?IB�,�m��*����>�0��וf�����m���5-˂��Jɨb�1S.Z�W%O��������px�s���/�{�ٷ�-�<�����o�� �g�ԧ���x�|��� rxn�,�����6�<S8�J�U��o"z��o�N�Ts���(��yO
�jz6O���"������
�6C����ܭ-nk�$))aۤ>�i�2"��2%%NB����J�f%>�
����K�ӗ�����qY꧙���F�^|I_��R�L�Uo{���ѷﷄfw�/|�v�j5��@� /����#K]�&�h�Y[M�IRQ6�g"�邈n�-�iOL;UL
ͤH`Ndc���X��J�d�G�*T�`�FB��5���B}�+��De�8-3��#�*�2�~�'�V�J�����<����������O������/�u�4��|��ѷ"�JT�}�8�M����p��~�N��p:ͻZka���:�D�ۙ���������nI�Q�h�k�y^��T91133)"�b��f��@�Y�Z�\r΀���W��X))1	@ں�-�1QQc�
�
�3���9�gN���U��N���,���>+���S�S^��N������¯��'�
�����w?�Y�؏��}�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��1�Ӓ������   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X    IEND�B`�PK
     w�O\d��   �   /   images/a262aa33-74c4-460b-b0ad-c746896f6744.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK 
     w�O\���gm gm                  cirkitFile.jsonPK 
     w�O\                        �m jsons/PK 
     w�O\�'���d  �d               �m jsons/user_defined.jsonPK 
     w�O\                        �� images/PK 
     w�O\��;�. �. /             �� images/03bee633-62f2-4ed0-b5c1-e772de98cfcb.pngPK 
     w�O\j���  �  /             � images/85ff3ff6-223b-4d64-b6b1-3b6b2877ae4f.pngPK 
     w�O\���� � /             � images/bb2d2ee4-fa83-49b1-89fe-70727f49c778.pngPK 
     w�O\����  �  /             � images/32487380-bef1-4e4f-8e56-19d5eed1120c.pngPK 
     w�O\��=Y3  Y3  /             ö images/3d684ffe-1f74-462a-8eb5-42254bda90cd.pngPK 
     w�O\���|  |  /             i� images/6fad6c1f-1fec-41b3-8a64-12aeedea4fac.pngPK 
     w�O\tX�K�~  �~  /             2� images/80e9010a-c477-4737-bb01-43c9d75c1ab5.pngPK 
     w�O\ےtR�2  �2  /             Qz images/6a650d67-2f6f-4705-ba20-a1e007a57e5c.pngPK 
     w�O\��_oLM LM /             O� images/a65aebfd-90e6-4215-8cb5-f5692b012cc2.pngPK 
     w�O\Z���N� N� /             �� images/7e39c2f4-a1af-49ff-bc26-783004b83469.pngPK 
     w�O\�c��f  �f  /             �� images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     w�O\��EM  M  /             �a images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK 
     w�O\acO��� �� /             Ku images/90a26a0e-dc54-4725-bfe3-cfd4e64c35ea.pngPK 
     w�O\4	sj�i  �i  /             JD# images/5c3bf32d-6880-4472-891e-2d4d904f1ad6.pngPK 
     w�O\	��} } /             ��# images/bbfae99c-8036-4c5e-89fd-a87441410720.pngPK 
     w�O\d��   �   /             �+% images/a262aa33-74c4-460b-b0ad-c746896f6744.pngPK      �  �L%   